
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire _44061_;
  wire _44062_;
  wire _44063_;
  wire _44064_;
  wire _44065_;
  wire _44066_;
  wire _44067_;
  wire _44068_;
  wire _44069_;
  wire _44070_;
  wire _44071_;
  wire _44072_;
  wire _44073_;
  wire _44074_;
  wire _44075_;
  wire _44076_;
  wire _44077_;
  wire _44078_;
  wire _44079_;
  wire _44080_;
  wire _44081_;
  wire _44082_;
  wire _44083_;
  wire _44084_;
  wire _44085_;
  wire _44086_;
  wire _44087_;
  wire _44088_;
  wire _44089_;
  wire _44090_;
  wire _44091_;
  wire _44092_;
  wire _44093_;
  wire _44094_;
  wire _44095_;
  wire _44096_;
  wire _44097_;
  wire _44098_;
  wire _44099_;
  wire _44100_;
  wire _44101_;
  wire _44102_;
  wire _44103_;
  wire _44104_;
  wire _44105_;
  wire _44106_;
  wire _44107_;
  wire _44108_;
  wire _44109_;
  wire _44110_;
  wire _44111_;
  wire _44112_;
  wire _44113_;
  wire _44114_;
  wire _44115_;
  wire _44116_;
  wire _44117_;
  wire _44118_;
  wire _44119_;
  wire _44120_;
  wire _44121_;
  wire _44122_;
  wire _44123_;
  wire _44124_;
  wire _44125_;
  wire _44126_;
  wire _44127_;
  wire _44128_;
  wire _44129_;
  wire _44130_;
  wire _44131_;
  wire _44132_;
  wire _44133_;
  wire _44134_;
  wire _44135_;
  wire _44136_;
  wire _44137_;
  wire _44138_;
  wire _44139_;
  wire _44140_;
  wire _44141_;
  wire _44142_;
  wire _44143_;
  wire _44144_;
  wire _44145_;
  wire _44146_;
  wire _44147_;
  wire _44148_;
  wire _44149_;
  wire _44150_;
  wire _44151_;
  wire _44152_;
  wire _44153_;
  wire _44154_;
  wire _44155_;
  wire _44156_;
  wire _44157_;
  wire _44158_;
  wire _44159_;
  wire _44160_;
  wire _44161_;
  wire _44162_;
  wire _44163_;
  wire _44164_;
  wire _44165_;
  wire _44166_;
  wire _44167_;
  wire _44168_;
  wire _44169_;
  wire _44170_;
  wire _44171_;
  wire _44172_;
  wire _44173_;
  wire _44174_;
  wire _44175_;
  wire _44176_;
  wire _44177_;
  wire _44178_;
  wire _44179_;
  wire _44180_;
  wire _44181_;
  wire _44182_;
  wire _44183_;
  wire _44184_;
  wire _44185_;
  wire _44186_;
  wire _44187_;
  wire _44188_;
  wire _44189_;
  wire _44190_;
  wire _44191_;
  wire _44192_;
  wire _44193_;
  wire _44194_;
  wire _44195_;
  wire _44196_;
  wire _44197_;
  wire _44198_;
  wire _44199_;
  wire _44200_;
  wire _44201_;
  wire _44202_;
  wire _44203_;
  wire _44204_;
  wire _44205_;
  wire _44206_;
  wire _44207_;
  wire _44208_;
  wire _44209_;
  wire _44210_;
  wire _44211_;
  wire _44212_;
  wire _44213_;
  wire _44214_;
  wire _44215_;
  wire _44216_;
  wire _44217_;
  wire _44218_;
  wire _44219_;
  wire _44220_;
  wire _44221_;
  wire _44222_;
  wire _44223_;
  wire _44224_;
  wire _44225_;
  wire _44226_;
  wire _44227_;
  wire _44228_;
  wire _44229_;
  wire _44230_;
  wire _44231_;
  wire _44232_;
  wire _44233_;
  wire _44234_;
  wire _44235_;
  wire _44236_;
  wire _44237_;
  wire _44238_;
  wire _44239_;
  wire _44240_;
  wire _44241_;
  wire _44242_;
  wire _44243_;
  wire _44244_;
  wire _44245_;
  wire _44246_;
  wire _44247_;
  wire _44248_;
  wire _44249_;
  wire _44250_;
  wire _44251_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire [7:0] ie_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [6:0] \oc8051_golden_model_1.n0988 ;
  wire \oc8051_golden_model_1.n0989 ;
  wire \oc8051_golden_model_1.n0990 ;
  wire \oc8051_golden_model_1.n0991 ;
  wire \oc8051_golden_model_1.n0992 ;
  wire \oc8051_golden_model_1.n0993 ;
  wire \oc8051_golden_model_1.n0994 ;
  wire \oc8051_golden_model_1.n0995 ;
  wire \oc8051_golden_model_1.n0996 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire [7:0] \oc8051_golden_model_1.n1004 ;
  wire [7:0] \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire \oc8051_golden_model_1.n1018 ;
  wire \oc8051_golden_model_1.n1019 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire [7:0] \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1043 ;
  wire [7:0] \oc8051_golden_model_1.n1044 ;
  wire [3:0] \oc8051_golden_model_1.n1137 ;
  wire [3:0] \oc8051_golden_model_1.n1139 ;
  wire [3:0] \oc8051_golden_model_1.n1141 ;
  wire [3:0] \oc8051_golden_model_1.n1142 ;
  wire [3:0] \oc8051_golden_model_1.n1143 ;
  wire [3:0] \oc8051_golden_model_1.n1144 ;
  wire [3:0] \oc8051_golden_model_1.n1145 ;
  wire [3:0] \oc8051_golden_model_1.n1146 ;
  wire [3:0] \oc8051_golden_model_1.n1147 ;
  wire \oc8051_golden_model_1.n1194 ;
  wire \oc8051_golden_model_1.n1239 ;
  wire [8:0] \oc8051_golden_model_1.n1240 ;
  wire [8:0] \oc8051_golden_model_1.n1241 ;
  wire [7:0] \oc8051_golden_model_1.n1242 ;
  wire \oc8051_golden_model_1.n1243 ;
  wire [2:0] \oc8051_golden_model_1.n1244 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [1:0] \oc8051_golden_model_1.n1246 ;
  wire [7:0] \oc8051_golden_model_1.n1247 ;
  wire [6:0] \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1251 ;
  wire \oc8051_golden_model_1.n1252 ;
  wire \oc8051_golden_model_1.n1253 ;
  wire \oc8051_golden_model_1.n1254 ;
  wire \oc8051_golden_model_1.n1255 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [7:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1280 ;
  wire [7:0] \oc8051_golden_model_1.n1281 ;
  wire [15:0] \oc8051_golden_model_1.n1323 ;
  wire [7:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1328 ;
  wire \oc8051_golden_model_1.n1329 ;
  wire \oc8051_golden_model_1.n1330 ;
  wire \oc8051_golden_model_1.n1331 ;
  wire \oc8051_golden_model_1.n1332 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire \oc8051_golden_model_1.n1340 ;
  wire [7:0] \oc8051_golden_model_1.n1341 ;
  wire [8:0] \oc8051_golden_model_1.n1343 ;
  wire [8:0] \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire [3:0] \oc8051_golden_model_1.n1349 ;
  wire [4:0] \oc8051_golden_model_1.n1350 ;
  wire [4:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [8:0] \oc8051_golden_model_1.n1356 ;
  wire \oc8051_golden_model_1.n1364 ;
  wire [7:0] \oc8051_golden_model_1.n1365 ;
  wire [6:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1381 ;
  wire [7:0] \oc8051_golden_model_1.n1382 ;
  wire [8:0] \oc8051_golden_model_1.n1404 ;
  wire \oc8051_golden_model_1.n1405 ;
  wire [4:0] \oc8051_golden_model_1.n1410 ;
  wire \oc8051_golden_model_1.n1411 ;
  wire \oc8051_golden_model_1.n1419 ;
  wire [7:0] \oc8051_golden_model_1.n1420 ;
  wire [6:0] \oc8051_golden_model_1.n1421 ;
  wire \oc8051_golden_model_1.n1436 ;
  wire [7:0] \oc8051_golden_model_1.n1437 ;
  wire [8:0] \oc8051_golden_model_1.n1439 ;
  wire [8:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1442 ;
  wire [3:0] \oc8051_golden_model_1.n1443 ;
  wire [4:0] \oc8051_golden_model_1.n1444 ;
  wire [4:0] \oc8051_golden_model_1.n1446 ;
  wire \oc8051_golden_model_1.n1447 ;
  wire [8:0] \oc8051_golden_model_1.n1448 ;
  wire \oc8051_golden_model_1.n1455 ;
  wire [7:0] \oc8051_golden_model_1.n1456 ;
  wire [6:0] \oc8051_golden_model_1.n1457 ;
  wire \oc8051_golden_model_1.n1472 ;
  wire [7:0] \oc8051_golden_model_1.n1473 ;
  wire [8:0] \oc8051_golden_model_1.n1476 ;
  wire \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1484 ;
  wire [7:0] \oc8051_golden_model_1.n1485 ;
  wire [6:0] \oc8051_golden_model_1.n1486 ;
  wire [7:0] \oc8051_golden_model_1.n1487 ;
  wire [8:0] \oc8051_golden_model_1.n1489 ;
  wire [8:0] \oc8051_golden_model_1.n1491 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [4:0] \oc8051_golden_model_1.n1493 ;
  wire [4:0] \oc8051_golden_model_1.n1495 ;
  wire \oc8051_golden_model_1.n1496 ;
  wire [8:0] \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire [4:0] \oc8051_golden_model_1.n1524 ;
  wire \oc8051_golden_model_1.n1525 ;
  wire [7:0] \oc8051_golden_model_1.n1526 ;
  wire [6:0] \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [8:0] \oc8051_golden_model_1.n1530 ;
  wire \oc8051_golden_model_1.n1531 ;
  wire \oc8051_golden_model_1.n1538 ;
  wire [7:0] \oc8051_golden_model_1.n1539 ;
  wire [6:0] \oc8051_golden_model_1.n1540 ;
  wire [7:0] \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [6:0] \oc8051_golden_model_1.n1543 ;
  wire [7:0] \oc8051_golden_model_1.n1544 ;
  wire [8:0] \oc8051_golden_model_1.n1547 ;
  wire [8:0] \oc8051_golden_model_1.n1548 ;
  wire [7:0] \oc8051_golden_model_1.n1549 ;
  wire [7:0] \oc8051_golden_model_1.n1550 ;
  wire [6:0] \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1552 ;
  wire \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire \oc8051_golden_model_1.n1555 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1559 ;
  wire \oc8051_golden_model_1.n1566 ;
  wire [7:0] \oc8051_golden_model_1.n1567 ;
  wire [7:0] \oc8051_golden_model_1.n1568 ;
  wire [8:0] \oc8051_golden_model_1.n1571 ;
  wire [8:0] \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire [4:0] \oc8051_golden_model_1.n1575 ;
  wire [4:0] \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1585 ;
  wire [7:0] \oc8051_golden_model_1.n1586 ;
  wire [6:0] \oc8051_golden_model_1.n1587 ;
  wire \oc8051_golden_model_1.n1602 ;
  wire [7:0] \oc8051_golden_model_1.n1603 ;
  wire [8:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1608 ;
  wire [4:0] \oc8051_golden_model_1.n1610 ;
  wire \oc8051_golden_model_1.n1611 ;
  wire \oc8051_golden_model_1.n1618 ;
  wire [7:0] \oc8051_golden_model_1.n1619 ;
  wire [6:0] \oc8051_golden_model_1.n1620 ;
  wire \oc8051_golden_model_1.n1635 ;
  wire [7:0] \oc8051_golden_model_1.n1636 ;
  wire [8:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1641 ;
  wire [4:0] \oc8051_golden_model_1.n1643 ;
  wire \oc8051_golden_model_1.n1644 ;
  wire \oc8051_golden_model_1.n1651 ;
  wire [7:0] \oc8051_golden_model_1.n1652 ;
  wire [6:0] \oc8051_golden_model_1.n1653 ;
  wire \oc8051_golden_model_1.n1668 ;
  wire [7:0] \oc8051_golden_model_1.n1669 ;
  wire [8:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1674 ;
  wire [4:0] \oc8051_golden_model_1.n1676 ;
  wire \oc8051_golden_model_1.n1677 ;
  wire \oc8051_golden_model_1.n1684 ;
  wire [7:0] \oc8051_golden_model_1.n1685 ;
  wire [6:0] \oc8051_golden_model_1.n1686 ;
  wire \oc8051_golden_model_1.n1701 ;
  wire [7:0] \oc8051_golden_model_1.n1702 ;
  wire [7:0] \oc8051_golden_model_1.n1727 ;
  wire [6:0] \oc8051_golden_model_1.n1728 ;
  wire [7:0] \oc8051_golden_model_1.n1729 ;
  wire \oc8051_golden_model_1.n1784 ;
  wire [7:0] \oc8051_golden_model_1.n1785 ;
  wire \oc8051_golden_model_1.n1801 ;
  wire [7:0] \oc8051_golden_model_1.n1802 ;
  wire \oc8051_golden_model_1.n1818 ;
  wire [7:0] \oc8051_golden_model_1.n1819 ;
  wire \oc8051_golden_model_1.n1835 ;
  wire [7:0] \oc8051_golden_model_1.n1836 ;
  wire [7:0] \oc8051_golden_model_1.n1859 ;
  wire [6:0] \oc8051_golden_model_1.n1860 ;
  wire [7:0] \oc8051_golden_model_1.n1861 ;
  wire \oc8051_golden_model_1.n1916 ;
  wire [7:0] \oc8051_golden_model_1.n1917 ;
  wire \oc8051_golden_model_1.n1933 ;
  wire [7:0] \oc8051_golden_model_1.n1934 ;
  wire \oc8051_golden_model_1.n1950 ;
  wire [7:0] \oc8051_golden_model_1.n1951 ;
  wire \oc8051_golden_model_1.n1967 ;
  wire [7:0] \oc8051_golden_model_1.n1968 ;
  wire \oc8051_golden_model_1.n2065 ;
  wire [7:0] \oc8051_golden_model_1.n2066 ;
  wire \oc8051_golden_model_1.n2082 ;
  wire [7:0] \oc8051_golden_model_1.n2083 ;
  wire \oc8051_golden_model_1.n2099 ;
  wire [7:0] \oc8051_golden_model_1.n2100 ;
  wire \oc8051_golden_model_1.n2116 ;
  wire [7:0] \oc8051_golden_model_1.n2117 ;
  wire \oc8051_golden_model_1.n2121 ;
  wire [6:0] \oc8051_golden_model_1.n2122 ;
  wire [7:0] \oc8051_golden_model_1.n2123 ;
  wire [6:0] \oc8051_golden_model_1.n2124 ;
  wire [7:0] \oc8051_golden_model_1.n2125 ;
  wire \oc8051_golden_model_1.n2140 ;
  wire [7:0] \oc8051_golden_model_1.n2141 ;
  wire \oc8051_golden_model_1.n2180 ;
  wire [7:0] \oc8051_golden_model_1.n2181 ;
  wire [6:0] \oc8051_golden_model_1.n2182 ;
  wire [7:0] \oc8051_golden_model_1.n2183 ;
  wire [3:0] \oc8051_golden_model_1.n2190 ;
  wire \oc8051_golden_model_1.n2191 ;
  wire [7:0] \oc8051_golden_model_1.n2192 ;
  wire [6:0] \oc8051_golden_model_1.n2193 ;
  wire \oc8051_golden_model_1.n2208 ;
  wire [7:0] \oc8051_golden_model_1.n2209 ;
  wire [7:0] \oc8051_golden_model_1.n2421 ;
  wire \oc8051_golden_model_1.n2424 ;
  wire \oc8051_golden_model_1.n2426 ;
  wire \oc8051_golden_model_1.n2432 ;
  wire [7:0] \oc8051_golden_model_1.n2433 ;
  wire [6:0] \oc8051_golden_model_1.n2434 ;
  wire \oc8051_golden_model_1.n2449 ;
  wire [7:0] \oc8051_golden_model_1.n2450 ;
  wire \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2456 ;
  wire \oc8051_golden_model_1.n2462 ;
  wire [7:0] \oc8051_golden_model_1.n2463 ;
  wire [6:0] \oc8051_golden_model_1.n2464 ;
  wire \oc8051_golden_model_1.n2479 ;
  wire [7:0] \oc8051_golden_model_1.n2480 ;
  wire \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2486 ;
  wire \oc8051_golden_model_1.n2492 ;
  wire [7:0] \oc8051_golden_model_1.n2493 ;
  wire [6:0] \oc8051_golden_model_1.n2494 ;
  wire \oc8051_golden_model_1.n2509 ;
  wire [7:0] \oc8051_golden_model_1.n2510 ;
  wire \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2516 ;
  wire \oc8051_golden_model_1.n2522 ;
  wire [7:0] \oc8051_golden_model_1.n2523 ;
  wire [6:0] \oc8051_golden_model_1.n2524 ;
  wire \oc8051_golden_model_1.n2539 ;
  wire [7:0] \oc8051_golden_model_1.n2540 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire [7:0] \oc8051_golden_model_1.n2545 ;
  wire [7:0] \oc8051_golden_model_1.n2546 ;
  wire [6:0] \oc8051_golden_model_1.n2547 ;
  wire [7:0] \oc8051_golden_model_1.n2548 ;
  wire [15:0] \oc8051_golden_model_1.n2552 ;
  wire \oc8051_golden_model_1.n2558 ;
  wire [7:0] \oc8051_golden_model_1.n2559 ;
  wire [6:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2575 ;
  wire [7:0] \oc8051_golden_model_1.n2576 ;
  wire \oc8051_golden_model_1.n2579 ;
  wire [7:0] \oc8051_golden_model_1.n2580 ;
  wire [6:0] \oc8051_golden_model_1.n2581 ;
  wire [7:0] \oc8051_golden_model_1.n2582 ;
  wire \oc8051_golden_model_1.n2614 ;
  wire [7:0] \oc8051_golden_model_1.n2615 ;
  wire [6:0] \oc8051_golden_model_1.n2616 ;
  wire [7:0] \oc8051_golden_model_1.n2617 ;
  wire \oc8051_golden_model_1.n2622 ;
  wire [7:0] \oc8051_golden_model_1.n2623 ;
  wire [6:0] \oc8051_golden_model_1.n2624 ;
  wire [7:0] \oc8051_golden_model_1.n2625 ;
  wire \oc8051_golden_model_1.n2630 ;
  wire [7:0] \oc8051_golden_model_1.n2631 ;
  wire [6:0] \oc8051_golden_model_1.n2632 ;
  wire [7:0] \oc8051_golden_model_1.n2633 ;
  wire \oc8051_golden_model_1.n2638 ;
  wire [7:0] \oc8051_golden_model_1.n2639 ;
  wire [6:0] \oc8051_golden_model_1.n2640 ;
  wire [7:0] \oc8051_golden_model_1.n2641 ;
  wire \oc8051_golden_model_1.n2646 ;
  wire [7:0] \oc8051_golden_model_1.n2647 ;
  wire [6:0] \oc8051_golden_model_1.n2648 ;
  wire [7:0] \oc8051_golden_model_1.n2649 ;
  wire [7:0] \oc8051_golden_model_1.n2674 ;
  wire [6:0] \oc8051_golden_model_1.n2675 ;
  wire [7:0] \oc8051_golden_model_1.n2676 ;
  wire [3:0] \oc8051_golden_model_1.n2677 ;
  wire [7:0] \oc8051_golden_model_1.n2678 ;
  wire \oc8051_golden_model_1.n2679 ;
  wire \oc8051_golden_model_1.n2680 ;
  wire \oc8051_golden_model_1.n2681 ;
  wire \oc8051_golden_model_1.n2682 ;
  wire \oc8051_golden_model_1.n2683 ;
  wire \oc8051_golden_model_1.n2684 ;
  wire \oc8051_golden_model_1.n2685 ;
  wire \oc8051_golden_model_1.n2686 ;
  wire \oc8051_golden_model_1.n2693 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [6:0] \oc8051_golden_model_1.n2715 ;
  wire [7:0] \oc8051_golden_model_1.n2731 ;
  wire \oc8051_golden_model_1.n2732 ;
  wire \oc8051_golden_model_1.n2733 ;
  wire \oc8051_golden_model_1.n2734 ;
  wire \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2736 ;
  wire \oc8051_golden_model_1.n2737 ;
  wire \oc8051_golden_model_1.n2738 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire \oc8051_golden_model_1.n2746 ;
  wire [7:0] \oc8051_golden_model_1.n2747 ;
  wire \oc8051_golden_model_1.n2748 ;
  wire \oc8051_golden_model_1.n2749 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2762 ;
  wire [7:0] \oc8051_golden_model_1.n2763 ;
  wire [7:0] \oc8051_golden_model_1.n2795 ;
  wire [6:0] \oc8051_golden_model_1.n2796 ;
  wire [7:0] \oc8051_golden_model_1.n2797 ;
  wire \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire [6:0] \oc8051_golden_model_1.n2818 ;
  wire \oc8051_golden_model_1.n2833 ;
  wire [7:0] \oc8051_golden_model_1.n2834 ;
  wire [7:0] \oc8051_golden_model_1.n2838 ;
  wire [3:0] \oc8051_golden_model_1.n2839 ;
  wire [7:0] \oc8051_golden_model_1.n2840 ;
  wire \oc8051_golden_model_1.n2841 ;
  wire \oc8051_golden_model_1.n2842 ;
  wire \oc8051_golden_model_1.n2843 ;
  wire \oc8051_golden_model_1.n2844 ;
  wire \oc8051_golden_model_1.n2845 ;
  wire \oc8051_golden_model_1.n2846 ;
  wire \oc8051_golden_model_1.n2847 ;
  wire \oc8051_golden_model_1.n2848 ;
  wire \oc8051_golden_model_1.n2855 ;
  wire [7:0] \oc8051_golden_model_1.n2856 ;
  wire \oc8051_golden_model_1.n2874 ;
  wire [7:0] \oc8051_golden_model_1.n2875 ;
  wire \oc8051_golden_model_1.n2891 ;
  wire [7:0] \oc8051_golden_model_1.n2892 ;
  wire [7:0] \oc8051_golden_model_1.n2893 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  wire property_invalid_psw_1_r;
  output property_invalid_sp;
  wire property_invalid_sp_1_r;
  wire [7:0] psw_impl;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_41991_, rst);
  not (_15613_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_15624_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15635_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15624_);
  and (_15646_, _15635_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_15657_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15624_);
  and (_15668_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _15624_);
  nor (_15679_, _15668_, _15657_);
  and (_15690_, _15679_, _15646_);
  nor (_15701_, _15690_, _15613_);
  and (_15712_, _15613_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15723_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_15734_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _15723_);
  nor (_15745_, _15734_, _15712_);
  not (_15756_, _15745_);
  and (_15767_, _15756_, _15690_);
  or (_15778_, _15767_, _15701_);
  and (_22423_, _15778_, _41991_);
  nor (_15799_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15810_, _15799_);
  and (_15821_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_15832_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_15842_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_15853_, _15842_);
  not (_15864_, _15734_);
  nor (_15875_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_15886_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_15897_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _15886_);
  nor (_15908_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_15919_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_15930_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _15919_);
  nor (_15941_, _15930_, _15908_);
  nor (_15952_, _15941_, _15897_);
  not (_15963_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_15974_, _15897_, _15963_);
  nor (_15985_, _15974_, _15952_);
  and (_15996_, _15985_, _15875_);
  not (_16007_, _15996_);
  and (_16018_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16029_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_16040_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_16051_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _16040_);
  and (_16062_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_16073_, _16062_, _16029_);
  and (_16084_, _16073_, _16007_);
  nor (_16095_, _16084_, _15864_);
  not (_16106_, _15712_);
  nor (_16117_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_16128_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _15919_);
  nor (_16139_, _16128_, _16117_);
  nor (_16150_, _16139_, _15897_);
  not (_16161_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_16171_, _15897_, _16161_);
  nor (_16182_, _16171_, _16150_);
  and (_16193_, _16182_, _15875_);
  not (_16204_, _16193_);
  and (_16215_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_16226_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_16237_, _16226_, _16215_);
  and (_16248_, _16237_, _16204_);
  nor (_16259_, _16248_, _16106_);
  nor (_16270_, _16259_, _16095_);
  nor (_16281_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_16292_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _15919_);
  nor (_16303_, _16292_, _16281_);
  nor (_16314_, _16303_, _15897_);
  not (_16325_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_16336_, _15897_, _16325_);
  nor (_16347_, _16336_, _16314_);
  and (_16358_, _16347_, _15875_);
  not (_16369_, _16358_);
  and (_16380_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_16391_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_16402_, _16391_, _16380_);
  and (_16413_, _16402_, _16369_);
  nor (_16424_, _16413_, _15756_);
  nor (_16435_, _16424_, _15799_);
  and (_16446_, _16435_, _16270_);
  nor (_16457_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_16468_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _15919_);
  nor (_16479_, _16468_, _16457_);
  nor (_16489_, _16479_, _15897_);
  not (_16500_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_16511_, _15897_, _16500_);
  nor (_16522_, _16511_, _16489_);
  and (_16544_, _16522_, _15875_);
  not (_16545_, _16544_);
  and (_16556_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_16567_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16578_, _16567_, _16556_);
  and (_16589_, _16578_, _16545_);
  and (_16600_, _16589_, _15799_);
  nor (_16611_, _16600_, _16446_);
  not (_16622_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16633_, _16622_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16644_, _16633_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16655_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_16666_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16677_, _16666_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16688_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_16699_, _16688_, _16655_);
  nor (_16710_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16721_, _16710_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16732_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_16743_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16754_, _16633_, _16743_);
  and (_16765_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_16776_, _16765_, _16732_);
  and (_16787_, _16776_, _16699_);
  and (_16798_, _16710_, _16622_);
  and (_16808_, _16798_, _16522_);
  and (_16819_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16830_, _16819_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16841_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_16852_, _16819_, _16743_);
  and (_16863_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16874_, _16863_, _16841_);
  not (_16885_, _16874_);
  nor (_16896_, _16885_, _16808_);
  and (_16907_, _16896_, _16787_);
  not (_16918_, _16907_);
  and (_16929_, _16918_, _16611_);
  not (_16940_, _16929_);
  nor (_16951_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_16962_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _15919_);
  nor (_16973_, _16962_, _16951_);
  nor (_16984_, _16973_, _15897_);
  not (_16995_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_17006_, _15897_, _16995_);
  nor (_17017_, _17006_, _16984_);
  and (_17028_, _17017_, _15875_);
  not (_17039_, _17028_);
  and (_17050_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_17061_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_17072_, _17061_, _17050_);
  and (_17083_, _17072_, _17039_);
  nor (_17094_, _17083_, _15864_);
  nor (_17105_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_17116_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _15919_);
  nor (_17127_, _17116_, _17105_);
  nor (_17138_, _17127_, _15897_);
  not (_17148_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_17159_, _15897_, _17148_);
  nor (_17170_, _17159_, _17138_);
  and (_17181_, _17170_, _15875_);
  not (_17192_, _17181_);
  and (_17203_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_17214_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17225_, _17214_, _17203_);
  and (_17235_, _17225_, _17192_);
  nor (_17246_, _17235_, _16106_);
  nor (_17267_, _17246_, _17094_);
  nor (_17268_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_17289_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _15919_);
  nor (_17290_, _17289_, _17268_);
  nor (_17301_, _17290_, _15897_);
  not (_17312_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_17323_, _15897_, _17312_);
  nor (_17333_, _17323_, _17301_);
  and (_17344_, _17333_, _15875_);
  not (_17355_, _17344_);
  and (_17366_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_17377_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_17388_, _17377_, _17366_);
  and (_17399_, _17388_, _17355_);
  nor (_17410_, _17399_, _15756_);
  nor (_17420_, _17410_, _15799_);
  and (_17431_, _17420_, _17267_);
  nor (_17442_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_17453_, _15919_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_17464_, _17453_, _17442_);
  nor (_17475_, _17464_, _15897_);
  not (_17486_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_17497_, _15897_, _17486_);
  nor (_17508_, _17497_, _17475_);
  and (_17518_, _17508_, _15875_);
  not (_17529_, _17518_);
  and (_17540_, _16018_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_17551_, _16051_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_17562_, _17551_, _17540_);
  and (_17573_, _17562_, _17529_);
  and (_17584_, _17573_, _15799_);
  or (_17595_, _17584_, _17431_);
  and (_17606_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_17616_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_17627_, _17616_, _17606_);
  and (_17638_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_17649_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_17660_, _17649_, _17638_);
  and (_17671_, _17660_, _17627_);
  and (_17682_, _17508_, _16798_);
  and (_17693_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_17703_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_17714_, _17703_, _17693_);
  not (_17725_, _17714_);
  nor (_17736_, _17725_, _17682_);
  and (_17747_, _17736_, _17671_);
  nor (_17758_, _17747_, _17595_);
  and (_17769_, _17758_, _16940_);
  not (_17780_, _17769_);
  and (_17791_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_17801_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_17812_, _17801_, _17791_);
  and (_17823_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_17834_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_17845_, _17834_, _17823_);
  and (_17856_, _17845_, _17812_);
  and (_17867_, _17170_, _16798_);
  and (_17878_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_17888_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17899_, _17888_, _17878_);
  not (_17910_, _17899_);
  nor (_17921_, _17910_, _17867_);
  and (_17932_, _17921_, _17856_);
  nor (_17943_, _17932_, _17595_);
  and (_17954_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_17965_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_17976_, _17965_, _17954_);
  and (_17986_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_17997_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_18008_, _17997_, _17986_);
  and (_18019_, _18008_, _17976_);
  and (_18030_, _16798_, _16182_);
  and (_18041_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_18052_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_18063_, _18052_, _18041_);
  not (_18073_, _18063_);
  nor (_18084_, _18073_, _18030_);
  and (_18095_, _18084_, _18019_);
  not (_18106_, _18095_);
  and (_18117_, _18106_, _16611_);
  and (_18128_, _17943_, _18117_);
  and (_18139_, _16918_, _18128_);
  nor (_18150_, _16929_, _18128_);
  nor (_18161_, _18150_, _18139_);
  and (_18171_, _18161_, _17943_);
  and (_18182_, _17758_, _16929_);
  nor (_18193_, _16907_, _17595_);
  not (_18204_, _17747_);
  and (_18215_, _18204_, _16611_);
  nor (_18226_, _18215_, _18193_);
  nor (_18237_, _18226_, _18182_);
  and (_18248_, _18237_, _18171_);
  nor (_18258_, _18237_, _18171_);
  nor (_18269_, _18258_, _18248_);
  and (_18280_, _18269_, _18139_);
  nor (_18291_, _18280_, _18248_);
  nor (_18302_, _18291_, _17780_);
  nor (_18313_, _17595_, _18095_);
  and (_18324_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_18335_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_18346_, _18335_, _18324_);
  and (_18356_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_18367_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_18378_, _18367_, _18356_);
  and (_18389_, _18378_, _18346_);
  and (_18400_, _17017_, _16798_);
  and (_18411_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_18422_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_18433_, _18422_, _18411_);
  not (_18444_, _18433_);
  nor (_18454_, _18444_, _18400_);
  and (_18465_, _18454_, _18389_);
  not (_18476_, _18465_);
  and (_18487_, _18476_, _16611_);
  and (_18498_, _18487_, _18313_);
  not (_18509_, _17932_);
  and (_18520_, _18509_, _16611_);
  nor (_18531_, _18520_, _18313_);
  nor (_18542_, _18531_, _18128_);
  and (_18552_, _18542_, _18498_);
  nor (_18563_, _16929_, _17943_);
  nor (_18574_, _18563_, _18171_);
  and (_18585_, _18574_, _18552_);
  nor (_18596_, _18269_, _18139_);
  nor (_18607_, _18596_, _18280_);
  and (_18618_, _18607_, _18585_);
  nor (_18629_, _18607_, _18585_);
  nor (_18640_, _18629_, _18618_);
  not (_18651_, _18640_);
  and (_18662_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_18672_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_18683_, _18672_, _18662_);
  and (_18694_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_18705_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_18716_, _18705_, _18694_);
  and (_18727_, _18716_, _18683_);
  and (_18738_, _17333_, _16798_);
  and (_18749_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_18760_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_18771_, _18760_, _18749_);
  not (_18781_, _18771_);
  nor (_18792_, _18781_, _18738_);
  and (_18803_, _18792_, _18727_);
  nor (_18814_, _18803_, _17595_);
  and (_18825_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_18836_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_18847_, _18836_, _18825_);
  and (_18858_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_18869_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_18880_, _18869_, _18858_);
  and (_18891_, _18880_, _18847_);
  and (_18901_, _16798_, _15985_);
  and (_18912_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_18923_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_18934_, _18923_, _18912_);
  not (_18945_, _18934_);
  nor (_18956_, _18945_, _18901_);
  and (_18967_, _18956_, _18891_);
  not (_18978_, _18967_);
  and (_18989_, _18978_, _16611_);
  and (_19000_, _18989_, _18814_);
  not (_19011_, _18803_);
  and (_19021_, _19011_, _16611_);
  not (_19032_, _19021_);
  nor (_19043_, _18967_, _17595_);
  and (_19054_, _19043_, _19032_);
  and (_19065_, _19054_, _18487_);
  nor (_19076_, _19065_, _19000_);
  nor (_19087_, _18465_, _17595_);
  nor (_19098_, _19087_, _18117_);
  nor (_19109_, _19098_, _18498_);
  not (_19120_, _19109_);
  nor (_19130_, _19120_, _19076_);
  nor (_19141_, _18542_, _18498_);
  nor (_19152_, _19141_, _18552_);
  and (_19163_, _19152_, _19130_);
  nor (_19174_, _18574_, _18552_);
  nor (_19185_, _19174_, _18585_);
  and (_19196_, _19185_, _19163_);
  and (_19207_, _16644_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_19218_, _16677_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_19229_, _19218_, _19207_);
  and (_19240_, _16721_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_19250_, _16754_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_19261_, _19250_, _19240_);
  and (_19272_, _19261_, _19229_);
  and (_19283_, _16798_, _16347_);
  and (_19294_, _16852_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_19305_, _16830_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_19316_, _19305_, _19294_);
  not (_19327_, _19316_);
  nor (_19338_, _19327_, _19283_);
  and (_19348_, _19338_, _19272_);
  nor (_19359_, _19348_, _17595_);
  and (_19370_, _19359_, _19021_);
  nor (_19381_, _18989_, _18814_);
  nor (_19392_, _19381_, _19000_);
  and (_19403_, _19392_, _19370_);
  nor (_19414_, _19054_, _18487_);
  nor (_19425_, _19414_, _19065_);
  and (_19436_, _19425_, _19403_);
  and (_19447_, _19120_, _19076_);
  nor (_19458_, _19447_, _19130_);
  and (_19468_, _19458_, _19436_);
  nor (_19479_, _19152_, _19130_);
  nor (_19490_, _19479_, _19163_);
  and (_19501_, _19490_, _19468_);
  nor (_19512_, _19185_, _19163_);
  nor (_19523_, _19512_, _19196_);
  and (_19534_, _19523_, _19501_);
  nor (_19545_, _19534_, _19196_);
  nor (_19556_, _19545_, _18651_);
  nor (_19567_, _19556_, _18618_);
  and (_19577_, _18291_, _17780_);
  nor (_19588_, _19577_, _18302_);
  not (_19599_, _19588_);
  nor (_19610_, _19599_, _19567_);
  or (_19621_, _19610_, _18182_);
  nor (_19632_, _19621_, _18302_);
  nor (_19643_, _19632_, _15853_);
  and (_19654_, _19632_, _15853_);
  nor (_19665_, _19654_, _19643_);
  not (_19676_, _19665_);
  and (_19687_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_19697_, _19599_, _19567_);
  nor (_19708_, _19697_, _19610_);
  and (_19719_, _19708_, _19687_);
  and (_19730_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_19741_, _19545_, _18651_);
  nor (_19752_, _19741_, _19556_);
  and (_19763_, _19752_, _19730_);
  nor (_19774_, _19752_, _19730_);
  nor (_19785_, _19774_, _19763_);
  not (_19796_, _19785_);
  and (_19807_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_19817_, _19523_, _19501_);
  nor (_19828_, _19817_, _19534_);
  and (_19839_, _19828_, _19807_);
  nor (_19850_, _19828_, _19807_);
  nor (_19861_, _19850_, _19839_);
  not (_19872_, _19861_);
  and (_19883_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_19894_, _19490_, _19468_);
  nor (_19905_, _19894_, _19501_);
  and (_19916_, _19905_, _19883_);
  nor (_19926_, _19905_, _19883_);
  nor (_19937_, _19926_, _19916_);
  not (_19948_, _19937_);
  and (_19959_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_19970_, _19458_, _19436_);
  nor (_19981_, _19970_, _19468_);
  and (_19992_, _19981_, _19959_);
  and (_20003_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_20014_, _19425_, _19403_);
  nor (_20025_, _20014_, _19436_);
  and (_20035_, _20025_, _20003_);
  and (_20046_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_20057_, _19392_, _19370_);
  nor (_20068_, _20057_, _19403_);
  and (_20079_, _20068_, _20046_);
  nor (_20090_, _20025_, _20003_);
  nor (_20101_, _20090_, _20035_);
  and (_20112_, _20101_, _20079_);
  nor (_20123_, _20112_, _20035_);
  not (_20134_, _20123_);
  nor (_20145_, _19981_, _19959_);
  nor (_20156_, _20145_, _19992_);
  and (_20166_, _20156_, _20134_);
  nor (_20177_, _20166_, _19992_);
  nor (_20188_, _20177_, _19948_);
  nor (_20199_, _20188_, _19916_);
  nor (_20210_, _20199_, _19872_);
  nor (_20221_, _20210_, _19839_);
  nor (_20232_, _20221_, _19796_);
  nor (_20243_, _20232_, _19763_);
  nor (_20254_, _19708_, _19687_);
  nor (_20265_, _20254_, _19719_);
  not (_20276_, _20265_);
  nor (_20287_, _20276_, _20243_);
  nor (_20297_, _20287_, _19719_);
  nor (_20308_, _20297_, _19676_);
  nor (_20319_, _20308_, _19643_);
  not (_20330_, _20319_);
  and (_20341_, _20330_, _15832_);
  and (_20352_, _20341_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_20363_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_20374_, _20363_, _20352_);
  and (_20385_, _20374_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_20396_, _20385_, _15821_);
  and (_20407_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20417_, _20407_, _20396_);
  and (_20428_, _20396_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_20439_, _20428_, _20417_);
  and (_24609_, _20439_, _41991_);
  nor (_20460_, _15690_, _15723_);
  and (_20471_, _15690_, _15723_);
  or (_20482_, _20471_, _20460_);
  and (_02454_, _20482_, _41991_);
  not (_20503_, _19348_);
  and (_20514_, _20503_, _16611_);
  and (_02649_, _20514_, _41991_);
  nor (_20535_, _19359_, _19021_);
  nor (_20545_, _20535_, _19370_);
  and (_02844_, _20545_, _41991_);
  nor (_20566_, _20068_, _20046_);
  nor (_20577_, _20566_, _20079_);
  and (_03045_, _20577_, _41991_);
  nor (_20598_, _20101_, _20079_);
  nor (_20609_, _20598_, _20112_);
  and (_03256_, _20609_, _41991_);
  nor (_20630_, _20156_, _20134_);
  nor (_20641_, _20630_, _20166_);
  and (_03457_, _20641_, _41991_);
  and (_20661_, _20177_, _19948_);
  nor (_20672_, _20661_, _20188_);
  and (_03658_, _20672_, _41991_);
  and (_20693_, _20199_, _19872_);
  nor (_20704_, _20693_, _20210_);
  and (_03859_, _20704_, _41991_);
  and (_20725_, _20221_, _19796_);
  nor (_20736_, _20725_, _20232_);
  and (_04060_, _20736_, _41991_);
  and (_20757_, _20276_, _20243_);
  nor (_20768_, _20757_, _20287_);
  and (_04161_, _20768_, _41991_);
  and (_20788_, _20297_, _19676_);
  nor (_20799_, _20788_, _20308_);
  and (_04262_, _20799_, _41991_);
  nor (_20820_, _20330_, _15832_);
  nor (_20831_, _20820_, _20341_);
  and (_04363_, _20831_, _41991_);
  and (_20852_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_20863_, _20852_, _20341_);
  nor (_20874_, _20863_, _20352_);
  and (_04464_, _20874_, _41991_);
  nor (_20895_, _20363_, _20352_);
  nor (_20905_, _20895_, _20374_);
  and (_04565_, _20905_, _41991_);
  and (_20926_, _15810_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_20937_, _20926_, _20374_);
  nor (_20948_, _20937_, _20385_);
  and (_04666_, _20948_, _41991_);
  nor (_20969_, _20385_, _15821_);
  nor (_20980_, _20969_, _20396_);
  and (_04767_, _20980_, _41991_);
  and (_21001_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15624_);
  nor (_21011_, _21001_, _15635_);
  not (_21022_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_21033_, _15657_, _21022_);
  and (_21044_, _21033_, _21011_);
  and (_21055_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_21066_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21077_, _21055_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21088_, _21077_, _21066_);
  and (_00850_, _21088_, _41991_);
  and (_00881_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _41991_);
  not (_21118_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_21129_, _17399_, _21118_);
  and (_21140_, _17083_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21151_, _21140_, _21129_);
  nor (_21162_, _21151_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21173_, _17235_, _21118_);
  and (_21184_, _17573_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_21195_, _21184_, _21173_);
  and (_21206_, _21195_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_21217_, _21206_, _21162_);
  nor (_21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_21238_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and (_21249_, _21227_, _17747_);
  nor (_21260_, _21249_, _21238_);
  not (_21271_, _21260_);
  and (_21282_, _16413_, _21118_);
  and (_21293_, _16084_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21304_, _21293_, _21282_);
  nor (_21315_, _21304_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21326_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21337_, _16248_, _21118_);
  and (_21347_, _16589_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21358_, _21347_, _21337_);
  nor (_21369_, _21358_, _21326_);
  nor (_21380_, _21369_, _21315_);
  nor (_21391_, _21380_, _21271_);
  and (_21402_, _21380_, _21271_);
  nor (_21413_, _21402_, _21391_);
  nor (_21424_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_21435_, _21227_, _16907_);
  nor (_21446_, _21435_, _21424_);
  not (_21456_, _21446_);
  nor (_21478_, _17399_, _21118_);
  nor (_21490_, _21478_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21502_, _17083_, _21118_);
  and (_21514_, _17235_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21526_, _21514_, _21502_);
  nor (_21538_, _21526_, _21326_);
  nor (_21539_, _21538_, _21490_);
  nor (_21550_, _21539_, _21456_);
  and (_21561_, _21539_, _21456_);
  nor (_21571_, _21561_, _21550_);
  not (_21582_, _21571_);
  and (_21593_, _21227_, _17932_);
  nor (_21604_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor (_21615_, _21604_, _21593_);
  not (_21626_, _21615_);
  nor (_21637_, _16413_, _21118_);
  nor (_21648_, _21637_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21659_, _16084_, _21118_);
  and (_21670_, _16248_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21680_, _21670_, _21659_);
  nor (_21691_, _21680_, _21326_);
  nor (_21702_, _21691_, _21648_);
  nor (_21713_, _21702_, _21626_);
  and (_21724_, _21702_, _21626_);
  nor (_21735_, _21724_, _21713_);
  not (_21746_, _21735_);
  and (_21757_, _21151_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21768_, _21757_);
  nor (_21779_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_21789_, _21227_, _18095_);
  nor (_21800_, _21789_, _21779_);
  and (_21811_, _21800_, _21768_);
  and (_21822_, _21304_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21833_, _21822_);
  and (_21844_, _21227_, _18465_);
  nor (_21855_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_21866_, _21855_, _21844_);
  and (_21877_, _21866_, _21833_);
  nor (_21888_, _21866_, _21833_);
  nor (_21898_, _21888_, _21877_);
  not (_21909_, _21898_);
  and (_21920_, _21478_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21931_, _21920_);
  and (_21942_, _21227_, _18967_);
  nor (_21953_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_21964_, _21953_, _21942_);
  and (_21975_, _21964_, _21931_);
  and (_21986_, _21637_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21997_, _21986_);
  and (_22007_, _21227_, _18803_);
  nor (_22018_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  nor (_22029_, _22018_, _22007_);
  nor (_22050_, _22029_, _21997_);
  not (_22051_, _22050_);
  nor (_22062_, _21964_, _21931_);
  nor (_22073_, _22062_, _21975_);
  and (_22084_, _22073_, _22051_);
  nor (_22095_, _22084_, _21975_);
  nor (_22106_, _22095_, _21909_);
  nor (_22116_, _22106_, _21877_);
  nor (_22127_, _21800_, _21768_);
  nor (_22138_, _22127_, _21811_);
  not (_22149_, _22138_);
  nor (_22160_, _22149_, _22116_);
  nor (_22171_, _22160_, _21811_);
  nor (_22182_, _22171_, _21746_);
  nor (_22193_, _22182_, _21713_);
  nor (_22204_, _22193_, _21582_);
  nor (_22215_, _22204_, _21550_);
  not (_22225_, _22215_);
  and (_22236_, _22225_, _21413_);
  or (_22247_, _22236_, _21391_);
  and (_22258_, _17573_, _16589_);
  or (_22269_, _22258_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_22280_, _21526_);
  and (_22291_, _21195_, _22280_);
  nor (_22313_, _21680_, _21358_);
  and (_22314_, _22313_, _22291_);
  or (_22325_, _22314_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_22335_, _22325_, _22269_);
  and (_22346_, _22335_, _22247_);
  and (_22357_, _22346_, _21217_);
  nor (_22368_, _22225_, _21413_);
  or (_22379_, _22368_, _22236_);
  and (_22390_, _22379_, _22357_);
  nor (_22401_, _22357_, _21260_);
  nor (_22412_, _22401_, _22390_);
  not (_22424_, _22412_);
  and (_22435_, _22412_, _21217_);
  not (_22446_, _21380_);
  and (_22456_, _22193_, _21582_);
  or (_22467_, _22456_, _22204_);
  and (_22478_, _22467_, _22357_);
  nor (_22489_, _22357_, _21446_);
  nor (_22500_, _22489_, _22478_);
  and (_22511_, _22500_, _22446_);
  nor (_22522_, _22500_, _22446_);
  nor (_22533_, _22522_, _22511_);
  not (_22544_, _22533_);
  not (_22554_, _21539_);
  nor (_22565_, _22357_, _21626_);
  and (_22576_, _22171_, _21746_);
  nor (_22587_, _22576_, _22182_);
  and (_22598_, _22587_, _22357_);
  or (_22609_, _22598_, _22565_);
  and (_22620_, _22609_, _22554_);
  nor (_22631_, _22609_, _22554_);
  not (_22642_, _21702_);
  and (_22653_, _22149_, _22116_);
  or (_22663_, _22653_, _22160_);
  and (_22674_, _22663_, _22357_);
  nor (_22685_, _22357_, _21800_);
  nor (_22696_, _22685_, _22674_);
  and (_22707_, _22696_, _22642_);
  and (_22718_, _22095_, _21909_);
  nor (_22729_, _22718_, _22106_);
  not (_22740_, _22729_);
  and (_22751_, _22740_, _22357_);
  nor (_22762_, _22357_, _21866_);
  nor (_22773_, _22762_, _22751_);
  and (_22783_, _22773_, _21768_);
  nor (_22794_, _22773_, _21768_);
  nor (_22805_, _22794_, _22783_);
  not (_22816_, _22805_);
  nor (_22827_, _22073_, _22051_);
  nor (_22838_, _22827_, _22084_);
  not (_22849_, _22838_);
  and (_22860_, _22849_, _22357_);
  nor (_22871_, _22357_, _21964_);
  nor (_22882_, _22871_, _22860_);
  and (_22892_, _22882_, _21833_);
  not (_22903_, _22029_);
  and (_22914_, _22357_, _21986_);
  or (_22925_, _22914_, _22903_);
  nand (_22936_, _22357_, _21986_);
  or (_22947_, _22936_, _22029_);
  and (_22958_, _22947_, _22925_);
  nor (_22969_, _22958_, _21920_);
  and (_22990_, _22958_, _21920_);
  nor (_22991_, _22990_, _22969_);
  and (_23001_, _21227_, _19348_);
  nor (_23022_, _21227_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_23023_, _23022_, _23001_);
  nor (_23034_, _23023_, _21997_);
  not (_23055_, _23034_);
  and (_23056_, _23055_, _22991_);
  nor (_23067_, _23056_, _22969_);
  nor (_23088_, _22882_, _21833_);
  nor (_23089_, _23088_, _22892_);
  not (_23100_, _23089_);
  nor (_23120_, _23100_, _23067_);
  nor (_23121_, _23120_, _22892_);
  nor (_23132_, _23121_, _22816_);
  nor (_23153_, _23132_, _22783_);
  nor (_23154_, _22696_, _22642_);
  nor (_23165_, _23154_, _22707_);
  not (_23186_, _23165_);
  nor (_23187_, _23186_, _23153_);
  nor (_23198_, _23187_, _22707_);
  nor (_23209_, _23198_, _22631_);
  nor (_23219_, _23209_, _22620_);
  nor (_23230_, _23219_, _22544_);
  or (_23241_, _23230_, _22511_);
  or (_23252_, _23241_, _22435_);
  and (_23263_, _23252_, _22335_);
  nor (_23274_, _23263_, _22424_);
  and (_23285_, _22435_, _22335_);
  and (_23296_, _23285_, _23241_);
  or (_23307_, _23296_, _23274_);
  and (_00902_, _23307_, _41991_);
  or (_23328_, _22412_, _21217_);
  and (_23339_, _23328_, _23263_);
  and (_03002_, _23339_, _41991_);
  and (_03013_, _22357_, _41991_);
  and (_03034_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _41991_);
  and (_03056_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _41991_);
  and (_03077_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _41991_);
  or (_23400_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_23411_, _21055_, rst);
  and (_03088_, _23411_, _23400_);
  and (_23432_, _23339_, _21986_);
  or (_23443_, _23432_, _23023_);
  nand (_23454_, _23432_, _23023_);
  and (_23465_, _23454_, _23443_);
  and (_03099_, _23465_, _41991_);
  nor (_23486_, _23339_, _22958_);
  nor (_23497_, _23055_, _22991_);
  nor (_23508_, _23497_, _23056_);
  and (_23519_, _23508_, _23339_);
  or (_23530_, _23519_, _23486_);
  and (_03110_, _23530_, _41991_);
  and (_23551_, _23100_, _23067_);
  or (_23562_, _23551_, _23120_);
  nand (_23573_, _23562_, _23339_);
  or (_23584_, _23339_, _22882_);
  and (_23595_, _23584_, _23573_);
  and (_03121_, _23595_, _41991_);
  and (_23616_, _23121_, _22816_);
  or (_23627_, _23616_, _23132_);
  nand (_23638_, _23627_, _23339_);
  or (_23649_, _23339_, _22773_);
  and (_23660_, _23649_, _23638_);
  and (_03132_, _23660_, _41991_);
  and (_23681_, _23186_, _23153_);
  or (_23692_, _23681_, _23187_);
  nand (_23703_, _23692_, _23339_);
  or (_23714_, _23339_, _22696_);
  and (_23725_, _23714_, _23703_);
  and (_03143_, _23725_, _41991_);
  or (_23746_, _22631_, _22620_);
  and (_23757_, _23746_, _23198_);
  nor (_23768_, _23746_, _23198_);
  or (_23779_, _23768_, _23757_);
  nand (_23790_, _23779_, _23339_);
  or (_23801_, _23339_, _22609_);
  and (_23812_, _23801_, _23790_);
  and (_03154_, _23812_, _41991_);
  and (_23833_, _23219_, _22544_);
  or (_23844_, _23833_, _23230_);
  nand (_23855_, _23844_, _23339_);
  or (_23866_, _23339_, _22500_);
  and (_23877_, _23866_, _23855_);
  and (_03165_, _23877_, _41991_);
  not (_23898_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23909_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15624_);
  and (_23920_, _23909_, _23898_);
  and (_23931_, _23920_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23942_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23953_, _23942_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_23964_, _23942_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_23975_, _23964_, _23953_);
  and (_23986_, _23975_, _23931_);
  not (_23997_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_24008_, _23920_, _23997_);
  and (_24019_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24030_, _24019_, _23986_);
  not (_24041_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24052_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15624_);
  and (_24063_, _24052_, _24041_);
  and (_24074_, _24063_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24085_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24096_, _24063_, _23898_);
  and (_24107_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_24118_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24129_, _24118_, _15624_);
  nor (_24140_, _24129_, _24052_);
  and (_24151_, _24140_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24173_, _24151_, _24107_);
  nor (_24185_, _24173_, _24085_);
  and (_24197_, _24185_, _24030_);
  nor (_24209_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24221_, _24209_, _23942_);
  and (_24233_, _24221_, _23931_);
  and (_24245_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_24246_, _24245_, _24233_);
  and (_24257_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_24268_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_24279_, _24140_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_24290_, _24279_, _24268_);
  nor (_24301_, _24290_, _24257_);
  and (_24312_, _24301_, _24246_);
  and (_24323_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_24334_, _24140_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24345_, _24334_, _24323_);
  not (_24356_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24367_, _23931_, _24356_);
  not (_24378_, _24367_);
  and (_24389_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_24400_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_24411_, _24400_, _24389_);
  and (_24422_, _24411_, _24378_);
  and (_24433_, _24422_, _24345_);
  and (_24444_, _24433_, _24312_);
  and (_24455_, _24444_, _24197_);
  and (_24466_, _23953_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_24477_, _24466_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_24488_, _24477_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_24499_, _24488_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_24510_, _24499_);
  not (_24521_, _23931_);
  nor (_24532_, _24488_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_24543_, _24532_, _24521_);
  and (_24554_, _24543_, _24510_);
  not (_24565_, _24554_);
  and (_24576_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24587_, _24576_, _23909_);
  and (_24598_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_24610_, _24598_, _24587_);
  and (_24621_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_24632_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_24643_, _24632_, _24621_);
  and (_24654_, _24643_, _24610_);
  and (_24665_, _24654_, _24565_);
  nor (_24676_, _24477_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_24686_, _24676_);
  nor (_24697_, _24488_, _24521_);
  and (_24708_, _24697_, _24686_);
  not (_24719_, _24708_);
  and (_24730_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_24741_, _24730_, _24587_);
  and (_24752_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_24763_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_24774_, _24763_, _24752_);
  and (_24785_, _24774_, _24741_);
  and (_24795_, _24785_, _24719_);
  nor (_24806_, _24795_, _24665_);
  not (_24817_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_24828_, _24499_, _24817_);
  and (_24839_, _24499_, _24817_);
  nor (_24850_, _24839_, _24828_);
  nor (_24861_, _24850_, _24521_);
  not (_24872_, _24861_);
  and (_24883_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_24894_, _24883_, _24587_);
  and (_24905_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_24916_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_24927_, _24916_, _24905_);
  and (_24938_, _24927_, _24894_);
  and (_24949_, _24938_, _24872_);
  not (_24960_, _24949_);
  and (_24971_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_24982_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_24993_, _24982_, _24971_);
  not (_25004_, _24466_);
  nor (_25015_, _23953_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_25026_, _25015_, _24521_);
  and (_25036_, _25026_, _25004_);
  and (_25047_, _24140_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_25058_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_25069_, _25058_, _25047_);
  not (_25080_, _25069_);
  nor (_25101_, _25080_, _25036_);
  and (_25102_, _25101_, _24993_);
  not (_25113_, _25102_);
  and (_25124_, _24008_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_25145_, _25124_, _24587_);
  and (_25146_, _24074_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_25156_, _25146_);
  and (_25177_, _25156_, _25145_);
  nor (_25178_, _24466_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_25189_, _25178_);
  nor (_25200_, _24477_, _24521_);
  and (_25211_, _25200_, _25189_);
  and (_25232_, _24096_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_25233_, _24140_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_25244_, _25233_, _25232_);
  not (_25255_, _25244_);
  nor (_25265_, _25255_, _25211_);
  and (_25276_, _25265_, _25177_);
  nor (_25287_, _25276_, _25113_);
  and (_25298_, _25287_, _24960_);
  and (_25309_, _25298_, _24806_);
  nand (_25320_, _25309_, _24455_);
  and (_25331_, _23307_, _21044_);
  not (_25342_, _25331_);
  and (_25363_, _20439_, _15690_);
  not (_25364_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_25375_, _15635_, _25364_);
  and (_25385_, _25375_, _15679_);
  not (_25396_, _25385_);
  nor (_25407_, _17747_, _17573_);
  and (_25418_, _17747_, _17573_);
  nor (_25429_, _25418_, _25407_);
  not (_25440_, _16589_);
  nor (_25451_, _16907_, _25440_);
  nor (_25462_, _16907_, _16589_);
  and (_25473_, _16907_, _16589_);
  nor (_25484_, _25473_, _25462_);
  not (_25495_, _17235_);
  nor (_25506_, _17932_, _25495_);
  nor (_25517_, _17932_, _17235_);
  and (_25538_, _17932_, _17235_);
  nor (_25539_, _25538_, _25517_);
  not (_25550_, _16248_);
  and (_25561_, _18095_, _25550_);
  nor (_25571_, _25561_, _25539_);
  nor (_25582_, _25571_, _25506_);
  nor (_25593_, _25582_, _25484_);
  nor (_25604_, _25593_, _25451_);
  and (_25615_, _25582_, _25484_);
  nor (_25626_, _25615_, _25593_);
  not (_25637_, _25626_);
  and (_25647_, _25561_, _25539_);
  nor (_25658_, _25647_, _25571_);
  not (_25669_, _25658_);
  nor (_25680_, _18095_, _16248_);
  and (_25691_, _18095_, _16248_);
  nor (_25702_, _25691_, _25680_);
  not (_25713_, _25702_);
  and (_25733_, _18465_, _17083_);
  nor (_25734_, _18465_, _17083_);
  nor (_25745_, _25734_, _25733_);
  nor (_25756_, _18967_, _16084_);
  and (_25767_, _18967_, _16084_);
  nor (_25778_, _25767_, _25756_);
  nor (_25789_, _18803_, _17399_);
  and (_25800_, _18803_, _17399_);
  nor (_25811_, _25800_, _25789_);
  not (_25822_, _16413_);
  and (_25832_, _19348_, _25822_);
  nor (_25843_, _25832_, _25811_);
  not (_25854_, _17399_);
  nor (_25865_, _18803_, _25854_);
  nor (_25876_, _25865_, _25843_);
  nor (_25887_, _25876_, _25778_);
  not (_25898_, _16084_);
  nor (_25909_, _18967_, _25898_);
  nor (_25919_, _25909_, _25887_);
  nor (_25930_, _25919_, _25745_);
  and (_25941_, _25919_, _25745_);
  nor (_25952_, _25941_, _25930_);
  not (_25963_, _25952_);
  and (_25974_, _25876_, _25778_);
  nor (_25985_, _25974_, _25887_);
  not (_25996_, _25985_);
  and (_26006_, _25832_, _25811_);
  nor (_26017_, _26006_, _25843_);
  not (_26028_, _26017_);
  nor (_26039_, _19348_, _16413_);
  and (_26050_, _19348_, _16413_);
  nor (_26061_, _26050_, _26039_);
  not (_26082_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_26083_, _15897_, _26082_);
  not (_26093_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26104_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26115_, _26104_, _17464_);
  nor (_26126_, _26115_, _26093_);
  nor (_26137_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26148_, _26137_, _16139_);
  not (_26159_, _26148_);
  not (_26170_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26190_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _26170_);
  and (_26191_, _26190_, _17127_);
  not (_26202_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_26213_, _26202_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26224_, _26213_, _16479_);
  nor (_26235_, _26224_, _26191_);
  and (_26246_, _26235_, _26159_);
  and (_26256_, _26246_, _26126_);
  and (_26267_, _26104_, _16973_);
  nor (_26278_, _26267_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26289_, _26213_, _15941_);
  not (_26300_, _26289_);
  and (_26311_, _26190_, _17290_);
  and (_26322_, _26137_, _16303_);
  nor (_26333_, _26322_, _26311_);
  and (_26343_, _26333_, _26300_);
  and (_26354_, _26343_, _26278_);
  nor (_26365_, _26354_, _26256_);
  nor (_26376_, _26365_, _15897_);
  nor (_26387_, _26376_, _26083_);
  and (_26398_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_26409_, _26398_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_26420_, _26409_);
  and (_26431_, _26420_, _26387_);
  and (_26441_, _26420_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_26452_, _26441_, _26431_);
  nor (_26463_, _26452_, _26061_);
  and (_26474_, _26463_, _26028_);
  and (_26485_, _26474_, _25996_);
  and (_26496_, _26485_, _25963_);
  not (_26507_, _17083_);
  or (_26518_, _18465_, _26507_);
  and (_26528_, _18465_, _26507_);
  or (_26539_, _25919_, _26528_);
  and (_26550_, _26539_, _26518_);
  or (_26561_, _26550_, _26496_);
  and (_26572_, _26561_, _25713_);
  and (_26583_, _26572_, _25669_);
  and (_26594_, _26583_, _25637_);
  nor (_26605_, _26594_, _25604_);
  nor (_26615_, _26605_, _25429_);
  and (_26636_, _26605_, _25429_);
  nor (_26637_, _26636_, _26615_);
  nor (_26648_, _26637_, _25396_);
  not (_26659_, _26648_);
  not (_26670_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_26681_, _21001_, _26670_);
  and (_26692_, _26681_, _15679_);
  not (_26702_, _25484_);
  and (_26713_, _25680_, _25539_);
  nor (_26724_, _26713_, _25517_);
  nor (_26735_, _26724_, _26702_);
  not (_26746_, _25778_);
  and (_26757_, _26039_, _25811_);
  nor (_26768_, _26757_, _25789_);
  nor (_26779_, _26768_, _26746_);
  nor (_26789_, _26779_, _25756_);
  nor (_26800_, _26789_, _25745_);
  and (_26811_, _26789_, _25745_);
  nor (_26822_, _26811_, _26800_);
  not (_26833_, _26061_);
  nor (_26844_, _26452_, _26833_);
  and (_26855_, _26844_, _25811_);
  and (_26866_, _26768_, _26746_);
  nor (_26877_, _26866_, _26779_);
  and (_26888_, _26877_, _26855_);
  not (_26898_, _26888_);
  nor (_26909_, _26898_, _26822_);
  nor (_26930_, _26789_, _25733_);
  or (_26931_, _26930_, _25734_);
  or (_26942_, _26931_, _26909_);
  and (_26953_, _26942_, _25702_);
  and (_26964_, _26953_, _25539_);
  and (_26975_, _26724_, _26702_);
  nor (_26986_, _26975_, _26735_);
  and (_26997_, _26986_, _26964_);
  or (_27007_, _26997_, _26735_);
  nor (_27018_, _27007_, _25462_);
  and (_27039_, _27018_, _25429_);
  nor (_27040_, _27018_, _25429_);
  or (_27051_, _27040_, _27039_);
  and (_27062_, _27051_, _26692_);
  and (_27073_, _15668_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27084_, _27073_, _25375_);
  nor (_27095_, _19348_, _18803_);
  and (_27106_, _27095_, _18978_);
  and (_27117_, _27106_, _18476_);
  and (_27127_, _27117_, _18106_);
  and (_27138_, _27127_, _18509_);
  and (_27149_, _27138_, _16918_);
  and (_27160_, _27149_, _26452_);
  not (_27171_, _26452_);
  and (_27182_, _16907_, _17932_);
  and (_27193_, _19348_, _18803_);
  and (_27204_, _27193_, _18967_);
  and (_27215_, _27204_, _18465_);
  and (_27226_, _27215_, _18095_);
  and (_27236_, _27226_, _27182_);
  and (_27257_, _27236_, _27171_);
  nor (_27258_, _27257_, _27160_);
  and (_27269_, _27258_, _17747_);
  nor (_27280_, _27258_, _17747_);
  nor (_27291_, _27280_, _27269_);
  and (_27302_, _27291_, _27084_);
  not (_27313_, _17573_);
  nor (_27324_, _26452_, _27313_);
  not (_27335_, _27324_);
  and (_27346_, _26452_, _17747_);
  and (_27356_, _27073_, _15646_);
  not (_27367_, _27356_);
  nor (_27378_, _27367_, _27346_);
  and (_27389_, _27378_, _27335_);
  nor (_27400_, _27389_, _27302_);
  and (_27411_, _26681_, _21033_);
  not (_27422_, _27411_);
  and (_27433_, _18967_, _18803_);
  nor (_27444_, _27433_, _18465_);
  and (_27455_, _27444_, _27411_);
  and (_27466_, _27455_, _18106_);
  not (_27476_, _27466_);
  and (_27487_, _27476_, _27182_);
  nor (_27498_, _27182_, _17747_);
  nor (_27519_, _27498_, _27455_);
  and (_27520_, _27519_, _26452_);
  nor (_27531_, _27520_, _27487_);
  and (_27542_, _27531_, _17747_);
  nor (_27553_, _27531_, _17747_);
  nor (_27564_, _27553_, _27542_);
  nor (_27575_, _27564_, _27422_);
  not (_27585_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_27596_, _15668_, _27585_);
  and (_27607_, _27596_, _26681_);
  not (_27618_, _27607_);
  nor (_27629_, _27618_, _25418_);
  and (_27640_, _27596_, _21011_);
  and (_27651_, _27640_, _25429_);
  nor (_27662_, _27651_, _27629_);
  and (_27672_, _27073_, _21011_);
  not (_27683_, _27672_);
  nor (_27694_, _27683_, _19348_);
  and (_27705_, _27596_, _15635_);
  not (_27716_, _27705_);
  nor (_27727_, _27716_, _16907_);
  nor (_27738_, _27727_, _27694_);
  and (_27749_, _27073_, _26681_);
  not (_27760_, _27749_);
  nor (_27771_, _27760_, _26452_);
  and (_27782_, _21033_, _15646_);
  and (_27802_, _27782_, _25407_);
  and (_27803_, _25375_, _21033_);
  and (_27814_, _27803_, _17747_);
  nor (_27825_, _27814_, _27802_);
  and (_27836_, _21011_, _15679_);
  not (_27847_, _27836_);
  nor (_27858_, _27847_, _17747_);
  not (_27869_, _27858_);
  nand (_27880_, _27869_, _27825_);
  nor (_27891_, _27880_, _27771_);
  and (_27902_, _27891_, _27738_);
  and (_27913_, _27902_, _27662_);
  not (_27923_, _27913_);
  nor (_27934_, _27923_, _27575_);
  and (_27945_, _27934_, _27400_);
  not (_27956_, _27945_);
  nor (_27967_, _27956_, _27062_);
  and (_27978_, _27967_, _26659_);
  not (_27989_, _27978_);
  nor (_28000_, _27989_, _25363_);
  and (_28011_, _28000_, _25342_);
  not (_28022_, _28011_);
  or (_28033_, _28022_, _25320_);
  and (_28043_, \oc8051_top_1.oc8051_decoder1.wr , _15624_);
  not (_28054_, _28043_);
  nor (_28065_, _28054_, _23920_);
  not (_28076_, _28065_);
  nor (_28087_, _28076_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not (_28098_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_28109_, _25320_, _28098_);
  and (_28120_, _28109_, _28087_);
  and (_28131_, _28120_, _28033_);
  nor (_28142_, _28065_, _28098_);
  not (_28153_, _26692_);
  nor (_28164_, _27018_, _25418_);
  nor (_28175_, _28164_, _25407_);
  nor (_28185_, _28175_, _28153_);
  not (_28196_, _28185_);
  and (_28207_, _17747_, _27313_);
  nor (_28218_, _28207_, _26615_);
  nor (_28239_, _28218_, _25396_);
  nor (_28240_, _27466_, _18509_);
  and (_28251_, _26452_, _16907_);
  and (_28262_, _28251_, _28240_);
  nor (_28273_, _28262_, _27346_);
  nor (_28284_, _26452_, _17747_);
  not (_28295_, _28284_);
  nor (_28306_, _28295_, _27487_);
  nor (_28316_, _28306_, _27422_);
  and (_28327_, _28316_, _28273_);
  not (_28338_, _28327_);
  nor (_28349_, _27803_, _27171_);
  and (_28360_, _27683_, _26441_);
  nor (_28371_, _28360_, _26431_);
  nor (_28382_, _28371_, _27836_);
  nor (_28393_, _28382_, _28349_);
  not (_28404_, _28393_);
  nor (_28425_, _26441_, _26387_);
  not (_28426_, _27640_);
  nor (_28437_, _28426_, _26431_);
  nor (_28447_, _28437_, _27607_);
  nor (_28458_, _28447_, _28425_);
  not (_28469_, _28458_);
  and (_28480_, _26409_, _26387_);
  and (_28491_, _27596_, _25375_);
  and (_28502_, _27782_, _26387_);
  nor (_28513_, _28502_, _28491_);
  nor (_28524_, _28513_, _28480_);
  not (_28535_, _28524_);
  and (_28546_, _27596_, _15646_);
  not (_28556_, _28546_);
  nor (_28567_, _28556_, _17747_);
  not (_28578_, _28567_);
  nor (_28589_, _27760_, _19348_);
  nor (_28600_, _28589_, _27455_);
  and (_28611_, _28600_, _28578_);
  and (_28622_, _28611_, _28535_);
  and (_28633_, _28622_, _28469_);
  and (_28644_, _28633_, _28404_);
  and (_28655_, _28644_, _28338_);
  not (_28665_, _28655_);
  nor (_28676_, _28665_, _28239_);
  and (_28687_, _28676_, _28196_);
  not (_28698_, _24197_);
  nor (_28709_, _24433_, _24312_);
  and (_28720_, _28709_, _28698_);
  and (_28731_, _28720_, _25309_);
  nand (_28742_, _28731_, _28687_);
  and (_28753_, _28065_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_28764_, _28731_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_28775_, _28764_, _28753_);
  and (_28785_, _28775_, _28742_);
  or (_28796_, _28785_, _28142_);
  or (_28807_, _28796_, _28131_);
  and (_06683_, _28807_, _41991_);
  and (_28828_, _23465_, _21044_);
  not (_28839_, _28828_);
  and (_28850_, _20768_, _15690_);
  and (_28861_, _26452_, _26833_);
  nor (_28872_, _28861_, _26844_);
  nor (_28883_, _26692_, _25385_);
  not (_28893_, _28883_);
  and (_28904_, _28893_, _28872_);
  not (_28915_, _28904_);
  nor (_28926_, _28556_, _26452_);
  not (_28937_, _28926_);
  nor (_28958_, _28426_, _26039_);
  nor (_28959_, _28958_, _27607_);
  or (_28970_, _28959_, _26050_);
  and (_28981_, _28491_, _18204_);
  and (_28992_, _27073_, _26670_);
  not (_29003_, _28992_);
  nor (_29013_, _29003_, _18803_);
  nor (_29024_, _29013_, _28981_);
  and (_29035_, _27782_, _26039_);
  and (_29046_, _27803_, _19348_);
  nor (_29057_, _29046_, _29035_);
  nor (_29068_, _27367_, _16413_);
  and (_29079_, _27084_, _19348_);
  nor (_29090_, _29079_, _29068_);
  nor (_29101_, _27836_, _27411_);
  nor (_29112_, _29101_, _19348_);
  not (_29122_, _29112_);
  and (_29133_, _29122_, _29090_);
  and (_29144_, _29133_, _29057_);
  and (_29155_, _29144_, _29024_);
  and (_29166_, _29155_, _28970_);
  and (_29177_, _29166_, _28937_);
  and (_29188_, _29177_, _28915_);
  not (_29199_, _29188_);
  nor (_29210_, _29199_, _28850_);
  and (_29221_, _29210_, _28839_);
  not (_29232_, _29221_);
  or (_29242_, _29232_, _25320_);
  not (_29253_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_29264_, _25320_, _29253_);
  and (_29275_, _29264_, _28087_);
  and (_29286_, _29275_, _29242_);
  nor (_29297_, _28065_, _29253_);
  not (_29308_, _28687_);
  or (_29319_, _29308_, _25320_);
  and (_29329_, _29264_, _28753_);
  and (_29340_, _29329_, _29319_);
  or (_29351_, _29340_, _29297_);
  or (_29362_, _29351_, _29286_);
  and (_08921_, _29362_, _41991_);
  and (_29383_, _23530_, _21044_);
  not (_29394_, _29383_);
  and (_29405_, _20799_, _15690_);
  nor (_29415_, _26039_, _25811_);
  or (_29426_, _29415_, _26757_);
  and (_29437_, _29426_, _26844_);
  nor (_29448_, _29426_, _26844_);
  or (_29459_, _29448_, _29437_);
  and (_29470_, _29459_, _26692_);
  nor (_29481_, _26463_, _26028_);
  nor (_29501_, _29481_, _26474_);
  nor (_29502_, _29501_, _25396_);
  nor (_29513_, _29502_, _29470_);
  nor (_29524_, _27367_, _17399_);
  nor (_29535_, _27193_, _27095_);
  not (_29546_, _29535_);
  nor (_29557_, _29546_, _26452_);
  and (_29568_, _29546_, _26452_);
  nor (_29579_, _29568_, _29557_);
  and (_29589_, _29579_, _27084_);
  nor (_29600_, _29589_, _29524_);
  nor (_29611_, _27444_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_29622_, _29611_, _19011_);
  nor (_29633_, _29611_, _19011_);
  nor (_29644_, _29633_, _29622_);
  nor (_29655_, _29644_, _27422_);
  not (_29666_, _29655_);
  and (_29676_, _27640_, _25811_);
  nor (_29687_, _27618_, _25800_);
  not (_29698_, _29687_);
  and (_29709_, _27782_, _25789_);
  and (_29720_, _27803_, _18803_);
  nor (_29731_, _29720_, _29709_);
  nand (_29742_, _29731_, _29698_);
  nor (_29762_, _29742_, _29676_);
  nor (_29763_, _27847_, _18803_);
  not (_29774_, _29763_);
  nor (_29785_, _29003_, _18967_);
  nor (_29796_, _27716_, _19348_);
  nor (_29807_, _29796_, _29785_);
  and (_29818_, _29807_, _29774_);
  and (_29829_, _29818_, _29762_);
  and (_29840_, _29829_, _29666_);
  and (_29850_, _29840_, _29600_);
  and (_29861_, _29850_, _29513_);
  not (_29872_, _29861_);
  nor (_29883_, _29872_, _29405_);
  and (_29894_, _29883_, _29394_);
  not (_29905_, _29894_);
  or (_29916_, _29905_, _25320_);
  not (_29926_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_29937_, _25320_, _29926_);
  and (_29948_, _29937_, _28087_);
  and (_29959_, _29948_, _29916_);
  nor (_29970_, _28065_, _29926_);
  not (_29981_, _24433_);
  and (_29992_, _29981_, _24312_);
  and (_30003_, _29992_, _24197_);
  and (_30013_, _30003_, _25309_);
  or (_30024_, _30013_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_30035_, _30024_, _28753_);
  nand (_30046_, _30013_, _28687_);
  and (_30067_, _30046_, _30035_);
  or (_30068_, _30067_, _29970_);
  or (_30079_, _30068_, _29959_);
  and (_08932_, _30079_, _41991_);
  and (_30099_, _20831_, _15690_);
  not (_30110_, _30099_);
  and (_30121_, _23595_, _21044_);
  nor (_30132_, _27367_, _16084_);
  and (_30143_, _27193_, _27171_);
  and (_30154_, _27095_, _26452_);
  nor (_30165_, _30154_, _30143_);
  nor (_30176_, _30165_, _18967_);
  not (_30186_, _27084_);
  and (_30197_, _30165_, _18967_);
  or (_30208_, _30197_, _30186_);
  nor (_30219_, _30208_, _30176_);
  nor (_30230_, _30219_, _30132_);
  nor (_30241_, _26474_, _25996_);
  nor (_30252_, _30241_, _26485_);
  nor (_30263_, _30252_, _25396_);
  not (_30274_, _30263_);
  nor (_30284_, _29003_, _18465_);
  and (_30295_, _27782_, _25756_);
  and (_30306_, _27803_, _18967_);
  nor (_30317_, _30306_, _30295_);
  nor (_30328_, _27618_, _25767_);
  and (_30339_, _27640_, _25778_);
  nor (_30350_, _30339_, _30328_);
  nor (_30361_, _27716_, _18803_);
  nor (_30371_, _27847_, _18967_);
  nor (_30392_, _30371_, _30361_);
  and (_30393_, _30392_, _30350_);
  nand (_30404_, _30393_, _30317_);
  nor (_30415_, _30404_, _30284_);
  and (_30426_, _30415_, _30274_);
  nor (_30437_, _26877_, _26855_);
  nor (_30448_, _30437_, _28153_);
  and (_30459_, _30448_, _26898_);
  and (_30480_, _27433_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30491_, _29633_, _18967_);
  nor (_30502_, _30491_, _30480_);
  nor (_30513_, _30502_, _27422_);
  nor (_30524_, _30513_, _30459_);
  and (_30535_, _30524_, _30426_);
  and (_30546_, _30535_, _30230_);
  not (_30556_, _30546_);
  nor (_30567_, _30556_, _30121_);
  and (_30578_, _30567_, _30110_);
  not (_30589_, _30578_);
  or (_30600_, _30589_, _25320_);
  not (_30611_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_30622_, _25320_, _30611_);
  and (_30633_, _30622_, _28087_);
  and (_30643_, _30633_, _30600_);
  nor (_30654_, _28065_, _30611_);
  nand (_30665_, _25309_, _24197_);
  or (_30676_, _28709_, _30665_);
  and (_30687_, _30676_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_30698_, _24312_);
  and (_30709_, _24197_, _24433_);
  and (_30720_, _30709_, _30698_);
  and (_30730_, _30720_, _29308_);
  and (_30741_, _24197_, _24312_);
  and (_30752_, _30741_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_30763_, _30752_, _30730_);
  and (_30774_, _30763_, _25309_);
  or (_30785_, _30774_, _30687_);
  and (_30796_, _30785_, _28753_);
  or (_30807_, _30796_, _30654_);
  or (_30817_, _30807_, _30643_);
  and (_08943_, _30817_, _41991_);
  and (_30838_, _20874_, _15690_);
  not (_30849_, _30838_);
  and (_30860_, _23660_, _21044_);
  nor (_30881_, _26485_, _25963_);
  nor (_30882_, _30881_, _26496_);
  nor (_30893_, _30882_, _25396_);
  not (_30903_, _30893_);
  and (_30914_, _27640_, _25745_);
  nor (_30925_, _27618_, _25733_);
  or (_30936_, _30925_, _30914_);
  not (_30947_, _30936_);
  and (_30958_, _26898_, _26822_);
  or (_30969_, _30958_, _28153_);
  nor (_30980_, _30969_, _26909_);
  nor (_30990_, _27367_, _17083_);
  and (_31001_, _27106_, _26452_);
  and (_31012_, _27204_, _27171_);
  nor (_31023_, _31012_, _31001_);
  nor (_31034_, _31023_, _18465_);
  and (_31045_, _31023_, _18465_);
  or (_31056_, _31045_, _30186_);
  nor (_31067_, _31056_, _31034_);
  nor (_31077_, _31067_, _30990_);
  nor (_31088_, _27716_, _18967_);
  nor (_31109_, _27847_, _18465_);
  nor (_31110_, _31109_, _31088_);
  not (_31121_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_31132_, _27433_, _31121_);
  nor (_31143_, _31132_, _18476_);
  or (_31153_, _31143_, _27422_);
  or (_31164_, _31153_, _27444_);
  nor (_31175_, _29003_, _18095_);
  not (_31186_, _31175_);
  and (_31197_, _27782_, _25734_);
  and (_31208_, _27803_, _18465_);
  nor (_31219_, _31208_, _31197_);
  and (_31230_, _31219_, _31186_);
  and (_31240_, _31230_, _31164_);
  and (_31251_, _31240_, _31110_);
  nand (_31262_, _31251_, _31077_);
  nor (_31273_, _31262_, _30980_);
  and (_31284_, _31273_, _30947_);
  and (_31295_, _31284_, _30903_);
  not (_31306_, _31295_);
  nor (_31317_, _31306_, _30860_);
  and (_31327_, _31317_, _30849_);
  not (_31338_, _31327_);
  or (_31349_, _31338_, _25320_);
  not (_31360_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_31371_, _25320_, _31360_);
  and (_31382_, _31371_, _28087_);
  and (_31393_, _31382_, _31349_);
  nor (_31404_, _28065_, _31360_);
  and (_31414_, _30665_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_31425_, _28709_, _24197_);
  not (_31436_, _31425_);
  nor (_31447_, _31436_, _28687_);
  nor (_31458_, _30741_, _30709_);
  nor (_31469_, _31458_, _31360_);
  or (_31480_, _31469_, _31447_);
  and (_31491_, _31480_, _25309_);
  or (_31502_, _31491_, _31414_);
  and (_31512_, _31502_, _28753_);
  or (_31523_, _31512_, _31404_);
  or (_31534_, _31523_, _31393_);
  and (_08954_, _31534_, _41991_);
  and (_31555_, _23725_, _21044_);
  not (_31566_, _31555_);
  and (_31577_, _20905_, _15690_);
  or (_31588_, _26942_, _25702_);
  nor (_31598_, _28153_, _26953_);
  and (_31609_, _31598_, _31588_);
  nor (_31620_, _26561_, _25702_);
  and (_31631_, _26561_, _25702_);
  nor (_31642_, _31631_, _31620_);
  and (_31653_, _31642_, _25385_);
  or (_31664_, _27455_, _18106_);
  and (_31684_, _31664_, _27411_);
  and (_31685_, _31684_, _27476_);
  and (_31696_, _27117_, _26452_);
  and (_31707_, _27215_, _27171_);
  nor (_31718_, _31707_, _31696_);
  and (_31729_, _31718_, _18095_);
  nor (_31740_, _31718_, _18095_);
  nor (_31751_, _31740_, _31729_);
  and (_31761_, _31751_, _27084_);
  nor (_31772_, _26452_, _16248_);
  and (_31783_, _26452_, _18106_);
  nor (_31794_, _31783_, _31772_);
  nor (_31805_, _31794_, _27367_);
  nor (_31816_, _31805_, _31761_);
  and (_31827_, _27782_, _25680_);
  and (_31838_, _27803_, _18095_);
  nor (_31848_, _31838_, _31827_);
  or (_31859_, _29003_, _17932_);
  nand (_31870_, _31859_, _31848_);
  and (_31881_, _27640_, _25702_);
  nor (_31892_, _27618_, _25691_);
  or (_31903_, _31892_, _31881_);
  nor (_31914_, _27847_, _18095_);
  nor (_31925_, _27716_, _18465_);
  or (_31935_, _31925_, _31914_);
  or (_31946_, _31935_, _31903_);
  nor (_31957_, _31946_, _31870_);
  nand (_31968_, _31957_, _31816_);
  or (_31979_, _31968_, _31685_);
  or (_31990_, _31979_, _31653_);
  or (_32001_, _31990_, _31609_);
  nor (_32012_, _32001_, _31577_);
  and (_32022_, _32012_, _31566_);
  not (_32033_, _32022_);
  or (_32044_, _32033_, _25320_);
  not (_32055_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_32066_, _25320_, _32055_);
  and (_32077_, _32066_, _28087_);
  and (_32088_, _32077_, _32044_);
  nor (_32099_, _28065_, _32055_);
  not (_32109_, _25309_);
  and (_32120_, _24444_, _28698_);
  nor (_32131_, _24444_, _28698_);
  nor (_32142_, _32131_, _32120_);
  or (_32153_, _32142_, _32109_);
  and (_32164_, _32153_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_32175_, _32120_, _29308_);
  and (_32186_, _32131_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_32196_, _32186_, _32175_);
  and (_32207_, _32196_, _25309_);
  or (_32218_, _32207_, _32164_);
  and (_32229_, _32218_, _28753_);
  or (_32240_, _32229_, _32099_);
  or (_32251_, _32240_, _32088_);
  and (_08964_, _32251_, _41991_);
  and (_32272_, _23812_, _21044_);
  not (_32282_, _32272_);
  and (_32293_, _20948_, _15690_);
  nor (_32314_, _25680_, _25539_);
  nor (_32315_, _32314_, _26713_);
  nor (_32326_, _32315_, _26953_);
  nor (_32337_, _32326_, _26964_);
  and (_32348_, _32337_, _26692_);
  not (_32359_, _32348_);
  nor (_32370_, _26572_, _25669_);
  nor (_32381_, _32370_, _26583_);
  nor (_32392_, _32381_, _25396_);
  nor (_32403_, _26452_, _17235_);
  and (_32414_, _26452_, _18509_);
  nor (_32425_, _32414_, _32403_);
  nor (_32436_, _32425_, _27367_);
  and (_32447_, _27127_, _26452_);
  and (_32458_, _27226_, _27171_);
  nor (_32469_, _32458_, _32447_);
  and (_32480_, _32469_, _17932_);
  nor (_32491_, _32469_, _17932_);
  or (_32502_, _32491_, _30186_);
  nor (_32513_, _32502_, _32480_);
  nor (_32524_, _32513_, _32436_);
  not (_32535_, _27520_);
  and (_32545_, _32535_, _28240_);
  nor (_32556_, _27520_, _27466_);
  nor (_32567_, _32556_, _17932_);
  nor (_32578_, _32567_, _32545_);
  nor (_32589_, _32578_, _27422_);
  and (_32600_, _27640_, _25539_);
  and (_32621_, _27782_, _25517_);
  nor (_32622_, _27618_, _25538_);
  and (_32633_, _27803_, _17932_);
  or (_32644_, _32633_, _32622_);
  or (_32655_, _32644_, _32621_);
  nor (_32666_, _32655_, _32600_);
  nor (_32677_, _29003_, _16907_);
  not (_32688_, _32677_);
  nor (_32699_, _27847_, _17932_);
  nor (_32710_, _27716_, _18095_);
  nor (_32721_, _32710_, _32699_);
  and (_32732_, _32721_, _32688_);
  and (_32743_, _32732_, _32666_);
  not (_32754_, _32743_);
  nor (_32765_, _32754_, _32589_);
  and (_32776_, _32765_, _32524_);
  not (_32787_, _32776_);
  nor (_32798_, _32787_, _32392_);
  and (_32809_, _32798_, _32359_);
  not (_32820_, _32809_);
  nor (_32831_, _32820_, _32293_);
  and (_32842_, _32831_, _32282_);
  not (_32853_, _32842_);
  or (_32864_, _32853_, _25320_);
  not (_32875_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_32886_, _25320_, _32875_);
  and (_32897_, _32886_, _28087_);
  and (_32908_, _32897_, _32864_);
  nor (_32919_, _28065_, _32875_);
  and (_32930_, _29992_, _28698_);
  and (_32940_, _32930_, _25309_);
  nand (_32951_, _32940_, _28687_);
  or (_32972_, _32940_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_32973_, _32972_, _28753_);
  and (_32984_, _32973_, _32951_);
  or (_32995_, _32984_, _32919_);
  or (_33006_, _32995_, _32908_);
  and (_08975_, _33006_, _41991_);
  and (_33027_, _23877_, _21044_);
  not (_33038_, _33027_);
  and (_33049_, _20980_, _15690_);
  nor (_33060_, _26986_, _26964_);
  not (_33071_, _33060_);
  nor (_33082_, _28153_, _26997_);
  and (_33093_, _33082_, _33071_);
  not (_33104_, _33093_);
  nor (_33115_, _26583_, _25637_);
  nor (_33126_, _33115_, _26594_);
  nor (_33137_, _33126_, _25396_);
  nor (_33148_, _26452_, _25440_);
  or (_33159_, _33148_, _27367_);
  nor (_33170_, _33159_, _28251_);
  or (_33181_, _26452_, _17932_);
  or (_33192_, _32458_, _27138_);
  and (_33203_, _33192_, _33181_);
  nor (_33214_, _33203_, _16918_);
  and (_33225_, _33203_, _16918_);
  or (_33236_, _33225_, _30186_);
  nor (_33247_, _33236_, _33214_);
  nor (_33258_, _33247_, _33170_);
  nor (_33269_, _32545_, _16907_);
  and (_33280_, _32545_, _16907_);
  nor (_33291_, _33280_, _33269_);
  nor (_33301_, _33291_, _27422_);
  nor (_33312_, _27618_, _25473_);
  and (_33323_, _27640_, _25484_);
  nor (_33344_, _33323_, _33312_);
  and (_33345_, _27782_, _25462_);
  and (_33356_, _27803_, _16907_);
  nor (_33367_, _33356_, _33345_);
  nor (_33378_, _29003_, _17747_);
  not (_33389_, _33378_);
  nor (_33400_, _27847_, _16907_);
  nor (_33411_, _27716_, _17932_);
  nor (_33422_, _33411_, _33400_);
  and (_33433_, _33422_, _33389_);
  and (_33444_, _33433_, _33367_);
  and (_33455_, _33444_, _33344_);
  not (_33466_, _33455_);
  nor (_33477_, _33466_, _33301_);
  and (_33488_, _33477_, _33258_);
  not (_33499_, _33488_);
  nor (_33510_, _33499_, _33137_);
  and (_33521_, _33510_, _33104_);
  not (_33532_, _33521_);
  nor (_33543_, _33532_, _33049_);
  and (_33554_, _33543_, _33038_);
  not (_33565_, _33554_);
  or (_33576_, _33565_, _25320_);
  not (_33587_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_33598_, _25320_, _33587_);
  and (_33609_, _33598_, _28087_);
  and (_33620_, _33609_, _33576_);
  nor (_33631_, _28065_, _33587_);
  nor (_33642_, _24197_, _24312_);
  and (_33652_, _33642_, _24433_);
  and (_33663_, _33652_, _25309_);
  nand (_33674_, _33663_, _28687_);
  or (_33685_, _33663_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_33696_, _33685_, _28753_);
  and (_33707_, _33696_, _33674_);
  or (_33718_, _33707_, _33631_);
  or (_33729_, _33718_, _33620_);
  and (_08986_, _33729_, _41991_);
  and (_33750_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33761_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_33772_, _15624_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_33783_, _33772_, _33761_);
  not (_33794_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_33805_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_33816_, _33805_, _33794_);
  nor (_33827_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_33838_, _33827_, _15624_);
  and (_33849_, _33838_, _33816_);
  not (_33870_, _33849_);
  and (_33871_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not (_33882_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_33893_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_33904_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_33915_, _33904_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_33926_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33937_, _33926_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_33948_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  not (_33959_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_33970_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_33981_, _33970_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33992_, _33981_, _33959_);
  and (_34002_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_34013_, _34002_, _33948_);
  and (_34024_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34035_, _34024_, _33959_);
  and (_34046_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not (_34057_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_34068_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _34057_);
  and (_34079_, _34068_, _33959_);
  and (_34090_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34101_, _34090_, _34046_);
  and (_34112_, _34101_, _34013_);
  nor (_34123_, _33926_, _33959_);
  and (_34144_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_34145_, _33926_, _33959_);
  and (_34156_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_34167_, _34156_, _34144_);
  and (_34178_, _34167_, _34112_);
  nor (_34189_, _34178_, _33915_);
  or (_34200_, _34189_, _33893_);
  and (_34211_, _34200_, _33882_);
  nor (_34222_, _34211_, _33871_);
  nor (_34233_, _34222_, _33870_);
  and (_34244_, _33816_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_34255_, _34244_, _33870_);
  nor (_34266_, _34255_, _34233_);
  not (_34277_, _34266_);
  and (_34288_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34299_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34310_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_34321_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_34332_, _34321_, _34310_);
  and (_34343_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_34353_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_34364_, _34353_, _34343_);
  and (_34375_, _34364_, _34332_);
  and (_34386_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34397_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_34408_, _34397_, _34386_);
  and (_34419_, _34408_, _34375_);
  nor (_34430_, _34419_, _33915_);
  nor (_34441_, _34430_, _34299_);
  nor (_34452_, _34441_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34463_, _34452_, _34288_);
  nor (_34474_, _34463_, _33870_);
  and (_34485_, _33816_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_34496_, _34485_, _33870_);
  nor (_34507_, _34496_, _34474_);
  nor (_34518_, _34507_, _34277_);
  and (_34529_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34540_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_34551_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34562_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_34573_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_34584_, _34573_, _34562_);
  and (_34595_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_34606_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_34617_, _34606_, _34595_);
  and (_34628_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_34639_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_34650_, _34639_, _34628_);
  and (_34661_, _34650_, _34617_);
  and (_34672_, _34661_, _34584_);
  nor (_34683_, _34672_, _33904_);
  and (_34694_, _34683_, _34551_);
  or (_34704_, _34694_, _34540_);
  and (_34715_, _34704_, _33882_);
  nor (_34726_, _34715_, _34529_);
  nor (_34737_, _34726_, _33870_);
  and (_34748_, _33816_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_34769_, _34748_, _33870_);
  nor (_34770_, _34769_, _34737_);
  and (_34781_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_34792_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_34803_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_34814_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_34825_, _34814_, _34803_);
  and (_34836_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_34847_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_34858_, _34847_, _34836_);
  and (_34869_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_34880_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_34891_, _34880_, _34869_);
  and (_34902_, _34891_, _34858_);
  and (_34913_, _34902_, _34825_);
  nor (_34924_, _34913_, _33915_);
  nor (_34935_, _34924_, _34792_);
  nor (_34946_, _34935_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_34957_, _34946_, _34781_);
  nor (_34968_, _34957_, _33870_);
  and (_34979_, _33816_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_34990_, _34979_, _33870_);
  nor (_35001_, _34990_, _34968_);
  and (_35012_, _35001_, _34770_);
  and (_35023_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_35034_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_35045_, _35034_, _35023_);
  and (_35055_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not (_35066_, _35055_);
  and (_35077_, _35066_, _35045_);
  and (_35088_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_35099_, _35088_, _33904_);
  and (_35110_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_35121_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_35132_, _35121_, _35110_);
  and (_35143_, _35132_, _35099_);
  and (_35154_, _35143_, _35077_);
  and (_35165_, _35154_, _34551_);
  nor (_35176_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _34551_);
  or (_35187_, _35176_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35198_, _35187_, _35165_);
  and (_35209_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_35220_, _35209_, _35198_);
  and (_35231_, _35220_, _33849_);
  and (_35242_, _33816_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_35253_, _35242_, _33870_);
  nor (_35264_, _35253_, _35231_);
  and (_35275_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35286_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35297_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_35308_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_35319_, _35308_, _35297_);
  and (_35330_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_35341_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_35352_, _35341_, _35330_);
  and (_35363_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_35373_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_35384_, _35373_, _35363_);
  and (_35395_, _35384_, _35352_);
  and (_35406_, _35395_, _35319_);
  nor (_35417_, _35406_, _33904_);
  and (_35428_, _35417_, _34551_);
  or (_35439_, _35428_, _35286_);
  and (_35450_, _35439_, _33882_);
  nor (_35461_, _35450_, _35275_);
  nor (_35483_, _35461_, _33870_);
  and (_35484_, _33816_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_35506_, _35484_, _33870_);
  nor (_35507_, _35506_, _35483_);
  and (_35529_, _35507_, _35264_);
  and (_35530_, _35529_, _35012_);
  and (_35552_, _35530_, _34518_);
  and (_35553_, _35552_, _33783_);
  nor (_35564_, _33827_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_35575_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_35586_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_35597_, _35586_, _35575_);
  and (_35608_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_35619_, _35608_, _33904_);
  and (_35630_, _35619_, _35597_);
  and (_35641_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_35652_, _35641_);
  and (_35663_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_35674_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_35685_, _35674_, _35663_);
  and (_35696_, _35685_, _35652_);
  and (_35706_, _35696_, _35630_);
  and (_35717_, _35706_, _34551_);
  nor (_35728_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _34551_);
  nor (_35739_, _35728_, _35717_);
  nor (_35750_, _35739_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_35761_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _33882_);
  nor (_35772_, _35761_, _35750_);
  and (_35783_, _35772_, _33849_);
  and (_35794_, _33816_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_35805_, _35794_, _33870_);
  nor (_35816_, _35805_, _35783_);
  and (_35827_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_35838_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_35849_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_35860_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_35871_, _35860_, _35849_);
  and (_35882_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_35893_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_35904_, _35893_, _35882_);
  and (_35915_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_35926_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_35937_, _35926_, _35915_);
  and (_35948_, _35937_, _35904_);
  and (_35959_, _35948_, _35871_);
  nor (_35970_, _35959_, _33904_);
  and (_35981_, _35970_, _34551_);
  or (_35992_, _35981_, _35838_);
  and (_36003_, _35992_, _33882_);
  nor (_36013_, _36003_, _35827_);
  nor (_36024_, _36013_, _33870_);
  and (_36035_, _33816_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_36046_, _36035_, _33870_);
  nor (_36057_, _36046_, _36024_);
  not (_36068_, _36057_);
  and (_36079_, _34507_, _34277_);
  and (_36090_, _36079_, _36068_);
  and (_36101_, _36090_, _35816_);
  not (_36112_, _35507_);
  not (_36123_, _35264_);
  and (_36134_, _35012_, _36123_);
  and (_36145_, _36134_, _36112_);
  and (_36156_, _36145_, _36101_);
  not (_36167_, _35816_);
  and (_36178_, _34507_, _36057_);
  and (_36189_, _36178_, _34277_);
  and (_36200_, _36189_, _36167_);
  and (_36211_, _36145_, _36200_);
  nor (_36222_, _34507_, _36057_);
  and (_36233_, _36222_, _34266_);
  and (_36244_, _36233_, _36167_);
  and (_36255_, _36145_, _36244_);
  nor (_36266_, _36255_, _36211_);
  not (_36277_, _36266_);
  nor (_36288_, _36277_, _36156_);
  and (_36299_, _36189_, _35816_);
  not (_36310_, _35001_);
  and (_36320_, _36310_, _34770_);
  and (_36331_, _35529_, _36320_);
  and (_36342_, _36331_, _36299_);
  and (_36353_, _36331_, _36101_);
  nor (_36364_, _36353_, _36342_);
  and (_36375_, _36364_, _36288_);
  nor (_36386_, _36375_, _35564_);
  or (_36397_, _36386_, _35553_);
  not (_36408_, _35564_);
  nor (_36419_, _36364_, _36408_);
  nor (_36430_, _36419_, _36397_);
  nor (_36441_, _36430_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36452_, _36441_, _33750_);
  and (_36463_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36474_, _35507_, _36123_);
  and (_36485_, _36474_, _36320_);
  and (_36496_, _36222_, _34277_);
  and (_36507_, _36496_, _35816_);
  and (_36518_, _36507_, _36485_);
  not (_36529_, _36518_);
  nor (_36540_, _35264_, _35001_);
  and (_36551_, _36540_, _34770_);
  and (_36562_, _36551_, _35816_);
  and (_36573_, _36562_, _36090_);
  and (_36584_, _36079_, _36167_);
  and (_36595_, _36584_, _36485_);
  nor (_36606_, _36595_, _36573_);
  and (_36616_, _36606_, _36529_);
  and (_36627_, _36134_, _35507_);
  and (_36638_, _36627_, _36200_);
  and (_36649_, _36299_, _36485_);
  nor (_36660_, _36649_, _36638_);
  and (_36671_, _34507_, _34266_);
  and (_36682_, _36671_, _36068_);
  and (_36693_, _36682_, _36627_);
  not (_36704_, _36693_);
  not (_36715_, _34770_);
  and (_36726_, _35816_, _36715_);
  and (_36737_, _36726_, _36090_);
  and (_36748_, _36671_, _36057_);
  and (_36759_, _36748_, _35816_);
  and (_36770_, _36759_, _36485_);
  nor (_36781_, _36770_, _36737_);
  and (_36792_, _36781_, _36704_);
  and (_36803_, _36792_, _36660_);
  and (_36814_, _36299_, _36627_);
  and (_36825_, _36057_, _36167_);
  and (_36836_, _34518_, _36825_);
  and (_36847_, _36836_, _36134_);
  nor (_36858_, _36847_, _36814_);
  and (_36869_, _35530_, _36682_);
  and (_36880_, _36869_, _35816_);
  and (_36891_, _36682_, _36167_);
  and (_36902_, _36671_, _36825_);
  or (_36913_, _36902_, _36891_);
  and (_36923_, _36913_, _35530_);
  nor (_36934_, _36923_, _36880_);
  and (_36945_, _36934_, _36858_);
  and (_36956_, _36945_, _36803_);
  and (_36967_, _36956_, _36616_);
  nor (_36978_, _34507_, _36068_);
  and (_36989_, _36978_, _34266_);
  and (_37000_, _36989_, _35816_);
  and (_37011_, _37000_, _36134_);
  not (_37022_, _37011_);
  and (_37033_, _36902_, _36485_);
  and (_37044_, _36090_, _36167_);
  and (_37055_, _35530_, _37044_);
  nor (_37066_, _37055_, _37033_);
  and (_37077_, _37066_, _37022_);
  and (_37088_, _36244_, _36627_);
  and (_37099_, _36978_, _34277_);
  and (_37110_, _37099_, _36167_);
  and (_37121_, _37110_, _36485_);
  nor (_37132_, _37121_, _37088_);
  and (_37143_, _37132_, _37077_);
  and (_37154_, _35530_, _36101_);
  and (_37165_, _37000_, _36485_);
  nor (_37176_, _37165_, _37154_);
  and (_37187_, _36627_, _37044_);
  and (_37198_, _37099_, _35816_);
  and (_37209_, _37198_, _36627_);
  nor (_37220_, _37209_, _37187_);
  and (_37229_, _37220_, _37176_);
  and (_37237_, _37229_, _37143_);
  not (_37245_, _36485_);
  nor (_37252_, _36836_, _36682_);
  nor (_37260_, _37252_, _37245_);
  and (_37268_, _37099_, _35530_);
  and (_37275_, _36233_, _35816_);
  and (_37283_, _37275_, _36134_);
  nor (_37291_, _37283_, _37268_);
  not (_37292_, _37291_);
  nor (_37293_, _37292_, _37260_);
  and (_37295_, _37275_, _36485_);
  and (_37306_, _37198_, _36485_);
  nor (_37317_, _37306_, _37295_);
  and (_37328_, _36101_, _36627_);
  and (_37339_, _37110_, _36627_);
  nor (_37350_, _37339_, _37328_);
  and (_37361_, _37350_, _37317_);
  and (_37372_, _37361_, _37293_);
  and (_37383_, _37372_, _37237_);
  and (_37394_, _37383_, _36967_);
  nor (_37405_, _37394_, _35564_);
  and (_37416_, _33772_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37427_, _37416_, _36693_);
  not (_37438_, _37427_);
  and (_37449_, _36682_, _35816_);
  and (_37460_, _37449_, _35530_);
  and (_37471_, _36902_, _35530_);
  nor (_37482_, _37471_, _37460_);
  not (_37493_, _33783_);
  nor (_37504_, _37493_, _37482_);
  nor (_37515_, _37504_, _35553_);
  and (_37526_, _37515_, _37438_);
  not (_37536_, _37526_);
  nor (_37547_, _37536_, _37405_);
  nor (_37558_, _37547_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37563_, _37558_, _36463_);
  and (_37573_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_37584_, _36167_, _34770_);
  and (_37595_, _37584_, _36540_);
  and (_37605_, _37595_, _36989_);
  and (_37616_, _36682_, _36551_);
  or (_37627_, _37616_, _37605_);
  not (_37637_, _37627_);
  and (_37648_, _36748_, _36551_);
  and (_37659_, _37595_, _36090_);
  nor (_37669_, _37659_, _37648_);
  not (_37680_, _37669_);
  and (_37691_, _36299_, _36551_);
  nor (_37701_, _37691_, _37680_);
  and (_37712_, _37099_, _36551_);
  and (_37723_, _36200_, _36551_);
  nor (_37733_, _37723_, _37712_);
  and (_37744_, _37733_, _36704_);
  and (_37755_, _37744_, _37701_);
  and (_37766_, _37755_, _37637_);
  and (_37777_, _37110_, _35530_);
  not (_37788_, _37777_);
  or (_37799_, _36989_, _36496_);
  and (_37810_, _37799_, _36562_);
  and (_37821_, _37275_, _36551_);
  nor (_37832_, _37821_, _37810_);
  and (_37843_, _37832_, _37788_);
  and (_37854_, _37843_, _36288_);
  and (_37865_, _37854_, _37766_);
  nor (_37876_, _37865_, _35564_);
  and (_37887_, _36693_, _33772_);
  and (_37898_, _37887_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37909_, _33783_, _36233_);
  and (_37920_, _37909_, _35530_);
  or (_37931_, _37920_, _37898_);
  nor (_37942_, _37931_, _37876_);
  nor (_37953_, _37942_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37964_, _37953_, _37573_);
  nor (_37975_, _37964_, _37563_);
  and (_37986_, _37975_, _36452_);
  and (_09532_, _37986_, _41991_);
  and (_38007_, _28087_, _25102_);
  and (_38018_, _24795_, _24665_);
  and (_38029_, _38018_, _25276_);
  and (_38040_, _38029_, _24960_);
  and (_38051_, _38040_, _30003_);
  and (_38062_, _38051_, _38007_);
  not (_38073_, _38062_);
  nor (_38084_, _21044_, _15690_);
  and (_38095_, _26681_, _21022_);
  nor (_38106_, _27705_, _38095_);
  and (_38117_, _38106_, _27847_);
  and (_38128_, _38117_, _38084_);
  and (_38139_, _38128_, _29003_);
  nor (_38150_, _38139_, _17747_);
  not (_38161_, _38150_);
  and (_38172_, _38161_, _27825_);
  and (_38183_, _38172_, _27662_);
  and (_38194_, _38183_, _27400_);
  nor (_38205_, _38194_, _38073_);
  and (_38216_, _38040_, _25102_);
  and (_38227_, _38216_, _24197_);
  and (_38238_, _38227_, _29992_);
  and (_38249_, _38238_, _28087_);
  and (_38260_, _38073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_38271_, _38249_);
  nor (_38282_, _38139_, _16907_);
  not (_38293_, _38282_);
  and (_38304_, _38293_, _33367_);
  and (_38315_, _38304_, _33344_);
  and (_38326_, _38315_, _33258_);
  nor (_38337_, _38326_, _38271_);
  nor (_38348_, _38337_, _38260_);
  and (_38359_, _38073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_38370_, _38139_, _17932_);
  not (_38381_, _38370_);
  and (_38391_, _38381_, _32666_);
  and (_38402_, _38391_, _32524_);
  nor (_38413_, _38402_, _38271_);
  nor (_38423_, _38413_, _38359_);
  and (_38434_, _38073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_38445_, _38139_, _18095_);
  nor (_38455_, _38445_, _31903_);
  and (_38466_, _38455_, _31848_);
  and (_38477_, _38466_, _31816_);
  nor (_38487_, _38477_, _38271_);
  nor (_38498_, _38487_, _38434_);
  and (_38509_, _38073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_38519_, _38139_, _18465_);
  nor (_38530_, _38519_, _30936_);
  and (_38541_, _38530_, _31219_);
  and (_38552_, _38541_, _31077_);
  nor (_38563_, _38552_, _38271_);
  nor (_38574_, _38563_, _38509_);
  and (_38585_, _38073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_38588_, _38139_, _18967_);
  not (_38589_, _38588_);
  and (_38590_, _38589_, _30317_);
  and (_38591_, _38590_, _30350_);
  and (_38592_, _38591_, _30230_);
  nor (_38593_, _38592_, _38271_);
  nor (_38594_, _38593_, _38585_);
  and (_38595_, _38073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_38596_, _38139_, _18803_);
  not (_38597_, _38596_);
  and (_38598_, _38597_, _29762_);
  and (_38599_, _38598_, _29600_);
  nor (_38600_, _38599_, _38073_);
  nor (_38601_, _38600_, _38595_);
  nor (_38602_, _38062_, _24356_);
  nor (_38603_, _38139_, _19348_);
  not (_38604_, _38603_);
  and (_38605_, _38604_, _29090_);
  and (_38606_, _38605_, _29057_);
  and (_38607_, _38606_, _28970_);
  not (_38608_, _38607_);
  and (_38609_, _38608_, _38062_);
  nor (_38610_, _38609_, _38602_);
  and (_38611_, _38610_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38612_, _38611_, _38601_);
  and (_38613_, _38612_, _38594_);
  and (_38614_, _38613_, _38574_);
  and (_38615_, _38614_, _38498_);
  and (_38616_, _38615_, _38423_);
  and (_38617_, _38616_, _38348_);
  nor (_38618_, _38062_, _24817_);
  and (_38619_, _38618_, _38617_);
  nor (_38620_, _38618_, _38617_);
  nor (_38621_, _38620_, _38619_);
  and (_38622_, _38621_, _24521_);
  nor (_38623_, _38622_, _24861_);
  nor (_38624_, _38623_, _38249_);
  nor (_38625_, _38624_, _38205_);
  nor (_09553_, _38625_, rst);
  not (_38626_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_38627_, _38610_, _38626_);
  nor (_38628_, _38610_, _38626_);
  nor (_38629_, _38628_, _38627_);
  and (_38630_, _38629_, _24521_);
  nor (_38631_, _38630_, _24367_);
  nor (_38632_, _38631_, _38249_);
  nor (_38633_, _38632_, _38609_);
  nand (_10678_, _38633_, _41991_);
  nor (_38634_, _38611_, _38601_);
  nor (_38635_, _38634_, _38612_);
  nor (_38636_, _38635_, _23931_);
  nor (_38637_, _38636_, _24233_);
  nor (_38638_, _38637_, _38249_);
  nor (_38639_, _38638_, _38600_);
  nand (_10689_, _38639_, _41991_);
  nor (_38640_, _38612_, _38594_);
  nor (_38641_, _38640_, _38613_);
  nor (_38642_, _38641_, _23931_);
  nor (_38643_, _38642_, _23986_);
  nor (_38644_, _38643_, _38249_);
  nor (_38645_, _38644_, _38593_);
  nand (_10700_, _38645_, _41991_);
  nor (_38646_, _38613_, _38574_);
  nor (_38647_, _38646_, _38614_);
  nor (_38648_, _38647_, _23931_);
  nor (_38649_, _38648_, _25036_);
  nor (_38650_, _38649_, _38249_);
  nor (_38651_, _38650_, _38563_);
  nor (_10711_, _38651_, rst);
  nor (_38652_, _38614_, _38498_);
  nor (_38653_, _38652_, _38615_);
  nor (_38654_, _38653_, _23931_);
  nor (_38655_, _38654_, _25211_);
  nor (_38656_, _38655_, _38249_);
  nor (_38657_, _38656_, _38487_);
  nor (_10722_, _38657_, rst);
  nor (_38658_, _38615_, _38423_);
  nor (_38659_, _38658_, _38616_);
  nor (_38660_, _38659_, _23931_);
  nor (_38661_, _38660_, _24708_);
  nor (_38662_, _38661_, _38249_);
  nor (_38663_, _38662_, _38413_);
  nor (_10733_, _38663_, rst);
  nor (_38664_, _38616_, _38348_);
  nor (_38665_, _38664_, _38617_);
  nor (_38666_, _38665_, _23931_);
  nor (_38667_, _38666_, _24554_);
  nor (_38668_, _38667_, _38249_);
  nor (_38669_, _38668_, _38337_);
  nor (_10744_, _38669_, rst);
  and (_38670_, _38007_, _31425_);
  nand (_38671_, _38670_, _38040_);
  nor (_38672_, _38671_, _28011_);
  and (_38673_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15624_);
  and (_38674_, _38673_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38675_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38676_, _38675_, _38674_);
  or (_38677_, _38676_, _38672_);
  nor (_38678_, _27847_, _17573_);
  nor (_38679_, _28556_, _18465_);
  nor (_38680_, _17747_, _16413_);
  and (_38681_, _38680_, _27149_);
  and (_38682_, _38681_, _25854_);
  and (_38683_, _38682_, _25898_);
  and (_38684_, _38683_, _26507_);
  and (_38685_, _38684_, _25550_);
  or (_38686_, _38685_, _27171_);
  and (_38687_, _27236_, _17747_);
  and (_38688_, _17083_, _16084_);
  and (_38689_, _17399_, _16413_);
  and (_38690_, _38689_, _38688_);
  and (_38691_, _38690_, _38687_);
  and (_38692_, _17235_, _16248_);
  and (_38693_, _38692_, _38691_);
  nor (_38694_, _38693_, _26452_);
  and (_38695_, _26452_, _17235_);
  nor (_38696_, _38695_, _38694_);
  and (_38697_, _38696_, _38686_);
  nor (_38698_, _26452_, _16589_);
  and (_38699_, _26452_, _16589_);
  nor (_38700_, _38699_, _38698_);
  and (_38701_, _38700_, _38697_);
  and (_38702_, _38701_, _27313_);
  nor (_38703_, _38701_, _27313_);
  nor (_38704_, _38703_, _38702_);
  and (_38705_, _38704_, _27084_);
  and (_38706_, _26452_, _27313_);
  nor (_38707_, _38706_, _28284_);
  nor (_38708_, _38707_, _27367_);
  or (_38709_, _38708_, _38705_);
  or (_38710_, _38709_, _38679_);
  and (_38711_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_38712_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38713_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38714_, _38713_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38715_, _38714_, _38712_);
  nor (_38716_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38717_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38718_, _38717_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38719_, _38718_, _38716_);
  nor (_38720_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38721_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38722_, _38721_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38723_, _38722_, _38720_);
  not (_38724_, _38723_);
  nor (_38725_, _38724_, _28175_);
  nor (_38726_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38727_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38728_, _38727_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38729_, _38728_, _38726_);
  and (_38730_, _38729_, _38725_);
  nor (_38731_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38732_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38733_, _38732_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38734_, _38733_, _38731_);
  and (_38735_, _38734_, _38730_);
  and (_38736_, _38735_, _38719_);
  nor (_38737_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38738_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38739_, _38738_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38740_, _38739_, _38737_);
  and (_38741_, _38740_, _38736_);
  and (_38742_, _38741_, _38715_);
  nor (_38743_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38744_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38745_, _38744_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38746_, _38745_, _38743_);
  and (_38747_, _38746_, _38742_);
  nor (_38748_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38749_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38750_, _38749_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38751_, _38750_, _38748_);
  nor (_38752_, _38751_, _38747_);
  and (_38753_, _38751_, _38747_);
  or (_38754_, _38753_, _38752_);
  nor (_38755_, _38754_, _28153_);
  and (_38756_, _20736_, _15690_);
  or (_38757_, _38756_, _38755_);
  or (_38758_, _38757_, _38711_);
  or (_38759_, _38758_, _38710_);
  nor (_38760_, _38759_, _38678_);
  nand (_38761_, _38760_, _38674_);
  and (_38762_, _38761_, _41991_);
  and (_12690_, _38762_, _38677_);
  and (_38763_, _38007_, _30720_);
  and (_38764_, _38763_, _38040_);
  nor (_38765_, _38764_, _38674_);
  not (_38766_, _38765_);
  nand (_38767_, _38766_, _28011_);
  not (_38768_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_38769_, _38765_, _38768_);
  and (_38770_, _38769_, _41991_);
  and (_12711_, _38770_, _38767_);
  nor (_38771_, _38671_, _29221_);
  and (_38772_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38773_, _38772_, _38674_);
  or (_38774_, _38773_, _38771_);
  nor (_38775_, _27847_, _16413_);
  nor (_38776_, _28556_, _18095_);
  nor (_38777_, _27367_, _19348_);
  nor (_38778_, _28284_, _27346_);
  not (_38779_, _38778_);
  nor (_38780_, _38779_, _27258_);
  nor (_38781_, _38780_, _25822_);
  and (_38782_, _38780_, _25822_);
  nor (_38783_, _38782_, _38781_);
  and (_38784_, _38783_, _27084_);
  or (_38785_, _38784_, _38777_);
  or (_38786_, _38785_, _38776_);
  and (_38787_, _23339_, _21044_);
  and (_38788_, _38724_, _28175_);
  nor (_38789_, _38788_, _38725_);
  and (_38790_, _38789_, _26692_);
  and (_38791_, _20514_, _15690_);
  or (_38792_, _38791_, _38790_);
  or (_38793_, _38792_, _38787_);
  or (_38794_, _38793_, _38786_);
  nor (_38795_, _38794_, _38775_);
  nand (_38796_, _38795_, _38674_);
  and (_38797_, _38796_, _41991_);
  and (_13606_, _38797_, _38774_);
  nor (_38798_, _38671_, _29894_);
  and (_38799_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38800_, _38799_, _38674_);
  or (_38801_, _38800_, _38798_);
  nor (_38802_, _27847_, _17399_);
  nor (_38803_, _28556_, _17932_);
  and (_38804_, _38681_, _26452_);
  and (_38805_, _38687_, _16413_);
  and (_38806_, _38805_, _27171_);
  nor (_38807_, _38806_, _38804_);
  and (_38808_, _38807_, _17399_);
  nor (_38809_, _38807_, _17399_);
  or (_38810_, _38809_, _30186_);
  nor (_38811_, _38810_, _38808_);
  nor (_38812_, _27367_, _18803_);
  or (_38813_, _38812_, _38811_);
  or (_38814_, _38813_, _38803_);
  and (_38815_, _22357_, _21044_);
  nor (_38816_, _38729_, _38725_);
  nor (_38817_, _38816_, _38730_);
  and (_38818_, _38817_, _26692_);
  and (_38819_, _20545_, _15690_);
  or (_38820_, _38819_, _38818_);
  or (_38821_, _38820_, _38815_);
  or (_38822_, _38821_, _38814_);
  nor (_38823_, _38822_, _38802_);
  nand (_38824_, _38823_, _38674_);
  and (_38825_, _38824_, _41991_);
  and (_13615_, _38825_, _38801_);
  nor (_38826_, _38671_, _30578_);
  and (_38827_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38828_, _38827_, _38674_);
  or (_38829_, _38828_, _38826_);
  nor (_38830_, _27847_, _16084_);
  nor (_38831_, _28556_, _16907_);
  and (_38832_, _38805_, _17399_);
  and (_38833_, _38832_, _27171_);
  and (_38834_, _38682_, _26452_);
  nor (_38835_, _38834_, _38833_);
  and (_38836_, _38835_, _16084_);
  nor (_38837_, _38835_, _16084_);
  nor (_38838_, _38837_, _38836_);
  and (_38839_, _38838_, _27084_);
  nor (_38840_, _27367_, _18967_);
  or (_38841_, _38840_, _38839_);
  or (_38842_, _38841_, _38831_);
  and (_38843_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38844_, _38734_, _38730_);
  nor (_38845_, _38844_, _38735_);
  and (_38846_, _38845_, _26692_);
  and (_38847_, _20577_, _15690_);
  or (_38848_, _38847_, _38846_);
  or (_38849_, _38848_, _38843_);
  or (_38850_, _38849_, _38842_);
  nor (_38851_, _38850_, _38830_);
  nand (_38852_, _38851_, _38674_);
  and (_38853_, _38852_, _41991_);
  and (_13625_, _38853_, _38829_);
  nor (_38854_, _38671_, _31327_);
  and (_38855_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38856_, _38855_, _38674_);
  or (_38857_, _38856_, _38854_);
  nor (_38858_, _27847_, _17083_);
  nor (_38859_, _38684_, _27171_);
  nor (_38860_, _38683_, _26507_);
  not (_38861_, _38860_);
  and (_38862_, _38861_, _38859_);
  and (_38863_, _38832_, _16084_);
  nor (_38864_, _38863_, _17083_);
  nor (_38865_, _38864_, _38691_);
  nor (_38866_, _38865_, _26452_);
  nor (_38867_, _38866_, _38862_);
  nor (_38868_, _38867_, _30186_);
  nor (_38869_, _27367_, _18465_);
  or (_38870_, _38869_, _38868_);
  or (_38871_, _38870_, _28567_);
  and (_38872_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_38873_, _38735_, _38719_);
  nor (_38874_, _38873_, _38736_);
  and (_38875_, _38874_, _26692_);
  and (_38876_, _20609_, _15690_);
  or (_38877_, _38876_, _38875_);
  or (_38878_, _38877_, _38872_);
  or (_38879_, _38878_, _38871_);
  nor (_38880_, _38879_, _38858_);
  nand (_38881_, _38880_, _38674_);
  and (_38882_, _38881_, _41991_);
  and (_13635_, _38882_, _38857_);
  nor (_38883_, _38671_, _32022_);
  and (_38884_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_38885_, _38884_, _38674_);
  or (_38886_, _38885_, _38883_);
  nor (_38887_, _27847_, _16248_);
  nor (_38888_, _28556_, _19348_);
  nor (_38889_, _38691_, _26452_);
  nor (_38890_, _38889_, _38859_);
  nor (_38891_, _38890_, _25550_);
  and (_38892_, _38890_, _25550_);
  nor (_38893_, _38892_, _38891_);
  and (_38894_, _38893_, _27084_);
  and (_38895_, _26452_, _16248_);
  nor (_38896_, _26452_, _18106_);
  or (_38897_, _38896_, _27367_);
  nor (_38898_, _38897_, _38895_);
  or (_38899_, _38898_, _38894_);
  or (_38900_, _38899_, _38888_);
  and (_38901_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_38902_, _38740_, _38736_);
  not (_38903_, _38902_);
  nor (_38904_, _38741_, _28153_);
  and (_38905_, _38904_, _38903_);
  and (_38906_, _20641_, _15690_);
  or (_38907_, _38906_, _38905_);
  or (_38908_, _38907_, _38901_);
  or (_38909_, _38908_, _38900_);
  nor (_38910_, _38909_, _38887_);
  nand (_38911_, _38910_, _38674_);
  and (_38912_, _38911_, _41991_);
  and (_13645_, _38912_, _38886_);
  nor (_38913_, _38671_, _32842_);
  and (_38914_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_38915_, _38914_, _38674_);
  or (_38916_, _38915_, _38913_);
  nor (_38917_, _27847_, _17235_);
  nor (_38918_, _28556_, _18803_);
  and (_38919_, _38691_, _16248_);
  nor (_38920_, _38919_, _26452_);
  not (_38921_, _38920_);
  and (_38922_, _38921_, _38686_);
  and (_38923_, _38922_, _17235_);
  nor (_38924_, _38922_, _17235_);
  or (_38925_, _38924_, _38923_);
  and (_38926_, _38925_, _27084_);
  nor (_38927_, _26452_, _18509_);
  or (_38928_, _38927_, _27367_);
  nor (_38929_, _38928_, _38695_);
  or (_38930_, _38929_, _38926_);
  or (_38931_, _38930_, _38918_);
  and (_38932_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_38933_, _38741_, _38715_);
  nor (_38934_, _38933_, _38742_);
  and (_38935_, _38934_, _26692_);
  and (_38936_, _20672_, _15690_);
  or (_38937_, _38936_, _38935_);
  or (_38938_, _38937_, _38932_);
  or (_38939_, _38938_, _38931_);
  nor (_38940_, _38939_, _38917_);
  nand (_38941_, _38940_, _38674_);
  and (_38942_, _38941_, _41991_);
  and (_13655_, _38942_, _38916_);
  nor (_38943_, _38671_, _33554_);
  and (_38944_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38945_, _38944_, _38674_);
  or (_38946_, _38945_, _38943_);
  nor (_38947_, _27847_, _16589_);
  nor (_38948_, _28556_, _18967_);
  and (_38949_, _38697_, _16589_);
  nor (_38950_, _38697_, _16589_);
  nor (_38951_, _38950_, _38949_);
  nor (_38952_, _38951_, _30186_);
  nor (_38953_, _26452_, _16918_);
  or (_38954_, _38953_, _27367_);
  nor (_38955_, _38954_, _38699_);
  or (_38956_, _38955_, _38952_);
  or (_38957_, _38956_, _38948_);
  and (_38958_, _21044_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_38959_, _38746_, _38742_);
  not (_38960_, _38959_);
  nor (_38961_, _38747_, _28153_);
  and (_38962_, _38961_, _38960_);
  and (_38963_, _20704_, _15690_);
  or (_38964_, _38963_, _38962_);
  or (_38965_, _38964_, _38958_);
  or (_38966_, _38965_, _38957_);
  nor (_38967_, _38966_, _38947_);
  nand (_38968_, _38967_, _38674_);
  and (_38969_, _38968_, _41991_);
  and (_13665_, _38969_, _38946_);
  nand (_38970_, _38766_, _29221_);
  not (_38971_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_38972_, _38765_, _38971_);
  and (_38973_, _38972_, _41991_);
  and (_13674_, _38973_, _38970_);
  nand (_38974_, _38766_, _29894_);
  not (_38975_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_38976_, _38765_, _38975_);
  and (_38977_, _38976_, _41991_);
  and (_13683_, _38977_, _38974_);
  nand (_38978_, _38766_, _30578_);
  not (_38979_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_38980_, _38765_, _38979_);
  and (_38981_, _38980_, _41991_);
  and (_13693_, _38981_, _38978_);
  nand (_38982_, _38766_, _31327_);
  or (_38983_, _38766_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38984_, _38983_, _41991_);
  and (_13703_, _38984_, _38982_);
  nand (_38985_, _38766_, _32022_);
  or (_38986_, _38766_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38987_, _38986_, _41991_);
  and (_13713_, _38987_, _38985_);
  nand (_38988_, _38766_, _32842_);
  or (_38989_, _38766_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38990_, _38989_, _41991_);
  and (_13722_, _38990_, _38988_);
  nand (_38994_, _38766_, _33554_);
  or (_38995_, _38766_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38996_, _38995_, _41991_);
  and (_13731_, _38996_, _38994_);
  not (_38997_, _24665_);
  and (_38998_, _25287_, _24795_);
  and (_38999_, _38998_, _38997_);
  not (_39000_, _28753_);
  nor (_39001_, _39000_, _24949_);
  and (_39002_, _39001_, _38999_);
  not (_39003_, _28720_);
  nor (_39012_, _39003_, _28687_);
  not (_39018_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_39024_, _28720_, _39018_);
  or (_39028_, _39024_, _39012_);
  and (_39029_, _39028_, _39002_);
  and (_39030_, _28087_, _24455_);
  nor (_39031_, _24665_, _24949_);
  and (_39032_, _38998_, _39031_);
  and (_39033_, _39032_, _39030_);
  nor (_39034_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_39035_, _39034_);
  nand (_39036_, _39035_, _28687_);
  and (_39037_, _39032_, _28753_);
  and (_39038_, _39034_, _39018_);
  nor (_39039_, _39038_, _39037_);
  and (_39040_, _39039_, _39036_);
  or (_39041_, _39040_, _39033_);
  or (_39042_, _39041_, _39029_);
  nand (_39043_, _39033_, _38194_);
  and (_39044_, _39043_, _39042_);
  and (_16533_, _39044_, _41991_);
  not (_39045_, _39033_);
  nor (_39046_, _39045_, _38599_);
  not (_39047_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_39048_, _39037_, _30003_);
  nand (_39049_, _39048_, _39047_);
  and (_39050_, _39049_, _39045_);
  or (_39051_, _39048_, _29308_);
  and (_39053_, _39051_, _39050_);
  or (_39055_, _39053_, _39046_);
  and (_21467_, _39055_, _41991_);
  nand (_39056_, _39033_, _38592_);
  or (_39057_, _20799_, _20768_);
  or (_39058_, _39057_, _20831_);
  or (_39059_, _39058_, _20874_);
  or (_39060_, _39059_, _20948_);
  or (_39061_, _39060_, _20980_);
  or (_39062_, _39061_, _20439_);
  and (_39063_, _39062_, _15690_);
  or (_39064_, _28218_, _26605_);
  not (_39065_, _28207_);
  nand (_39066_, _39065_, _26605_);
  and (_39067_, _39066_, _25385_);
  and (_39068_, _39067_, _39064_);
  not (_39069_, _25407_);
  nand (_39070_, _27018_, _39069_);
  nor (_39071_, _28153_, _28164_);
  and (_39072_, _39071_, _39070_);
  and (_39073_, _38692_, _22258_);
  and (_39074_, _38690_, _21044_);
  nand (_39075_, _39074_, _39073_);
  nand (_39076_, _39075_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_39077_, _39076_, _39072_);
  or (_39078_, _39077_, _39068_);
  or (_39079_, _39078_, _31577_);
  or (_39080_, _39079_, _39063_);
  nor (_39081_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_39082_, _39081_, _39037_);
  and (_39083_, _39082_, _39080_);
  not (_39084_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_39085_, _30720_, _39084_);
  or (_39086_, _39085_, _30730_);
  and (_39087_, _39086_, _39037_);
  or (_39088_, _39087_, _39033_);
  or (_39089_, _39088_, _39083_);
  and (_39090_, _39089_, _39056_);
  and (_21479_, _39090_, _41991_);
  nor (_39094_, _39045_, _38552_);
  and (_39100_, _39037_, _31425_);
  nand (_39105_, _39100_, _28687_);
  or (_39112_, _39100_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_39119_, _39112_, _39045_);
  and (_39129_, _39119_, _39105_);
  or (_39130_, _39129_, _39094_);
  and (_21491_, _39130_, _41991_);
  nor (_39131_, _39045_, _38477_);
  not (_39132_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_39133_, _39033_, _39132_);
  nor (_39134_, _39133_, _39131_);
  not (_39135_, _39037_);
  nor (_39136_, _39135_, _32142_);
  nor (_39137_, _39136_, _39134_);
  and (_39138_, _32131_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_39139_, _39138_, _32175_);
  and (_39140_, _39139_, _39037_);
  or (_39141_, _39140_, _39137_);
  and (_21503_, _39141_, _41991_);
  and (_39142_, _39002_, _32930_);
  nand (_39143_, _39142_, _28687_);
  or (_39144_, _39142_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_39145_, _39144_, _39143_);
  and (_39146_, _39145_, _39045_);
  nor (_39147_, _39045_, _38402_);
  or (_39148_, _39147_, _39146_);
  and (_21515_, _39148_, _41991_);
  nor (_39149_, _39045_, _38326_);
  and (_39150_, _33652_, _29308_);
  or (_39151_, _33652_, _31121_);
  nand (_39152_, _39151_, _39037_);
  or (_39153_, _39152_, _39150_);
  and (_39154_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_39155_, _26692_, _26942_);
  and (_39156_, _26561_, _25385_);
  or (_39157_, _39156_, _39155_);
  and (_39158_, _39157_, _39154_);
  nand (_39159_, _39154_, _27847_);
  and (_39160_, _39159_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_39161_, _39160_, _39037_);
  or (_39162_, _39161_, _39158_);
  and (_39163_, _39162_, _39045_);
  and (_39167_, _39163_, _39153_);
  or (_39178_, _39167_, _39149_);
  and (_21527_, _39178_, _41991_);
  not (_39181_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39182_, _38673_, _39181_);
  not (_39191_, _39182_);
  nor (_39199_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_39200_, _39199_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_39201_, _24455_, _25102_);
  not (_39202_, _24795_);
  and (_39203_, _25276_, _39202_);
  and (_39204_, _39203_, _28087_);
  and (_39205_, _39204_, _39201_);
  and (_39206_, _39205_, _39031_);
  nor (_39207_, _39206_, _39200_);
  nor (_39208_, _39207_, _28011_);
  and (_39209_, _25276_, _25102_);
  and (_39210_, _39209_, _24806_);
  and (_39211_, _39210_, _39001_);
  and (_39212_, _39211_, _28720_);
  and (_39213_, _39212_, _28687_);
  nor (_39214_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_39215_, _39200_, _39182_);
  nor (_39216_, _39215_, _39206_);
  not (_39217_, _39216_);
  nor (_39218_, _39217_, _39214_);
  not (_39219_, _39218_);
  nor (_39220_, _39219_, _39213_);
  or (_39221_, _39220_, _39208_);
  and (_39222_, _39221_, _39191_);
  nor (_39223_, _39191_, _38760_);
  or (_39224_, _39223_, _39222_);
  and (_22302_, _39224_, _41991_);
  nor (_39225_, _39207_, _29221_);
  and (_39226_, _39211_, _24455_);
  and (_39227_, _39226_, _28687_);
  nor (_39228_, _39226_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_39229_, _39228_, _39217_);
  not (_39230_, _39229_);
  nor (_39231_, _39230_, _39227_);
  or (_39232_, _39231_, _39225_);
  and (_39233_, _39232_, _39191_);
  nor (_39234_, _39191_, _38795_);
  or (_39235_, _39234_, _39233_);
  and (_24162_, _39235_, _41991_);
  and (_39236_, _39182_, _38823_);
  nor (_39237_, _39207_, _29894_);
  and (_39238_, _39211_, _30003_);
  and (_39239_, _39238_, _28687_);
  nor (_39240_, _39238_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_39241_, _39240_, _39217_);
  not (_39242_, _39241_);
  nor (_39243_, _39242_, _39239_);
  nor (_39244_, _39243_, _39182_);
  not (_39245_, _39244_);
  nor (_39246_, _39245_, _39237_);
  nor (_39247_, _39246_, _39236_);
  and (_24174_, _39247_, _41991_);
  nor (_39248_, _39207_, _30578_);
  nor (_39249_, _25113_, _24949_);
  and (_39250_, _39249_, _25276_);
  and (_39251_, _28753_, _24806_);
  and (_39252_, _39251_, _39250_);
  not (_39253_, _39252_);
  and (_39254_, _39216_, _39253_);
  and (_39255_, _39254_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_39256_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_39257_, _30720_, _39256_);
  nor (_39258_, _39257_, _30730_);
  and (_39259_, _39216_, _39252_);
  not (_39260_, _39259_);
  nor (_39261_, _39260_, _39258_);
  nor (_39262_, _39261_, _39255_);
  and (_39263_, _39262_, _39191_);
  not (_39264_, _39263_);
  nor (_39265_, _39264_, _39248_);
  and (_39266_, _39182_, _38851_);
  or (_39267_, _39266_, _39265_);
  nor (_24186_, _39267_, rst);
  nor (_39268_, _39207_, _31327_);
  and (_39269_, _39254_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_39270_, _31436_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_39271_, _39270_, _31447_);
  nor (_39272_, _39271_, _39260_);
  nor (_39273_, _39272_, _39269_);
  and (_39274_, _39273_, _39191_);
  not (_39275_, _39274_);
  nor (_39276_, _39275_, _39268_);
  and (_39277_, _39182_, _38880_);
  or (_39278_, _39277_, _39276_);
  nor (_24198_, _39278_, rst);
  nor (_39279_, _39207_, _32022_);
  and (_39280_, _39211_, _32120_);
  and (_39281_, _39280_, _28687_);
  nor (_39282_, _39280_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_39283_, _39282_, _39217_);
  not (_39284_, _39283_);
  nor (_39285_, _39284_, _39281_);
  or (_39286_, _39285_, _39279_);
  and (_39287_, _39286_, _39191_);
  nor (_39288_, _39191_, _38910_);
  or (_39289_, _39288_, _39287_);
  and (_24210_, _39289_, _41991_);
  nor (_39290_, _39207_, _32842_);
  and (_39291_, _39211_, _32930_);
  and (_39292_, _39291_, _28687_);
  nor (_39293_, _39291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_39294_, _39293_, _39217_);
  not (_39295_, _39294_);
  nor (_39296_, _39295_, _39292_);
  or (_39297_, _39296_, _39290_);
  and (_39298_, _39297_, _39191_);
  nor (_39299_, _39191_, _38940_);
  or (_39300_, _39299_, _39298_);
  and (_24222_, _39300_, _41991_);
  nor (_39301_, _39207_, _33554_);
  and (_39302_, _39211_, _33652_);
  and (_39303_, _39302_, _28687_);
  nor (_39304_, _39302_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_39305_, _39304_, _39217_);
  not (_39306_, _39305_);
  nor (_39307_, _39306_, _39303_);
  or (_39308_, _39307_, _39301_);
  and (_39309_, _39308_, _39191_);
  nor (_39310_, _39191_, _38967_);
  or (_39311_, _39310_, _39309_);
  and (_24234_, _39311_, _41991_);
  and (_39312_, _38216_, _28720_);
  nand (_39313_, _39312_, _28687_);
  or (_39314_, _39312_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39315_, _39314_, _28753_);
  and (_39316_, _39315_, _39313_);
  and (_39317_, _38040_, _39201_);
  nand (_39318_, _39317_, _38194_);
  or (_39319_, _39317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_39320_, _39319_, _28087_);
  and (_39321_, _39320_, _39318_);
  not (_39322_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_39323_, _28065_, _39322_);
  or (_39324_, _39323_, rst);
  or (_39325_, _39324_, _39321_);
  or (_35472_, _39325_, _39316_);
  nor (_39326_, _38997_, _24949_);
  and (_39327_, _38998_, _39326_);
  and (_39328_, _39327_, _28720_);
  nand (_39329_, _39328_, _28687_);
  or (_39330_, _39328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_39331_, _39330_, _28753_);
  and (_39332_, _39331_, _39329_);
  and (_39333_, _39327_, _24455_);
  not (_39334_, _39333_);
  nor (_39335_, _39334_, _38194_);
  not (_39336_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_39337_, _39333_, _39336_);
  or (_39338_, _39337_, _39335_);
  and (_39339_, _39338_, _28087_);
  nor (_39340_, _28065_, _39336_);
  or (_39341_, _39340_, rst);
  or (_39342_, _39341_, _39339_);
  or (_35495_, _39342_, _39332_);
  and (_39343_, _39202_, _24665_);
  and (_39344_, _39343_, _39250_);
  and (_39345_, _39344_, _28720_);
  nand (_39346_, _39345_, _28687_);
  or (_39347_, _39345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_39348_, _39347_, _28753_);
  and (_39349_, _39348_, _39346_);
  and (_39350_, _39203_, _39326_);
  and (_39351_, _39350_, _39201_);
  not (_39352_, _39351_);
  nor (_39353_, _39352_, _38194_);
  not (_39354_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_39355_, _39351_, _39354_);
  or (_39356_, _39355_, _39353_);
  and (_39357_, _39356_, _28087_);
  nor (_39358_, _28065_, _39354_);
  or (_39359_, _39358_, rst);
  or (_39360_, _39359_, _39357_);
  or (_35518_, _39360_, _39349_);
  and (_39361_, _39343_, _25298_);
  and (_39362_, _39361_, _28720_);
  nand (_39363_, _39362_, _28687_);
  or (_39364_, _39362_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_39365_, _39364_, _28753_);
  and (_39366_, _39365_, _39363_);
  nor (_39367_, _25276_, _24795_);
  and (_39368_, _39326_, _39367_);
  and (_39369_, _39368_, _39201_);
  not (_39370_, _39369_);
  nor (_39371_, _39370_, _38194_);
  not (_39372_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_39373_, _39369_, _39372_);
  or (_39374_, _39373_, _39371_);
  and (_39375_, _39374_, _28087_);
  nor (_39382_, _28065_, _39372_);
  or (_39393_, _39382_, rst);
  or (_39404_, _39393_, _39375_);
  or (_35541_, _39404_, _39366_);
  not (_39419_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_39429_, _39317_, _39419_);
  nand (_39440_, _38216_, _24455_);
  nor (_39451_, _39440_, _28687_);
  or (_39462_, _39451_, _39429_);
  and (_39473_, _39462_, _28753_);
  and (_39484_, _39317_, _38608_);
  or (_39495_, _39484_, _39429_);
  and (_39506_, _39495_, _28087_);
  nor (_39517_, _28065_, _39419_);
  or (_39528_, _39517_, rst);
  or (_39539_, _39528_, _39506_);
  or (_41393_, _39539_, _39473_);
  and (_39560_, _38216_, _30003_);
  nand (_39571_, _39560_, _28687_);
  or (_39582_, _39560_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39588_, _39582_, _28753_);
  and (_39589_, _39588_, _39571_);
  nand (_39590_, _39317_, _38599_);
  or (_39591_, _39317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39592_, _39591_, _28087_);
  and (_39593_, _39592_, _39590_);
  not (_39594_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_39595_, _28065_, _39594_);
  or (_39596_, _39595_, rst);
  or (_39597_, _39596_, _39593_);
  or (_41394_, _39597_, _39589_);
  not (_39598_, _31458_);
  nand (_39599_, _38216_, _39598_);
  and (_39600_, _39599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39601_, _30741_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_39602_, _39601_, _30730_);
  and (_39603_, _39602_, _38216_);
  or (_39604_, _39603_, _39600_);
  and (_39605_, _39604_, _28753_);
  nand (_39606_, _39317_, _38592_);
  or (_39607_, _39317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_39608_, _39607_, _28087_);
  and (_39609_, _39608_, _39606_);
  not (_39610_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_39611_, _28065_, _39610_);
  or (_39612_, _39611_, rst);
  or (_39613_, _39612_, _39609_);
  or (_41396_, _39613_, _39605_);
  not (_39614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_39615_, _38227_, _39614_);
  nor (_39616_, _31458_, _39614_);
  or (_39617_, _39616_, _31447_);
  and (_39618_, _39617_, _38216_);
  or (_39619_, _39618_, _39615_);
  and (_39620_, _39619_, _28753_);
  nand (_39621_, _39317_, _38552_);
  or (_39622_, _39317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39623_, _39622_, _28087_);
  and (_39624_, _39623_, _39621_);
  nor (_39625_, _28065_, _39614_);
  or (_39626_, _39625_, rst);
  or (_39627_, _39626_, _39624_);
  or (_41398_, _39627_, _39620_);
  not (_39628_, _38216_);
  or (_39629_, _39628_, _32142_);
  and (_39630_, _39629_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39631_, _32131_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39632_, _39631_, _32175_);
  and (_39633_, _39632_, _38216_);
  or (_39634_, _39633_, _39630_);
  and (_39635_, _39634_, _28753_);
  nand (_39636_, _39317_, _38477_);
  or (_39637_, _39317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_39638_, _39637_, _28087_);
  and (_39639_, _39638_, _39636_);
  and (_39640_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_39641_, _39640_, rst);
  or (_39642_, _39641_, _39639_);
  or (_41400_, _39642_, _39635_);
  and (_39643_, _38216_, _32930_);
  nand (_39644_, _39643_, _28687_);
  or (_39645_, _39643_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39646_, _39645_, _28753_);
  and (_39647_, _39646_, _39644_);
  nand (_39648_, _39317_, _38402_);
  or (_39649_, _39317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39650_, _39649_, _28087_);
  and (_39651_, _39650_, _39648_);
  and (_39652_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39653_, _39652_, rst);
  or (_39654_, _39653_, _39651_);
  or (_41401_, _39654_, _39647_);
  and (_39655_, _38216_, _33652_);
  nand (_39656_, _39655_, _28687_);
  or (_39657_, _39655_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39658_, _39657_, _28753_);
  and (_39659_, _39658_, _39656_);
  nand (_39660_, _39317_, _38326_);
  or (_39661_, _39317_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39662_, _39661_, _28087_);
  and (_39663_, _39662_, _39660_);
  not (_39664_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_39665_, _28065_, _39664_);
  or (_39666_, _39665_, rst);
  or (_39667_, _39666_, _39663_);
  or (_41403_, _39667_, _39659_);
  nand (_39668_, _39333_, _28687_);
  or (_39669_, _39333_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39670_, _39669_, _28753_);
  and (_39671_, _39670_, _39668_);
  and (_39672_, _39333_, _38608_);
  not (_39673_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39674_, _39333_, _39673_);
  or (_39675_, _39674_, _39672_);
  and (_39676_, _39675_, _28087_);
  nor (_39677_, _28065_, _39673_);
  or (_39678_, _39677_, rst);
  or (_39679_, _39678_, _39676_);
  or (_41405_, _39679_, _39671_);
  and (_39680_, _39327_, _30003_);
  nand (_39681_, _39680_, _28687_);
  or (_39682_, _39680_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39683_, _39682_, _28753_);
  and (_39684_, _39683_, _39681_);
  nor (_39685_, _39334_, _38599_);
  not (_39686_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_39687_, _39333_, _39686_);
  or (_39688_, _39687_, _39685_);
  and (_39689_, _39688_, _28087_);
  nor (_39690_, _28065_, _39686_);
  or (_39691_, _39690_, rst);
  or (_39692_, _39691_, _39689_);
  or (_41407_, _39692_, _39684_);
  and (_39693_, _39327_, _30720_);
  nand (_39694_, _39693_, _28687_);
  or (_39695_, _39693_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39696_, _39695_, _28753_);
  and (_39697_, _39696_, _39694_);
  nor (_39698_, _39334_, _38592_);
  not (_39699_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_39700_, _39333_, _39699_);
  or (_39701_, _39700_, _39698_);
  and (_39702_, _39701_, _28087_);
  nor (_39703_, _28065_, _39699_);
  or (_39704_, _39703_, rst);
  or (_39705_, _39704_, _39702_);
  or (_41408_, _39705_, _39697_);
  and (_39706_, _39327_, _31425_);
  nand (_39707_, _39706_, _28687_);
  or (_39708_, _39706_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39709_, _39708_, _28753_);
  and (_39710_, _39709_, _39707_);
  nor (_39711_, _39334_, _38552_);
  and (_39712_, _39334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39713_, _39712_, _39711_);
  and (_39714_, _39713_, _28087_);
  and (_39715_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39716_, _39715_, rst);
  or (_39717_, _39716_, _39714_);
  or (_41410_, _39717_, _39710_);
  and (_39718_, _39327_, _32120_);
  nand (_39719_, _39718_, _28687_);
  or (_39720_, _39718_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39721_, _39720_, _28753_);
  and (_39722_, _39721_, _39719_);
  nor (_39723_, _39334_, _38477_);
  and (_39724_, _39334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39725_, _39724_, _39723_);
  and (_39726_, _39725_, _28087_);
  and (_39727_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39728_, _39727_, rst);
  or (_39729_, _39728_, _39726_);
  or (_41412_, _39729_, _39722_);
  and (_39730_, _39327_, _32930_);
  nand (_39731_, _39730_, _28687_);
  or (_39732_, _39730_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39733_, _39732_, _28753_);
  and (_39734_, _39733_, _39731_);
  nor (_39735_, _39334_, _38402_);
  and (_39736_, _39334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39737_, _39736_, _39735_);
  and (_39738_, _39737_, _28087_);
  and (_39739_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39740_, _39739_, rst);
  or (_39741_, _39740_, _39738_);
  or (_41414_, _39741_, _39734_);
  and (_39742_, _39327_, _33652_);
  nand (_39743_, _39742_, _28687_);
  or (_39744_, _39742_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39745_, _39744_, _28753_);
  and (_39746_, _39745_, _39743_);
  nor (_39747_, _39334_, _38326_);
  not (_39748_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_39749_, _39333_, _39748_);
  or (_39750_, _39749_, _39747_);
  and (_39751_, _39750_, _28087_);
  nor (_39752_, _28065_, _39748_);
  or (_39753_, _39752_, rst);
  or (_39754_, _39753_, _39751_);
  or (_41415_, _39754_, _39746_);
  nand (_39755_, _39351_, _28687_);
  or (_39756_, _39351_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39757_, _39756_, _28753_);
  and (_39758_, _39757_, _39755_);
  and (_39759_, _39351_, _38608_);
  not (_39760_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_39761_, _39351_, _39760_);
  or (_39762_, _39761_, _39759_);
  and (_39763_, _39762_, _28087_);
  nor (_39764_, _28065_, _39760_);
  or (_39765_, _39764_, rst);
  or (_39766_, _39765_, _39763_);
  or (_41417_, _39766_, _39758_);
  and (_39767_, _39344_, _30003_);
  nand (_39768_, _39767_, _28687_);
  or (_39769_, _39767_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39770_, _39769_, _28753_);
  and (_39771_, _39770_, _39768_);
  nor (_39772_, _39352_, _38599_);
  not (_39773_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_39774_, _39351_, _39773_);
  or (_39775_, _39774_, _39772_);
  and (_39776_, _39775_, _28087_);
  nor (_39777_, _28065_, _39773_);
  or (_39778_, _39777_, rst);
  or (_39779_, _39778_, _39776_);
  or (_41419_, _39779_, _39771_);
  and (_39780_, _39344_, _30720_);
  nand (_39781_, _39780_, _28687_);
  or (_39782_, _39780_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39783_, _39782_, _28753_);
  and (_39784_, _39783_, _39781_);
  nor (_39785_, _39352_, _38592_);
  not (_39786_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_39787_, _39351_, _39786_);
  or (_39788_, _39787_, _39785_);
  and (_39789_, _39788_, _28087_);
  nor (_39790_, _28065_, _39786_);
  or (_39791_, _39790_, rst);
  or (_39792_, _39791_, _39789_);
  or (_41421_, _39792_, _39784_);
  and (_39793_, _39344_, _31425_);
  nand (_39794_, _39793_, _28687_);
  or (_39796_, _39793_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39797_, _39796_, _28753_);
  and (_39798_, _39797_, _39794_);
  nor (_39799_, _39352_, _38552_);
  and (_39800_, _39352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39801_, _39800_, _39799_);
  and (_39802_, _39801_, _28087_);
  and (_39803_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39804_, _39803_, rst);
  or (_39805_, _39804_, _39802_);
  or (_41422_, _39805_, _39798_);
  and (_39806_, _39344_, _32120_);
  nand (_39807_, _39806_, _28687_);
  or (_39808_, _39806_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39809_, _39808_, _28753_);
  and (_39810_, _39809_, _39807_);
  nor (_39811_, _39352_, _38477_);
  and (_39812_, _39352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39813_, _39812_, _39811_);
  and (_39814_, _39813_, _28087_);
  and (_39815_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39816_, _39815_, rst);
  or (_39817_, _39816_, _39814_);
  or (_41424_, _39817_, _39810_);
  and (_39818_, _39344_, _32930_);
  nand (_39819_, _39818_, _28687_);
  or (_39820_, _39818_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39821_, _39820_, _28753_);
  and (_39822_, _39821_, _39819_);
  nor (_39823_, _39352_, _38402_);
  and (_39824_, _39352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39825_, _39824_, _39823_);
  and (_39830_, _39825_, _28087_);
  and (_39831_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39832_, _39831_, rst);
  or (_39833_, _39832_, _39830_);
  or (_41426_, _39833_, _39822_);
  and (_39834_, _39344_, _33652_);
  nand (_39835_, _39834_, _28687_);
  or (_39836_, _39834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39837_, _39836_, _28753_);
  and (_39838_, _39837_, _39835_);
  nor (_39839_, _39352_, _38326_);
  not (_39840_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_39841_, _39351_, _39840_);
  or (_39842_, _39841_, _39839_);
  and (_39843_, _39842_, _28087_);
  nor (_39844_, _28065_, _39840_);
  or (_39845_, _39844_, rst);
  or (_39846_, _39845_, _39843_);
  or (_41428_, _39846_, _39838_);
  and (_39847_, _39361_, _24455_);
  nand (_39848_, _39847_, _28687_);
  or (_39849_, _39847_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39850_, _39849_, _28753_);
  and (_39851_, _39850_, _39848_);
  and (_39852_, _39369_, _38608_);
  not (_39853_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_39854_, _39369_, _39853_);
  or (_39855_, _39854_, _39852_);
  and (_39856_, _39855_, _28087_);
  nor (_39857_, _28065_, _39853_);
  or (_39858_, _39857_, rst);
  or (_39859_, _39858_, _39856_);
  or (_41429_, _39859_, _39851_);
  and (_39860_, _39361_, _30003_);
  nand (_39861_, _39860_, _28687_);
  or (_39862_, _39860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39863_, _39862_, _28753_);
  and (_39864_, _39863_, _39861_);
  nor (_39865_, _39370_, _38599_);
  not (_39866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_39867_, _39369_, _39866_);
  or (_39868_, _39867_, _39865_);
  and (_39869_, _39868_, _28087_);
  nor (_39870_, _28065_, _39866_);
  or (_39871_, _39870_, rst);
  or (_39872_, _39871_, _39869_);
  or (_41431_, _39872_, _39864_);
  and (_39873_, _39361_, _30720_);
  nand (_39874_, _39873_, _28687_);
  or (_39875_, _39873_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39876_, _39875_, _28753_);
  and (_39877_, _39876_, _39874_);
  nor (_39878_, _39370_, _38592_);
  not (_39879_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_39880_, _39369_, _39879_);
  or (_39881_, _39880_, _39878_);
  and (_39882_, _39881_, _28087_);
  nor (_39883_, _28065_, _39879_);
  or (_39884_, _39883_, rst);
  or (_39885_, _39884_, _39882_);
  or (_41433_, _39885_, _39877_);
  and (_39886_, _39361_, _31425_);
  nand (_39887_, _39886_, _28687_);
  or (_39888_, _39886_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39889_, _39888_, _28753_);
  and (_39890_, _39889_, _39887_);
  nor (_39898_, _39370_, _38552_);
  and (_39899_, _39370_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39900_, _39899_, _39898_);
  and (_39901_, _39900_, _28087_);
  and (_39902_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39903_, _39902_, rst);
  or (_39904_, _39903_, _39901_);
  or (_41435_, _39904_, _39890_);
  and (_39905_, _39361_, _32120_);
  nand (_39906_, _39905_, _28687_);
  or (_39907_, _39905_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39908_, _39907_, _28753_);
  and (_39909_, _39908_, _39906_);
  nor (_39910_, _39370_, _38477_);
  and (_39911_, _39370_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39912_, _39911_, _39910_);
  and (_39913_, _39912_, _28087_);
  and (_39914_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39915_, _39914_, rst);
  or (_39916_, _39915_, _39913_);
  or (_41436_, _39916_, _39909_);
  and (_39917_, _39361_, _32930_);
  nand (_39918_, _39917_, _28687_);
  or (_39919_, _39917_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39920_, _39919_, _28753_);
  and (_39921_, _39920_, _39918_);
  nor (_39922_, _39370_, _38402_);
  and (_39923_, _39370_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39924_, _39923_, _39922_);
  and (_39925_, _39924_, _28087_);
  and (_39926_, _28076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39927_, _39926_, rst);
  or (_39928_, _39927_, _39925_);
  or (_41438_, _39928_, _39921_);
  and (_39929_, _39361_, _33652_);
  nand (_39930_, _39929_, _28687_);
  or (_39931_, _39929_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39932_, _39931_, _28753_);
  and (_39933_, _39932_, _39930_);
  nor (_39934_, _39370_, _38326_);
  not (_39935_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_39936_, _39369_, _39935_);
  or (_39937_, _39936_, _39934_);
  and (_39938_, _39937_, _28087_);
  nor (_39939_, _28065_, _39935_);
  or (_39940_, _39939_, rst);
  or (_39941_, _39940_, _39938_);
  or (_41440_, _39941_, _39933_);
  nor (_39946_, _25276_, _25102_);
  and (_39947_, _39946_, _39343_);
  and (_39948_, _39947_, _39001_);
  and (_39949_, _39948_, _28720_);
  nand (_39950_, _39949_, _28687_);
  and (_39951_, _39030_, _25113_);
  and (_39952_, _39951_, _39368_);
  not (_39953_, _39952_);
  or (_39954_, _39949_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_39955_, _39954_, _39953_);
  and (_39956_, _39955_, _39950_);
  nor (_39957_, _39953_, _38194_);
  or (_39958_, _39957_, _39956_);
  and (_41933_, _39958_, _41991_);
  and (_39959_, _25276_, _25113_);
  and (_39969_, _39959_, _39001_);
  and (_39970_, _39969_, _39343_);
  and (_39971_, _39970_, _28720_);
  nand (_39972_, _39971_, _28687_);
  and (_39973_, _39951_, _39350_);
  not (_39974_, _39973_);
  or (_39975_, _39971_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_39976_, _39975_, _39974_);
  and (_39977_, _39976_, _39972_);
  nor (_39978_, _39974_, _38194_);
  or (_39979_, _39978_, _39977_);
  and (_41936_, _39979_, _41991_);
  or (_39980_, _24444_, _30709_);
  and (_39981_, _39980_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39982_, _39981_, _39150_);
  and (_39983_, _39969_, _38018_);
  and (_39984_, _39983_, _39982_);
  and (_39985_, _39951_, _38040_);
  nand (_39986_, _39983_, _24433_);
  and (_39987_, _39986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_39988_, _39987_, _39985_);
  or (_39989_, _39988_, _39984_);
  nand (_39990_, _39985_, _38326_);
  and (_39991_, _39990_, _41991_);
  and (_41938_, _39991_, _39989_);
  not (_39992_, _39985_);
  not (_39993_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_39994_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_39995_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_39996_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39995_);
  and (_39997_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_39998_, _39997_, _39996_);
  nor (_39999_, _39998_, _39994_);
  or (_40000_, _39999_, _39993_);
  and (_40001_, _39995_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40002_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40003_, _40002_, _40001_);
  nor (_40004_, _40003_, _39994_);
  and (_40005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39995_);
  and (_40006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40007_, _40006_, _40005_);
  nand (_40008_, _40007_, _40004_);
  or (_40009_, _40008_, _40000_);
  and (_40010_, _40009_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor (_40011_, _24197_, _25102_);
  and (_40012_, _28753_, _28709_);
  and (_40013_, _40012_, _38040_);
  and (_40014_, _40013_, _40011_);
  or (_40015_, _40014_, _40010_);
  and (_40016_, _40015_, _39992_);
  nand (_40017_, _40014_, _28687_);
  and (_40018_, _40017_, _40016_);
  nor (_40019_, _39992_, _38194_);
  or (_40020_, _40019_, _40018_);
  and (_41940_, _40020_, _41991_);
  nor (_40021_, _40007_, _39994_);
  nand (_40022_, _40021_, _40003_);
  or (_40023_, _40022_, _40000_);
  and (_40024_, _40023_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_40025_, _28753_, _29992_);
  and (_40026_, _40025_, _38040_);
  and (_40027_, _40026_, _40011_);
  or (_40028_, _40027_, _40024_);
  and (_40029_, _40028_, _39992_);
  nand (_40030_, _40027_, _28687_);
  and (_40031_, _40030_, _40029_);
  nor (_40032_, _39992_, _38402_);
  or (_40033_, _40032_, _40031_);
  and (_41942_, _40033_, _41991_);
  not (_40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_40035_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40034_);
  nand (_40036_, _39999_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_40037_, _40021_, _40004_);
  or (_40038_, _40037_, _40036_);
  and (_40039_, _40038_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_40040_, _40039_, _40035_);
  nor (_40041_, _28698_, _25102_);
  and (_40042_, _40026_, _40041_);
  or (_40043_, _40042_, _40040_);
  and (_40044_, _40043_, _39992_);
  nand (_40045_, _40042_, _28687_);
  and (_40046_, _40045_, _40044_);
  nor (_40047_, _39992_, _38599_);
  or (_40048_, _40047_, _40046_);
  and (_41944_, _40048_, _41991_);
  and (_40049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_40050_, _40036_, _40022_);
  and (_40051_, _40050_, _40049_);
  and (_40052_, _40013_, _40041_);
  or (_40053_, _40052_, _40051_);
  and (_40054_, _40053_, _39992_);
  nand (_40055_, _40052_, _28687_);
  and (_40056_, _40055_, _40054_);
  nor (_40057_, _39992_, _38552_);
  or (_40058_, _40057_, _40056_);
  and (_41946_, _40058_, _41991_);
  and (_40059_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40060_, _40059_, _39995_);
  and (_40061_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40062_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39995_);
  nor (_40063_, _40062_, _40061_);
  and (_40064_, _40063_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_40065_, _40064_, _39994_);
  and (_40066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40067_, _40066_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40069_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_40070_, _40069_, _40067_);
  and (_40071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40072_, _40071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40074_, _40073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_40075_, _40074_, _40072_);
  and (_40076_, _40075_, _40070_);
  nor (_40077_, _40076_, _40065_);
  and (_40078_, _40077_, _40060_);
  and (_40079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39994_);
  not (_40080_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40081_, _40066_, _40080_);
  not (_40082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40083_, _40068_, _40082_);
  nor (_40084_, _40083_, _40081_);
  not (_40085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40086_, _40071_, _40085_);
  not (_40087_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40088_, _40073_, _40087_);
  nor (_40089_, _40088_, _40086_);
  and (_40090_, _40089_, _40084_);
  not (_40091_, _40090_);
  and (_40092_, _40091_, _40079_);
  nand (_40093_, _40060_, _40092_);
  and (_40094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41991_);
  nand (_40095_, _40094_, _40093_);
  nor (_41978_, _40095_, _40078_);
  nor (_40096_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40097_, _40096_);
  nor (_40098_, _40077_, _40092_);
  nor (_40099_, _40098_, _40097_);
  nand (_40100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41991_);
  nor (_41980_, _40100_, _40099_);
  nor (_40101_, _40098_, _40059_);
  not (_40102_, _40101_);
  and (_40103_, _40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_40104_, _40059_);
  and (_40105_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40106_, _40070_);
  or (_40107_, _40106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_40108_, _40107_, _40105_);
  not (_40109_, _40072_);
  and (_40110_, _40109_, _40070_);
  or (_40111_, _40110_, _40001_);
  and (_40112_, _40111_, _40077_);
  and (_40113_, _40112_, _40108_);
  not (_40114_, _40077_);
  and (_40115_, _40114_, _40092_);
  and (_40116_, _40088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40117_, _40116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_40118_, _40084_);
  and (_40119_, _40086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40120_, _40119_, _40118_);
  and (_40121_, _40120_, _40117_);
  and (_40122_, _40118_, _40001_);
  or (_40123_, _40122_, _40121_);
  and (_40124_, _40123_, _40115_);
  or (_40125_, _40124_, _40113_);
  and (_40126_, _40125_, _40104_);
  or (_40127_, _40126_, _40103_);
  and (_41981_, _40127_, _41991_);
  and (_40128_, _40088_, _39995_);
  or (_40129_, _40128_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40130_, _40086_, _39995_);
  nor (_40131_, _40130_, _40118_);
  and (_40132_, _40131_, _40129_);
  and (_40133_, _40118_, _40002_);
  or (_40134_, _40133_, _40132_);
  and (_40135_, _40134_, _40115_);
  and (_40136_, _40098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_40137_, _40136_, _40135_);
  and (_40138_, _40074_, _39995_);
  or (_40139_, _40106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_40140_, _40139_, _40138_);
  or (_40141_, _40110_, _40002_);
  and (_40142_, _40141_, _40077_);
  and (_40143_, _40142_, _40140_);
  or (_40144_, _40143_, _40059_);
  or (_40145_, _40144_, _40137_);
  or (_40146_, _40104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40147_, _40146_, _41991_);
  and (_41983_, _40147_, _40145_);
  nand (_40148_, _40098_, _39994_);
  nor (_40149_, _39995_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40150_, _40149_, _40059_);
  and (_40151_, _40150_, _41991_);
  and (_41985_, _40151_, _40148_);
  and (_40152_, _40098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40153_, _39995_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40154_, _40153_, _40149_);
  nor (_40155_, _40154_, _40114_);
  or (_40156_, _40155_, _40059_);
  or (_40157_, _40156_, _40152_);
  or (_40158_, _40154_, _40104_);
  and (_40159_, _40158_, _41991_);
  and (_41987_, _40159_, _40157_);
  and (_40160_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41991_);
  and (_41989_, _40160_, _40059_);
  and (_40161_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40162_, _40161_, _40101_);
  and (_42909_, _40162_, _41991_);
  and (_40163_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40164_, _40163_, _40101_);
  and (_42911_, _40164_, _41991_);
  and (_40165_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _41991_);
  and (_42913_, _40165_, _40059_);
  not (_40166_, _40081_);
  nor (_40167_, _40088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40168_, _40167_, _40086_);
  or (_40169_, _40168_, _40083_);
  and (_40170_, _40169_, _40166_);
  and (_40171_, _40170_, _40115_);
  not (_40172_, _40067_);
  or (_40173_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40174_, _40173_, _40109_);
  or (_40175_, _40174_, _40069_);
  and (_40176_, _40175_, _40172_);
  and (_40177_, _40176_, _40077_);
  or (_40178_, _40177_, _40059_);
  or (_40179_, _40178_, _40171_);
  or (_40180_, _40104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40181_, _40180_, _41991_);
  and (_42915_, _40181_, _40179_);
  nand (_40182_, _40084_, _40079_);
  or (_40183_, _40182_, _40089_);
  nor (_40184_, _40183_, _40077_);
  or (_40185_, _40075_, _40106_);
  nor (_40186_, _40185_, _40065_);
  or (_40187_, _40186_, _40059_);
  or (_40188_, _40187_, _40184_);
  or (_40189_, _40104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40190_, _40189_, _41991_);
  and (_42917_, _40190_, _40188_);
  and (_40191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _41991_);
  and (_42919_, _40191_, _40059_);
  and (_40192_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _41991_);
  and (_42921_, _40192_, _40059_);
  nand (_40193_, _40098_, _40096_);
  nor (_40194_, _40077_, _40059_);
  or (_40195_, _40194_, _39995_);
  and (_40196_, _40195_, _41991_);
  and (_42923_, _40196_, _40193_);
  and (_40197_, _40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_40198_, _40138_);
  and (_40199_, _40198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40200_, _40072_, _39995_);
  or (_40201_, _40200_, _40069_);
  or (_40202_, _40201_, _40199_);
  not (_40203_, _40069_);
  or (_40204_, _40203_, _39997_);
  and (_40205_, _40204_, _40202_);
  or (_40206_, _40205_, _40067_);
  or (_40207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39995_);
  or (_40208_, _40207_, _40172_);
  and (_40209_, _40208_, _40077_);
  and (_40210_, _40209_, _40206_);
  not (_40211_, _40128_);
  and (_40212_, _40211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_40213_, _40130_, _40083_);
  or (_40214_, _40213_, _40212_);
  not (_40215_, _40083_);
  or (_40216_, _40215_, _39997_);
  and (_40217_, _40216_, _40214_);
  or (_40218_, _40217_, _40081_);
  or (_40219_, _40207_, _40166_);
  and (_40220_, _40219_, _40115_);
  and (_40221_, _40220_, _40218_);
  or (_40222_, _40221_, _40210_);
  and (_40223_, _40222_, _40104_);
  or (_40224_, _40223_, _40197_);
  and (_42925_, _40224_, _41991_);
  and (_40225_, _40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40226_, _40198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40227_, _40226_, _40201_);
  or (_40228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39995_);
  or (_40229_, _40228_, _40203_);
  and (_40230_, _40229_, _40227_);
  or (_40231_, _40230_, _40067_);
  or (_40232_, _40172_, _40006_);
  and (_40233_, _40232_, _40077_);
  and (_40234_, _40233_, _40231_);
  and (_40235_, _40211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_40236_, _40235_, _40213_);
  or (_40237_, _40228_, _40215_);
  and (_40238_, _40237_, _40236_);
  or (_40239_, _40238_, _40081_);
  or (_40240_, _40166_, _40006_);
  and (_40241_, _40240_, _40115_);
  and (_40242_, _40241_, _40239_);
  or (_40243_, _40242_, _40234_);
  and (_40244_, _40243_, _40104_);
  or (_40245_, _40244_, _40225_);
  and (_42927_, _40245_, _41991_);
  and (_40246_, _40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_40247_, _40105_);
  and (_40248_, _40247_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_40249_, _40072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40250_, _40249_, _40069_);
  or (_40251_, _40250_, _40248_);
  or (_40252_, _40203_, _39996_);
  and (_40253_, _40252_, _40251_);
  or (_40254_, _40253_, _40067_);
  or (_40255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40256_, _40255_, _40172_);
  and (_40257_, _40256_, _40077_);
  and (_40258_, _40257_, _40254_);
  not (_40259_, _40116_);
  and (_40260_, _40259_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_40261_, _40119_, _40083_);
  or (_40262_, _40261_, _40260_);
  or (_40263_, _40215_, _39996_);
  and (_40264_, _40263_, _40262_);
  or (_40265_, _40264_, _40081_);
  or (_40266_, _40255_, _40166_);
  and (_40267_, _40266_, _40115_);
  and (_40268_, _40267_, _40265_);
  or (_40269_, _40268_, _40258_);
  and (_40270_, _40269_, _40104_);
  or (_40271_, _40270_, _40246_);
  and (_42929_, _40271_, _41991_);
  and (_40272_, _40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40273_, _40247_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40274_, _40273_, _40250_);
  or (_40275_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40276_, _40275_, _40203_);
  and (_40277_, _40276_, _40274_);
  or (_40278_, _40277_, _40067_);
  or (_40279_, _40172_, _40005_);
  and (_40280_, _40279_, _40077_);
  and (_40281_, _40280_, _40278_);
  and (_40282_, _40259_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40283_, _40282_, _40261_);
  or (_40284_, _40275_, _40215_);
  and (_40285_, _40284_, _40283_);
  or (_40286_, _40285_, _40081_);
  or (_40287_, _40166_, _40005_);
  and (_40288_, _40287_, _40115_);
  and (_40289_, _40288_, _40286_);
  or (_40290_, _40289_, _40281_);
  and (_40291_, _40290_, _40104_);
  or (_40292_, _40291_, _40272_);
  and (_42931_, _40292_, _41991_);
  and (_40293_, _40096_, _40077_);
  nand (_40294_, _40096_, _40092_);
  and (_40295_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_40296_, _40295_, _40293_);
  and (_42933_, _40296_, _41991_);
  and (_40297_, _40093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_40298_, _40297_, _40078_);
  and (_42935_, _40298_, _41991_);
  and (_40299_, _39983_, _24455_);
  or (_40300_, _40299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40301_, _40300_, _39992_);
  nand (_40302_, _40299_, _28687_);
  and (_40303_, _40302_, _40301_);
  and (_40304_, _39985_, _38608_);
  or (_40305_, _40304_, _40303_);
  and (_42937_, _40305_, _41991_);
  and (_40306_, _39983_, _30720_);
  nand (_40307_, _40306_, _28687_);
  or (_40308_, _40306_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_40309_, _40308_, _39992_);
  and (_40310_, _40309_, _40307_);
  nor (_40311_, _39992_, _38592_);
  or (_40312_, _40311_, _40310_);
  and (_42939_, _40312_, _41991_);
  and (_40313_, _39983_, _32120_);
  nand (_40314_, _40313_, _28687_);
  or (_40315_, _40313_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_40316_, _40315_, _39992_);
  and (_40317_, _40316_, _40314_);
  nor (_40318_, _39992_, _38477_);
  or (_40319_, _40318_, _40317_);
  and (_42941_, _40319_, _41991_);
  and (_40320_, _39970_, _24455_);
  nand (_40321_, _40320_, _28687_);
  or (_40322_, _40320_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40323_, _40322_, _39974_);
  and (_40324_, _40323_, _40321_);
  and (_40325_, _39973_, _38608_);
  or (_40326_, _40325_, _40324_);
  and (_42943_, _40326_, _41991_);
  and (_40327_, _39970_, _30003_);
  nand (_40328_, _40327_, _28687_);
  or (_40329_, _40327_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40330_, _40329_, _39974_);
  and (_40331_, _40330_, _40328_);
  nor (_40332_, _39974_, _38599_);
  or (_40333_, _40332_, _40331_);
  and (_42945_, _40333_, _41991_);
  and (_40334_, _30741_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40335_, _40334_, _30730_);
  and (_40336_, _40335_, _39970_);
  nand (_40337_, _39970_, _39598_);
  and (_40338_, _40337_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40339_, _40338_, _39973_);
  or (_40340_, _40339_, _40336_);
  nand (_40341_, _39973_, _38592_);
  and (_40342_, _40341_, _41991_);
  and (_42947_, _40342_, _40340_);
  and (_40343_, _39970_, _31425_);
  nand (_40344_, _40343_, _28687_);
  or (_40345_, _40343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40346_, _40345_, _39974_);
  and (_40347_, _40346_, _40344_);
  nor (_40348_, _39974_, _38552_);
  or (_40349_, _40348_, _40347_);
  and (_42949_, _40349_, _41991_);
  and (_40350_, _39970_, _32120_);
  nand (_40351_, _40350_, _28687_);
  or (_40352_, _40350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40353_, _40352_, _39974_);
  and (_40354_, _40353_, _40351_);
  nor (_40355_, _39974_, _38477_);
  or (_40356_, _40355_, _40354_);
  and (_42951_, _40356_, _41991_);
  and (_40357_, _39970_, _32930_);
  nand (_40358_, _40357_, _28687_);
  or (_40359_, _40357_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40360_, _40359_, _39974_);
  and (_40361_, _40360_, _40358_);
  nor (_40362_, _39974_, _38402_);
  or (_40363_, _40362_, _40361_);
  and (_42953_, _40363_, _41991_);
  and (_40364_, _39970_, _33652_);
  nand (_40365_, _40364_, _28687_);
  or (_40366_, _40364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40367_, _40366_, _39974_);
  and (_40368_, _40367_, _40365_);
  nor (_40369_, _39974_, _38326_);
  or (_40370_, _40369_, _40368_);
  and (_42954_, _40370_, _41991_);
  and (_40371_, _39948_, _24455_);
  nand (_40372_, _40371_, _28687_);
  or (_40373_, _40371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40374_, _40373_, _39953_);
  and (_40375_, _40374_, _40372_);
  and (_40376_, _39952_, _38608_);
  or (_40377_, _40376_, _40375_);
  and (_42956_, _40377_, _41991_);
  and (_40378_, _39948_, _30003_);
  nand (_40379_, _40378_, _28687_);
  or (_40380_, _40378_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40381_, _40380_, _39953_);
  and (_40382_, _40381_, _40379_);
  nor (_40383_, _39953_, _38599_);
  or (_40384_, _40383_, _40382_);
  and (_42958_, _40384_, _41991_);
  and (_40385_, _30741_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40386_, _40385_, _30730_);
  and (_40387_, _40386_, _39948_);
  nand (_40388_, _39948_, _39598_);
  and (_40389_, _40388_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40390_, _40389_, _39952_);
  or (_40391_, _40390_, _40387_);
  nand (_40392_, _39952_, _38592_);
  and (_40393_, _40392_, _41991_);
  and (_42960_, _40393_, _40391_);
  and (_40394_, _39948_, _31425_);
  nand (_40395_, _40394_, _28687_);
  or (_40396_, _40394_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40397_, _40396_, _39953_);
  and (_40398_, _40397_, _40395_);
  nor (_40399_, _39953_, _38552_);
  or (_40400_, _40399_, _40398_);
  and (_42962_, _40400_, _41991_);
  and (_40401_, _39948_, _32120_);
  nand (_40402_, _40401_, _28687_);
  or (_40403_, _40401_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40404_, _40403_, _39953_);
  and (_40405_, _40404_, _40402_);
  nor (_40406_, _39953_, _38477_);
  or (_40407_, _40406_, _40405_);
  and (_42964_, _40407_, _41991_);
  and (_40408_, _39948_, _32930_);
  nand (_40409_, _40408_, _28687_);
  or (_40410_, _40408_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40411_, _40410_, _39953_);
  and (_40412_, _40411_, _40409_);
  nor (_40413_, _39953_, _38402_);
  or (_40414_, _40413_, _40412_);
  and (_42966_, _40414_, _41991_);
  and (_40415_, _39948_, _33652_);
  nand (_40416_, _40415_, _28687_);
  or (_40417_, _40415_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_40418_, _40417_, _40416_);
  or (_40419_, _40418_, _39952_);
  nand (_40420_, _39952_, _38326_);
  and (_40421_, _40420_, _41991_);
  and (_42968_, _40421_, _40419_);
  nor (_40422_, _24949_, _23920_);
  nor (_40423_, _40422_, _28054_);
  not (_40424_, _40423_);
  not (_40425_, _38625_);
  and (_40426_, _40425_, _37986_);
  not (_40427_, _40426_);
  not (_40428_, _37964_);
  and (_40429_, _40428_, _37563_);
  and (_40430_, _40429_, _36452_);
  not (_40431_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_40432_, _39033_, _40431_);
  nor (_40433_, _40432_, _39094_);
  nor (_40434_, _40433_, _35507_);
  and (_40435_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  not (_40436_, _40435_);
  and (_40437_, _40433_, _36112_);
  and (_40438_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_40439_, _40433_, _36112_);
  and (_40440_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_40441_, _40440_, _40438_);
  and (_40442_, _40441_, _40436_);
  nand (_40443_, _35507_, _29981_);
  or (_40444_, _35507_, _29981_);
  not (_40445_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_40446_, _30741_, _40445_);
  and (_40447_, _40446_, _40423_);
  and (_40448_, _40447_, _40444_);
  and (_40449_, _40448_, _40443_);
  and (_40450_, _40433_, _25113_);
  nor (_40451_, _40433_, _25113_);
  nor (_40452_, _40451_, _40450_);
  and (_40453_, _40452_, _40449_);
  and (_40454_, _40433_, _35507_);
  and (_40455_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_40456_, _40455_, _40453_);
  and (_40457_, _40456_, _40442_);
  and (_40458_, _40453_, _38194_);
  or (_40459_, _40458_, _40457_);
  not (_40460_, _40459_);
  and (_40461_, _40460_, _40430_);
  not (_40462_, _40461_);
  not (_40463_, _36452_);
  nor (_40464_, _40428_, _37563_);
  not (_40465_, _33838_);
  and (_40466_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_40467_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_40468_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_40469_, _40468_, _40467_);
  and (_40470_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_40471_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_40472_, _40471_, _40470_);
  and (_40473_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_40474_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_40475_, _40474_, _40473_);
  and (_40476_, _40475_, _40472_);
  and (_40477_, _40476_, _40469_);
  nor (_40478_, _33904_, _40465_);
  not (_40479_, _40478_);
  nor (_40480_, _40479_, _40477_);
  nor (_40481_, _40480_, _40466_);
  not (_40482_, _40481_);
  and (_40483_, _40482_, _40464_);
  nor (_40484_, _40483_, _40463_);
  and (_40485_, _40484_, _40462_);
  and (_40486_, _40485_, _40427_);
  not (_40487_, _36638_);
  and (_40488_, _37220_, _40487_);
  nor (_40489_, _37154_, _37088_);
  nor (_40490_, _37055_, _36814_);
  and (_40491_, _40490_, _40489_);
  and (_40492_, _37350_, _36934_);
  and (_40493_, _40492_, _40491_);
  and (_40494_, _40493_, _40488_);
  nor (_40495_, _40494_, _35564_);
  and (_40496_, _36891_, _35530_);
  nor (_40497_, _37471_, _40496_);
  nor (_40498_, _37493_, _40497_);
  nor (_40499_, _40498_, _40495_);
  not (_40500_, _40499_);
  and (_40501_, _40500_, _40486_);
  not (_40502_, _38651_);
  and (_40503_, _40502_, _37986_);
  and (_40504_, _40464_, _36452_);
  and (_40505_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_40506_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_40507_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_40508_, _40507_, _40506_);
  and (_40509_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_40510_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_40511_, _40510_, _40509_);
  and (_40512_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_40513_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_40514_, _40513_, _40512_);
  and (_40515_, _40514_, _40511_);
  and (_40516_, _40515_, _40508_);
  nor (_40517_, _40516_, _40479_);
  nor (_40518_, _40517_, _40505_);
  not (_40519_, _40518_);
  and (_40520_, _40519_, _40504_);
  nor (_40521_, _40520_, _40503_);
  not (_40522_, _40433_);
  and (_40523_, _37964_, _37563_);
  and (_40524_, _40523_, _36452_);
  and (_40525_, _40524_, _40522_);
  and (_40526_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  not (_40527_, _40526_);
  and (_40528_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_40529_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_40530_, _40529_, _40528_);
  and (_40531_, _40530_, _40527_);
  and (_40532_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_40533_, _40532_, _40453_);
  and (_40534_, _40533_, _40531_);
  and (_40535_, _40453_, _38552_);
  or (_40536_, _40535_, _40534_);
  not (_40537_, _40536_);
  and (_40538_, _40537_, _40430_);
  nor (_40539_, _40538_, _40525_);
  and (_40540_, _40539_, _40521_);
  not (_40541_, _40540_);
  and (_40542_, _40541_, _40501_);
  and (_40543_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_40544_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_40545_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_40546_, _40545_, _40544_);
  and (_40547_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_40548_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_40549_, _40548_, _40547_);
  and (_40550_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_40551_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_40552_, _40551_, _40550_);
  and (_40553_, _40552_, _40549_);
  and (_40554_, _40553_, _40546_);
  nor (_40555_, _40554_, _40479_);
  nor (_40556_, _40555_, _40543_);
  not (_40557_, _40556_);
  and (_40558_, _40557_, _40504_);
  and (_40559_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  not (_40560_, _40559_);
  and (_40561_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_40562_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_40563_, _40562_, _40561_);
  and (_40564_, _40563_, _40560_);
  and (_40565_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_40566_, _40565_, _40453_);
  and (_40567_, _40566_, _40564_);
  and (_40568_, _40453_, _38607_);
  or (_40569_, _40568_, _40567_);
  not (_40570_, _40569_);
  and (_40571_, _40570_, _40430_);
  nor (_40572_, _40571_, _40558_);
  not (_40573_, _38633_);
  and (_40574_, _40573_, _37986_);
  and (_40575_, _40524_, _36112_);
  nor (_40576_, _40575_, _40574_);
  and (_40577_, _40576_, _40572_);
  nor (_40578_, _40577_, _40500_);
  nor (_40579_, _40578_, _40542_);
  and (_40580_, _24949_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_40581_, _40580_, _25113_);
  nor (_40582_, _24433_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40583_, _40582_, _40581_);
  not (_40584_, _40583_);
  and (_40585_, _40584_, _40579_);
  nor (_40586_, _40585_, _40424_);
  not (_40587_, _38402_);
  and (_40588_, _40453_, _40587_);
  and (_40589_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_40590_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_40591_, _40590_, _40589_);
  and (_40592_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_40593_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_40594_, _40593_, _40592_);
  and (_40595_, _40594_, _40591_);
  nor (_40596_, _40595_, _40453_);
  nor (_40597_, _40596_, _40588_);
  not (_40598_, _40597_);
  and (_40599_, _40598_, _40430_);
  not (_40600_, _40599_);
  and (_40601_, _40463_, _37964_);
  and (_40602_, _40601_, _37563_);
  not (_40603_, _38663_);
  and (_40604_, _40603_, _37986_);
  nor (_40605_, _40604_, _40602_);
  and (_40606_, _40605_, _40600_);
  and (_40607_, _37975_, _40463_);
  and (_40608_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_40609_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_40610_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_40611_, _40610_, _40609_);
  and (_40612_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_40613_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_40614_, _40613_, _40612_);
  and (_40615_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_40616_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_40617_, _40616_, _40615_);
  and (_40618_, _40617_, _40614_);
  and (_40619_, _40618_, _40611_);
  nor (_40620_, _40619_, _40479_);
  nor (_40621_, _40620_, _40608_);
  not (_40622_, _40621_);
  and (_40623_, _40622_, _40504_);
  nor (_40624_, _40623_, _40607_);
  and (_40625_, _40624_, _40606_);
  not (_40626_, _40625_);
  and (_40627_, _40626_, _40501_);
  and (_40628_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_40629_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_40630_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_40631_, _40630_, _40629_);
  and (_40632_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_40633_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_40634_, _40633_, _40632_);
  and (_40635_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_40636_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_40637_, _40636_, _40635_);
  and (_40638_, _40637_, _40634_);
  and (_40639_, _40638_, _40631_);
  nor (_40640_, _40639_, _40479_);
  nor (_40641_, _40640_, _40628_);
  not (_40642_, _40641_);
  and (_40643_, _40642_, _40504_);
  and (_40644_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  not (_40645_, _40644_);
  and (_40646_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_40647_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_40648_, _40647_, _40646_);
  and (_40649_, _40648_, _40645_);
  and (_40650_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_40651_, _40650_, _40453_);
  and (_40652_, _40651_, _40649_);
  and (_40653_, _40453_, _38592_);
  or (_40654_, _40653_, _40652_);
  not (_40655_, _40654_);
  and (_40656_, _40655_, _40430_);
  nor (_40657_, _40656_, _40643_);
  not (_40658_, _38645_);
  and (_40659_, _40658_, _37986_);
  and (_40660_, _40524_, _36310_);
  nor (_40661_, _40660_, _40659_);
  and (_40662_, _40661_, _40657_);
  nor (_40663_, _40662_, _40500_);
  nor (_40664_, _40663_, _40627_);
  and (_40665_, _40580_, _39202_);
  nor (_40666_, _24197_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40667_, _40666_, _40665_);
  not (_40668_, _40667_);
  and (_40669_, _40668_, _40664_);
  nor (_40670_, _40584_, _40579_);
  nor (_40671_, _40670_, _40669_);
  and (_40672_, _40671_, _40586_);
  and (_40673_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_40674_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_40675_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_40676_, _40675_, _40674_);
  and (_40677_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_40678_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_40679_, _40678_, _40677_);
  and (_40680_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_40681_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_40682_, _40681_, _40680_);
  and (_40683_, _40682_, _40679_);
  and (_40684_, _40683_, _40676_);
  nor (_40685_, _40684_, _40479_);
  nor (_40686_, _40685_, _40673_);
  not (_40687_, _40686_);
  and (_40688_, _40687_, _40504_);
  not (_40689_, _39134_);
  and (_40690_, _40524_, _40689_);
  nor (_40691_, _40690_, _40688_);
  not (_40692_, _38477_);
  and (_40693_, _40453_, _40692_);
  and (_40694_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_40695_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_40696_, _40695_, _40694_);
  and (_40697_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_40698_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_40699_, _40698_, _40697_);
  and (_40700_, _40699_, _40696_);
  nor (_40701_, _40700_, _40453_);
  nor (_40702_, _40701_, _40693_);
  not (_40703_, _40702_);
  and (_40704_, _40703_, _40430_);
  not (_40705_, _40704_);
  not (_40706_, _38657_);
  and (_40707_, _40706_, _37986_);
  nor (_40708_, _40707_, _40601_);
  and (_40709_, _40708_, _40705_);
  and (_40710_, _40709_, _40691_);
  not (_40711_, _40710_);
  and (_40712_, _40711_, _40501_);
  and (_40713_, _40429_, _40463_);
  and (_40714_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_40715_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_40716_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_40717_, _40716_, _40715_);
  and (_40718_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_40719_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_40720_, _40719_, _40718_);
  and (_40721_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_40722_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_40723_, _40722_, _40721_);
  and (_40724_, _40723_, _40720_);
  and (_40725_, _40724_, _40717_);
  nor (_40726_, _40725_, _40479_);
  nor (_40727_, _40726_, _40714_);
  not (_40728_, _40727_);
  and (_40729_, _40728_, _40504_);
  nor (_40730_, _40729_, _40713_);
  not (_40731_, _38639_);
  and (_40732_, _40731_, _37986_);
  and (_40733_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_40734_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_40735_, _40734_, _40733_);
  and (_40736_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_40737_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_40738_, _40737_, _40736_);
  and (_40739_, _40738_, _40735_);
  nor (_40740_, _40739_, _40453_);
  not (_40741_, _38599_);
  and (_40742_, _40453_, _40741_);
  nor (_40743_, _40742_, _40740_);
  not (_40749_, _40743_);
  and (_40755_, _40749_, _40430_);
  and (_40761_, _40524_, _36123_);
  or (_40767_, _40761_, _40755_);
  nor (_40773_, _40767_, _40732_);
  and (_40776_, _40773_, _40730_);
  nor (_40777_, _40776_, _40500_);
  nor (_40778_, _40777_, _40712_);
  not (_40779_, _25276_);
  and (_40780_, _40580_, _40779_);
  nor (_40781_, _24312_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_40782_, _40781_, _40780_);
  nand (_40783_, _40782_, _40778_);
  or (_40784_, _40782_, _40778_);
  and (_40785_, _40784_, _40783_);
  not (_40786_, _40785_);
  nor (_40787_, _40668_, _40664_);
  not (_40788_, _40787_);
  not (_40789_, _38669_);
  and (_40791_, _40789_, _37986_);
  and (_40794_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_40798_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_40801_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_40802_, _40801_, _40798_);
  and (_40803_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_40805_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_40811_, _40805_, _40803_);
  and (_40814_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_40815_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_40816_, _40815_, _40814_);
  and (_40820_, _40816_, _40811_);
  and (_40826_, _40820_, _40802_);
  nor (_40827_, _40826_, _40479_);
  nor (_40828_, _40827_, _40794_);
  not (_40830_, _40828_);
  and (_40836_, _40830_, _40464_);
  nor (_40839_, _40836_, _40791_);
  nor (_40840_, _40429_, _36452_);
  not (_40841_, _38326_);
  and (_40845_, _40453_, _40841_);
  and (_40851_, _40437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_40852_, _40439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_40853_, _40852_, _40851_);
  and (_40856_, _40434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_40862_, _40454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_40864_, _40862_, _40856_);
  and (_40865_, _40864_, _40853_);
  nor (_40868_, _40865_, _40453_);
  nor (_40874_, _40868_, _40845_);
  not (_40876_, _40874_);
  and (_40877_, _40876_, _40430_);
  nor (_40879_, _40877_, _40840_);
  and (_40885_, _40879_, _40839_);
  and (_40888_, _40885_, _40501_);
  nor (_40889_, _40541_, _40501_);
  nor (_40890_, _40889_, _40888_);
  nor (_40894_, _40580_, _25113_);
  and (_40900_, _40580_, _24665_);
  nor (_40901_, _40900_, _40894_);
  not (_40902_, _40901_);
  and (_40905_, _40902_, _40890_);
  nor (_40911_, _40902_, _40890_);
  nor (_40913_, _40911_, _40905_);
  and (_40914_, _40913_, _40788_);
  and (_40917_, _40914_, _40786_);
  and (_40923_, _40917_, _40672_);
  not (_40925_, _40664_);
  and (_40926_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_40928_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_40934_, _40579_, _40928_);
  or (_40937_, _40934_, _40926_);
  and (_40938_, _40937_, _40778_);
  not (_40939_, _40778_);
  not (_40945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_40949_, _40579_, _40945_);
  and (_40950_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_40951_, _40950_, _40949_);
  and (_40956_, _40951_, _40939_);
  or (_40961_, _40956_, _40938_);
  or (_40962_, _40961_, _40925_);
  not (_40963_, _40890_);
  and (_40968_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_40973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_40974_, _40579_, _40973_);
  or (_40975_, _40974_, _40968_);
  and (_40980_, _40975_, _40778_);
  not (_40984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_40985_, _40579_, _40984_);
  and (_40986_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_40987_, _40986_, _40985_);
  and (_40988_, _40987_, _40939_);
  or (_40989_, _40988_, _40980_);
  or (_40990_, _40989_, _40664_);
  and (_40991_, _40990_, _40963_);
  and (_40992_, _40991_, _40962_);
  not (_40993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_40994_, _40579_, _40993_);
  or (_40995_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_40996_, _40995_, _40994_);
  and (_40997_, _40996_, _40778_);
  or (_40998_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_40999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_41000_, _40579_, _40999_);
  and (_41001_, _41000_, _40998_);
  and (_41002_, _41001_, _40939_);
  or (_41003_, _41002_, _40997_);
  or (_41004_, _41003_, _40925_);
  not (_41005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_41006_, _40579_, _41005_);
  or (_41007_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_41008_, _41007_, _41006_);
  and (_41009_, _41008_, _40778_);
  or (_41010_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_41011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_41012_, _40579_, _41011_);
  and (_41013_, _41012_, _41010_);
  and (_41014_, _41013_, _40939_);
  or (_41015_, _41014_, _41009_);
  or (_41016_, _41015_, _40664_);
  and (_41017_, _41016_, _40890_);
  and (_41018_, _41017_, _41004_);
  or (_41019_, _41018_, _40992_);
  or (_41020_, _41019_, _40923_);
  not (_41021_, _40923_);
  or (_41022_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_41023_, _41022_, _41991_);
  and (_43047_, _41023_, _41020_);
  nor (_41024_, _40583_, _40424_);
  nor (_41025_, _40782_, _40424_);
  and (_41026_, _41025_, _41024_);
  and (_41027_, _40901_, _40423_);
  nor (_41028_, _40667_, _40424_);
  and (_41029_, _41028_, _41027_);
  and (_41030_, _41029_, _41026_);
  and (_41031_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_41032_, _41031_, _26104_);
  nor (_41033_, _41032_, _28687_);
  nor (_41034_, _38194_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41035_, _26104_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41036_, _17464_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41037_, _41036_, _41035_);
  or (_41038_, _41037_, _41034_);
  or (_41039_, _41038_, _41033_);
  and (_41040_, _41039_, _40423_);
  and (_41041_, _41040_, _41030_);
  not (_41042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_41043_, _41030_, _41042_);
  or (_43059_, _41043_, _41041_);
  nor (_41044_, _41028_, _41027_);
  nor (_41045_, _41025_, _41024_);
  and (_41046_, _41045_, _40423_);
  and (_41047_, _41046_, _41044_);
  and (_41048_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _26093_);
  and (_41049_, _41048_, _26137_);
  not (_41050_, _41049_);
  nor (_41051_, _41050_, _28687_);
  not (_41052_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41053_, _38607_, _41052_);
  or (_41054_, _16303_, _41052_);
  and (_41055_, _41054_, _41050_);
  and (_41056_, _41055_, _41053_);
  or (_41057_, _41056_, _41051_);
  and (_41058_, _41057_, _41047_);
  not (_41059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_41060_, _41047_, _41059_);
  or (_43315_, _41060_, _41058_);
  not (_41061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_41062_, _41047_, _41061_);
  nand (_41063_, _41048_, _26190_);
  nor (_41064_, _41063_, _28687_);
  nor (_41065_, _38599_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41066_, _41048_, _26202_);
  and (_41067_, _41048_, _26104_);
  or (_41068_, _41067_, _41031_);
  or (_41069_, _41068_, _41066_);
  and (_41070_, _41069_, _17290_);
  or (_41071_, _41070_, _41065_);
  or (_41072_, _41071_, _41064_);
  and (_41073_, _41072_, _41047_);
  or (_43321_, _41073_, _41062_);
  not (_41074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_41075_, _41047_, _41074_);
  nand (_41076_, _41048_, _26213_);
  nor (_41077_, _41076_, _28687_);
  nor (_41078_, _38592_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41079_, _41048_, _26170_);
  or (_41080_, _41079_, _41068_);
  and (_41081_, _41080_, _15941_);
  or (_41082_, _41081_, _41078_);
  or (_41083_, _41082_, _41077_);
  and (_41084_, _41083_, _41047_);
  or (_43327_, _41084_, _41075_);
  not (_41085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_41086_, _41047_, _41085_);
  and (_41087_, _41067_, _29308_);
  nor (_41088_, _38552_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_41089_, _41066_, _41031_);
  or (_41090_, _41089_, _41079_);
  and (_41091_, _41090_, _16973_);
  or (_41092_, _41091_, _41088_);
  or (_41093_, _41092_, _41087_);
  and (_41094_, _41093_, _41047_);
  or (_43333_, _41094_, _41086_);
  nand (_41095_, _41031_, _26137_);
  nor (_41096_, _41095_, _28687_);
  nor (_41097_, _38477_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41098_, _26137_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41099_, _16139_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41100_, _41099_, _41098_);
  or (_41101_, _41100_, _41097_);
  or (_41102_, _41101_, _41096_);
  and (_41103_, _41102_, _41047_);
  not (_41104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41105_, _41047_, _41104_);
  or (_43339_, _41105_, _41103_);
  nand (_41106_, _41031_, _26190_);
  nor (_41107_, _41106_, _28687_);
  nor (_41108_, _38402_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41109_, _26190_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41110_, _17127_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41111_, _41110_, _41109_);
  or (_41112_, _41111_, _41108_);
  or (_41113_, _41112_, _41107_);
  and (_41114_, _41113_, _41047_);
  not (_41115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41116_, _41047_, _41115_);
  or (_43345_, _41116_, _41114_);
  nand (_41117_, _41031_, _26213_);
  nor (_41118_, _41117_, _28687_);
  nor (_41119_, _38326_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_41120_, _26213_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_41121_, _16479_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41122_, _41121_, _41120_);
  or (_41123_, _41122_, _41119_);
  or (_41124_, _41123_, _41118_);
  and (_41125_, _41124_, _41047_);
  not (_41126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_41127_, _41047_, _41126_);
  or (_43348_, _41127_, _41125_);
  and (_41128_, _41047_, _41039_);
  not (_41129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_41130_, _41047_, _41129_);
  or (_43351_, _41130_, _41128_);
  and (_41131_, _41057_, _40423_);
  and (_41132_, _41024_, _40782_);
  and (_41133_, _41132_, _41044_);
  and (_41134_, _41133_, _41131_);
  not (_41135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_41136_, _41133_, _41135_);
  or (_43359_, _41136_, _41134_);
  and (_41137_, _41072_, _40423_);
  and (_41138_, _41133_, _41137_);
  not (_41139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_41140_, _41133_, _41139_);
  or (_43363_, _41140_, _41138_);
  and (_41141_, _41083_, _40423_);
  and (_41142_, _41133_, _41141_);
  not (_41143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_41144_, _41133_, _41143_);
  or (_43367_, _41144_, _41142_);
  and (_41145_, _41093_, _40423_);
  and (_41146_, _41133_, _41145_);
  not (_41147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_41148_, _41133_, _41147_);
  or (_43371_, _41148_, _41146_);
  and (_41149_, _41102_, _40423_);
  and (_41150_, _41133_, _41149_);
  not (_41151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_41152_, _41133_, _41151_);
  or (_43375_, _41152_, _41150_);
  and (_41153_, _41113_, _40423_);
  and (_41154_, _41133_, _41153_);
  not (_41155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_41156_, _41133_, _41155_);
  or (_43379_, _41156_, _41154_);
  and (_41157_, _41124_, _40423_);
  and (_41158_, _41133_, _41157_);
  not (_41159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_41160_, _41133_, _41159_);
  or (_43383_, _41160_, _41158_);
  and (_41161_, _41133_, _41040_);
  nor (_41162_, _41133_, _40928_);
  or (_43386_, _41162_, _41161_);
  and (_41163_, _41025_, _40583_);
  and (_41164_, _41163_, _41044_);
  and (_41165_, _41164_, _41131_);
  not (_41166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_41167_, _41164_, _41166_);
  or (_43394_, _41167_, _41165_);
  and (_41168_, _41164_, _41137_);
  not (_41169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_41170_, _41164_, _41169_);
  or (_43398_, _41170_, _41168_);
  and (_41171_, _41164_, _41141_);
  not (_41172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_41173_, _41164_, _41172_);
  or (_43402_, _41173_, _41171_);
  and (_41174_, _41164_, _41145_);
  not (_41175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_41176_, _41164_, _41175_);
  or (_43406_, _41176_, _41174_);
  and (_41177_, _41164_, _41149_);
  not (_41178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_41179_, _41164_, _41178_);
  or (_43410_, _41179_, _41177_);
  and (_41180_, _41164_, _41153_);
  not (_41181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_41182_, _41164_, _41181_);
  or (_43414_, _41182_, _41180_);
  and (_41183_, _41164_, _41157_);
  not (_41184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_41185_, _41164_, _41184_);
  or (_43418_, _41185_, _41183_);
  and (_41186_, _41164_, _41040_);
  not (_41187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_41188_, _41164_, _41187_);
  or (_43421_, _41188_, _41186_);
  and (_41189_, _41044_, _41026_);
  and (_41190_, _41189_, _41131_);
  not (_41191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_41192_, _41189_, _41191_);
  or (_43446_, _41192_, _41190_);
  and (_41193_, _41189_, _41137_);
  not (_41194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_41195_, _41189_, _41194_);
  or (_43466_, _41195_, _41193_);
  and (_41196_, _41189_, _41141_);
  not (_41197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_41198_, _41189_, _41197_);
  or (_43484_, _41198_, _41196_);
  and (_41199_, _41189_, _41145_);
  not (_41200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_41201_, _41189_, _41200_);
  or (_43502_, _41201_, _41199_);
  and (_41202_, _41189_, _41149_);
  not (_41203_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_41204_, _41189_, _41203_);
  or (_43520_, _41204_, _41202_);
  and (_41205_, _41189_, _41153_);
  not (_41206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_41207_, _41189_, _41206_);
  or (_43539_, _41207_, _41205_);
  and (_41208_, _41189_, _41157_);
  not (_41209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_41210_, _41189_, _41209_);
  or (_43559_, _41210_, _41208_);
  and (_41211_, _41189_, _41040_);
  nor (_41212_, _41189_, _40945_);
  or (_43573_, _41212_, _41211_);
  and (_41213_, _41028_, _40902_);
  and (_41214_, _41213_, _41045_);
  and (_41215_, _41214_, _41131_);
  not (_41216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_41217_, _41214_, _41216_);
  or (_43610_, _41217_, _41215_);
  and (_41218_, _41214_, _41137_);
  not (_41219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_41220_, _41214_, _41219_);
  or (_43635_, _41220_, _41218_);
  and (_41221_, _41214_, _41141_);
  not (_41222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_41223_, _41214_, _41222_);
  or (_43653_, _41223_, _41221_);
  and (_41224_, _41214_, _41145_);
  not (_41225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_41226_, _41214_, _41225_);
  or (_43664_, _41226_, _41224_);
  and (_41227_, _41214_, _41149_);
  not (_41228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41229_, _41214_, _41228_);
  or (_43668_, _41229_, _41227_);
  and (_41230_, _41214_, _41153_);
  not (_41231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41232_, _41214_, _41231_);
  or (_43672_, _41232_, _41230_);
  and (_41233_, _41214_, _41157_);
  not (_41234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41235_, _41214_, _41234_);
  or (_43676_, _41235_, _41233_);
  and (_41236_, _41214_, _41040_);
  not (_41237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_41238_, _41214_, _41237_);
  or (_43679_, _41238_, _41236_);
  and (_41239_, _41213_, _41132_);
  and (_41240_, _41239_, _41131_);
  not (_41241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_41242_, _41239_, _41241_);
  or (_43684_, _41242_, _41240_);
  and (_41243_, _41239_, _41137_);
  not (_41244_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_41245_, _41239_, _41244_);
  or (_43688_, _41245_, _41243_);
  and (_41246_, _41239_, _41141_);
  not (_41247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_41248_, _41239_, _41247_);
  or (_43692_, _41248_, _41246_);
  and (_41249_, _41239_, _41145_);
  not (_41250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_41251_, _41239_, _41250_);
  or (_43696_, _41251_, _41249_);
  and (_41252_, _41239_, _41149_);
  not (_41253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_41254_, _41239_, _41253_);
  or (_43700_, _41254_, _41252_);
  and (_41255_, _41239_, _41153_);
  not (_41256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_41257_, _41239_, _41256_);
  or (_43704_, _41257_, _41255_);
  and (_41258_, _41239_, _41157_);
  not (_41259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_41260_, _41239_, _41259_);
  or (_43708_, _41260_, _41258_);
  and (_41261_, _41239_, _41040_);
  nor (_41262_, _41239_, _40973_);
  or (_43711_, _41262_, _41261_);
  and (_41263_, _41213_, _41163_);
  and (_41264_, _41263_, _41131_);
  not (_41265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_41266_, _41263_, _41265_);
  or (_43716_, _41266_, _41264_);
  and (_41267_, _41263_, _41137_);
  not (_41268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_41269_, _41263_, _41268_);
  or (_43720_, _41269_, _41267_);
  and (_41270_, _41263_, _41141_);
  not (_41271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_41272_, _41263_, _41271_);
  or (_43724_, _41272_, _41270_);
  and (_41273_, _41263_, _41145_);
  not (_41274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_41275_, _41263_, _41274_);
  or (_43728_, _41275_, _41273_);
  and (_41276_, _41263_, _41149_);
  not (_41277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_41278_, _41263_, _41277_);
  or (_43732_, _41278_, _41276_);
  and (_41279_, _41263_, _41153_);
  not (_41280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_41281_, _41263_, _41280_);
  or (_43736_, _41281_, _41279_);
  and (_41282_, _41263_, _41157_);
  not (_41283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_41284_, _41263_, _41283_);
  or (_43740_, _41284_, _41282_);
  and (_41285_, _41263_, _41040_);
  not (_41286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_41287_, _41263_, _41286_);
  or (_43743_, _41287_, _41285_);
  and (_41288_, _41213_, _41026_);
  and (_41289_, _41288_, _41131_);
  not (_41290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_41291_, _41288_, _41290_);
  or (_43748_, _41291_, _41289_);
  and (_41292_, _41288_, _41137_);
  not (_41293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_41294_, _41288_, _41293_);
  or (_43752_, _41294_, _41292_);
  and (_41295_, _41288_, _41141_);
  not (_41296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_41297_, _41288_, _41296_);
  or (_43756_, _41297_, _41295_);
  and (_41298_, _41288_, _41145_);
  not (_41299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_41300_, _41288_, _41299_);
  or (_43760_, _41300_, _41298_);
  and (_41301_, _41288_, _41149_);
  not (_41302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_41303_, _41288_, _41302_);
  or (_43764_, _41303_, _41301_);
  and (_41304_, _41288_, _41153_);
  not (_41305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_41306_, _41288_, _41305_);
  or (_43767_, _41306_, _41304_);
  and (_41307_, _41288_, _41157_);
  not (_41308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_41309_, _41288_, _41308_);
  or (_43771_, _41309_, _41307_);
  and (_41310_, _41288_, _41040_);
  nor (_41311_, _41288_, _40984_);
  or (_43774_, _41311_, _41310_);
  and (_41312_, _41027_, _40667_);
  and (_41313_, _41312_, _41045_);
  and (_41314_, _41313_, _41131_);
  not (_41315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_41316_, _41313_, _41315_);
  or (_43782_, _41316_, _41314_);
  and (_41317_, _41313_, _41137_);
  not (_41318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_41319_, _41313_, _41318_);
  or (_43786_, _41319_, _41317_);
  and (_41320_, _41313_, _41141_);
  not (_41321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_41322_, _41313_, _41321_);
  or (_43790_, _41322_, _41320_);
  and (_41323_, _41313_, _41145_);
  not (_41324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_41325_, _41313_, _41324_);
  or (_43794_, _41325_, _41323_);
  and (_41326_, _41313_, _41149_);
  not (_41327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_41328_, _41313_, _41327_);
  or (_43798_, _41328_, _41326_);
  and (_41329_, _41313_, _41153_);
  not (_41330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_41331_, _41313_, _41330_);
  or (_43802_, _41331_, _41329_);
  and (_41332_, _41313_, _41157_);
  not (_41333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_41334_, _41313_, _41333_);
  or (_43806_, _41334_, _41332_);
  and (_41335_, _41313_, _41040_);
  nor (_41336_, _41313_, _40993_);
  or (_43809_, _41336_, _41335_);
  and (_41337_, _41312_, _41132_);
  and (_41338_, _41337_, _41131_);
  not (_41339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_41340_, _41337_, _41339_);
  or (_43814_, _41340_, _41338_);
  and (_41341_, _41337_, _41137_);
  not (_41342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_41343_, _41337_, _41342_);
  or (_43818_, _41343_, _41341_);
  and (_41344_, _41337_, _41141_);
  not (_41345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_41346_, _41337_, _41345_);
  or (_43822_, _41346_, _41344_);
  and (_41347_, _41337_, _41145_);
  not (_41348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_41349_, _41337_, _41348_);
  or (_43826_, _41349_, _41347_);
  and (_41350_, _41337_, _41149_);
  not (_41351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_41352_, _41337_, _41351_);
  or (_43830_, _41352_, _41350_);
  and (_41353_, _41337_, _41153_);
  not (_41354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_41355_, _41337_, _41354_);
  or (_43834_, _41355_, _41353_);
  and (_41356_, _41337_, _41157_);
  not (_41357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_41358_, _41337_, _41357_);
  or (_43838_, _41358_, _41356_);
  and (_41359_, _41337_, _41040_);
  not (_41360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_41361_, _41337_, _41360_);
  or (_43841_, _41361_, _41359_);
  and (_41362_, _41312_, _41163_);
  and (_41363_, _41362_, _41131_);
  not (_41364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_41365_, _41362_, _41364_);
  or (_43846_, _41365_, _41363_);
  and (_41366_, _41362_, _41137_);
  not (_41367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_41368_, _41362_, _41367_);
  or (_43850_, _41368_, _41366_);
  and (_41369_, _41362_, _41141_);
  not (_41370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_41371_, _41362_, _41370_);
  or (_43854_, _41371_, _41369_);
  and (_41372_, _41362_, _41145_);
  not (_41373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_41374_, _41362_, _41373_);
  or (_43858_, _41374_, _41372_);
  and (_41375_, _41362_, _41149_);
  not (_41376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_41377_, _41362_, _41376_);
  or (_43862_, _41377_, _41375_);
  and (_41378_, _41362_, _41153_);
  not (_41379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_41380_, _41362_, _41379_);
  or (_43866_, _41380_, _41378_);
  and (_41381_, _41362_, _41157_);
  not (_41382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_41383_, _41362_, _41382_);
  or (_43870_, _41383_, _41381_);
  and (_41384_, _41362_, _41040_);
  nor (_41385_, _41362_, _40999_);
  or (_43873_, _41385_, _41384_);
  and (_41386_, _41312_, _41026_);
  and (_41387_, _41386_, _41131_);
  not (_41388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_41389_, _41386_, _41388_);
  or (_43878_, _41389_, _41387_);
  and (_41390_, _41386_, _41137_);
  not (_41391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_41392_, _41386_, _41391_);
  or (_43882_, _41392_, _41390_);
  and (_41395_, _41386_, _41141_);
  not (_41397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_41399_, _41386_, _41397_);
  or (_43886_, _41399_, _41395_);
  and (_41402_, _41386_, _41145_);
  not (_41404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_41406_, _41386_, _41404_);
  or (_43890_, _41406_, _41402_);
  and (_41409_, _41386_, _41149_);
  not (_41411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_41413_, _41386_, _41411_);
  or (_43894_, _41413_, _41409_);
  and (_41416_, _41386_, _41153_);
  not (_41418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_41420_, _41386_, _41418_);
  or (_43898_, _41420_, _41416_);
  and (_41423_, _41386_, _41157_);
  not (_41425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_41427_, _41386_, _41425_);
  or (_43902_, _41427_, _41423_);
  and (_41430_, _41386_, _41040_);
  not (_41432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_41434_, _41386_, _41432_);
  or (_43905_, _41434_, _41430_);
  and (_41437_, _41045_, _41029_);
  and (_41439_, _41437_, _41131_);
  not (_41441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_41442_, _41437_, _41441_);
  or (_43911_, _41442_, _41439_);
  and (_41443_, _41437_, _41137_);
  not (_41444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_41445_, _41437_, _41444_);
  or (_43915_, _41445_, _41443_);
  and (_41446_, _41437_, _41141_);
  not (_41447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_41448_, _41437_, _41447_);
  or (_43919_, _41448_, _41446_);
  and (_41449_, _41437_, _41145_);
  not (_41450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_41451_, _41437_, _41450_);
  or (_43923_, _41451_, _41449_);
  and (_41452_, _41437_, _41149_);
  not (_41453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_41454_, _41437_, _41453_);
  or (_43927_, _41454_, _41452_);
  and (_41455_, _41437_, _41153_);
  not (_41456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_41457_, _41437_, _41456_);
  or (_43931_, _41457_, _41455_);
  and (_41458_, _41437_, _41157_);
  not (_41459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_41460_, _41437_, _41459_);
  or (_43935_, _41460_, _41458_);
  and (_41461_, _41437_, _41040_);
  nor (_41462_, _41437_, _41005_);
  or (_43938_, _41462_, _41461_);
  and (_41463_, _41132_, _41029_);
  and (_41464_, _41463_, _41131_);
  not (_41465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_41466_, _41463_, _41465_);
  or (_43943_, _41466_, _41464_);
  and (_41467_, _41463_, _41137_);
  not (_41468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_41469_, _41463_, _41468_);
  or (_43947_, _41469_, _41467_);
  and (_41470_, _41463_, _41141_);
  not (_41471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_41472_, _41463_, _41471_);
  or (_43951_, _41472_, _41470_);
  and (_41473_, _41463_, _41145_);
  not (_41474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_41475_, _41463_, _41474_);
  or (_43955_, _41475_, _41473_);
  and (_41476_, _41463_, _41149_);
  not (_41477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_41478_, _41463_, _41477_);
  or (_43959_, _41478_, _41476_);
  and (_41479_, _41463_, _41153_);
  not (_41480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_41481_, _41463_, _41480_);
  or (_43963_, _41481_, _41479_);
  and (_41482_, _41463_, _41157_);
  not (_41483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_41484_, _41463_, _41483_);
  or (_43967_, _41484_, _41482_);
  and (_41485_, _41463_, _41040_);
  not (_41486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_41487_, _41463_, _41486_);
  or (_43970_, _41487_, _41485_);
  and (_41488_, _41163_, _41029_);
  and (_41489_, _41488_, _41131_);
  not (_41490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_41491_, _41488_, _41490_);
  or (_43975_, _41491_, _41489_);
  and (_41492_, _41488_, _41137_);
  not (_41493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_41494_, _41488_, _41493_);
  or (_43979_, _41494_, _41492_);
  and (_41495_, _41488_, _41141_);
  not (_41496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_41497_, _41488_, _41496_);
  or (_43983_, _41497_, _41495_);
  and (_41498_, _41488_, _41145_);
  not (_41499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_41500_, _41488_, _41499_);
  or (_43987_, _41500_, _41498_);
  and (_41501_, _41488_, _41149_);
  not (_41502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_41503_, _41488_, _41502_);
  or (_43991_, _41503_, _41501_);
  and (_41504_, _41488_, _41153_);
  not (_41505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_41506_, _41488_, _41505_);
  or (_43995_, _41506_, _41504_);
  and (_41507_, _41488_, _41157_);
  not (_41508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_41509_, _41488_, _41508_);
  or (_43999_, _41509_, _41507_);
  and (_41510_, _41488_, _41040_);
  nor (_41511_, _41488_, _41011_);
  or (_44002_, _41511_, _41510_);
  and (_41512_, _41131_, _41030_);
  not (_41513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_41514_, _41030_, _41513_);
  or (_44007_, _41514_, _41512_);
  and (_41515_, _41137_, _41030_);
  not (_41516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_41517_, _41030_, _41516_);
  or (_44011_, _41517_, _41515_);
  and (_41518_, _41141_, _41030_);
  not (_41519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_41520_, _41030_, _41519_);
  or (_44015_, _41520_, _41518_);
  and (_41521_, _41145_, _41030_);
  not (_41522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_41523_, _41030_, _41522_);
  or (_44019_, _41523_, _41521_);
  and (_41524_, _41149_, _41030_);
  not (_41525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_41526_, _41030_, _41525_);
  or (_44023_, _41526_, _41524_);
  and (_41527_, _41153_, _41030_);
  not (_41528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_41529_, _41030_, _41528_);
  or (_44027_, _41529_, _41527_);
  and (_41530_, _41157_, _41030_);
  not (_41531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_41532_, _41030_, _41531_);
  or (_44031_, _41532_, _41530_);
  and (_41533_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_41534_, _40579_, _41135_);
  or (_41535_, _41534_, _41533_);
  and (_41536_, _41535_, _40778_);
  nor (_41537_, _40579_, _41191_);
  and (_41538_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_41539_, _41538_, _41537_);
  and (_41540_, _41539_, _40939_);
  or (_41541_, _41540_, _41536_);
  or (_41542_, _41541_, _40925_);
  and (_41543_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_41544_, _40579_, _41241_);
  or (_41545_, _41544_, _41543_);
  and (_41546_, _41545_, _40778_);
  nor (_41547_, _40579_, _41290_);
  and (_41548_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_41549_, _41548_, _41547_);
  and (_41550_, _41549_, _40939_);
  or (_41551_, _41550_, _41546_);
  or (_41552_, _41551_, _40664_);
  and (_41553_, _41552_, _40963_);
  and (_41554_, _41553_, _41542_);
  nand (_41555_, _40579_, _41315_);
  or (_41556_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_41557_, _41556_, _41555_);
  and (_41558_, _41557_, _40778_);
  or (_41559_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_41560_, _40579_, _41364_);
  and (_41561_, _41560_, _41559_);
  and (_41562_, _41561_, _40939_);
  or (_41563_, _41562_, _41558_);
  or (_41564_, _41563_, _40925_);
  nand (_41565_, _40579_, _41441_);
  or (_41566_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_41567_, _41566_, _41565_);
  and (_41568_, _41567_, _40778_);
  or (_41569_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_41570_, _40579_, _41490_);
  and (_41571_, _41570_, _41569_);
  and (_41572_, _41571_, _40939_);
  or (_41573_, _41572_, _41568_);
  or (_41574_, _41573_, _40664_);
  and (_41575_, _41574_, _40890_);
  and (_41576_, _41575_, _41564_);
  or (_41577_, _41576_, _41554_);
  or (_41578_, _41577_, _40923_);
  or (_41579_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_41580_, _41579_, _41991_);
  and (_01396_, _41580_, _41578_);
  and (_41581_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_41582_, _40579_, _41139_);
  or (_41583_, _41582_, _41581_);
  and (_41584_, _41583_, _40778_);
  nor (_41585_, _40579_, _41194_);
  and (_41586_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_41587_, _41586_, _41585_);
  and (_41588_, _41587_, _40939_);
  or (_41589_, _41588_, _41584_);
  or (_41590_, _41589_, _40925_);
  and (_41591_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_41592_, _40579_, _41244_);
  or (_41593_, _41592_, _41591_);
  and (_41594_, _41593_, _40778_);
  nor (_41595_, _40579_, _41293_);
  and (_41596_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_41597_, _41596_, _41595_);
  and (_41598_, _41597_, _40939_);
  or (_41599_, _41598_, _41594_);
  or (_41600_, _41599_, _40664_);
  and (_41601_, _41600_, _40963_);
  and (_41602_, _41601_, _41590_);
  nand (_41603_, _40579_, _41318_);
  or (_41604_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_41605_, _41604_, _41603_);
  and (_41606_, _41605_, _40778_);
  or (_41607_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand (_41608_, _40579_, _41367_);
  and (_41609_, _41608_, _41607_);
  and (_41610_, _41609_, _40939_);
  or (_41611_, _41610_, _41606_);
  or (_41612_, _41611_, _40925_);
  nand (_41613_, _40579_, _41444_);
  or (_41614_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_41615_, _41614_, _41613_);
  and (_41616_, _41615_, _40778_);
  or (_41617_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand (_41618_, _40579_, _41493_);
  and (_41619_, _41618_, _41617_);
  and (_41620_, _41619_, _40939_);
  or (_41621_, _41620_, _41616_);
  or (_41622_, _41621_, _40664_);
  and (_41623_, _41622_, _40890_);
  and (_41624_, _41623_, _41612_);
  or (_41625_, _41624_, _41602_);
  or (_41626_, _41625_, _40923_);
  or (_41627_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_41628_, _41627_, _41991_);
  and (_01397_, _41628_, _41626_);
  and (_41629_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_41630_, _40579_, _41143_);
  or (_41631_, _41630_, _41629_);
  and (_41632_, _41631_, _40778_);
  nor (_41633_, _40579_, _41197_);
  and (_41634_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_41635_, _41634_, _41633_);
  and (_41636_, _41635_, _40939_);
  or (_41637_, _41636_, _41632_);
  or (_41638_, _41637_, _40925_);
  and (_41639_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_41640_, _40579_, _41247_);
  or (_41641_, _41640_, _41639_);
  and (_41642_, _41641_, _40778_);
  nor (_41643_, _40579_, _41296_);
  and (_41644_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_41645_, _41644_, _41643_);
  and (_41646_, _41645_, _40939_);
  or (_41647_, _41646_, _41642_);
  or (_41648_, _41647_, _40664_);
  and (_41649_, _41648_, _40963_);
  and (_41650_, _41649_, _41638_);
  nand (_41651_, _40579_, _41321_);
  or (_41652_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_41653_, _41652_, _41651_);
  and (_41654_, _41653_, _40778_);
  or (_41655_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_41656_, _40579_, _41370_);
  and (_41657_, _41656_, _41655_);
  and (_41658_, _41657_, _40939_);
  or (_41659_, _41658_, _41654_);
  or (_41660_, _41659_, _40925_);
  nand (_41661_, _40579_, _41447_);
  or (_41662_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_41663_, _41662_, _41661_);
  and (_41664_, _41663_, _40778_);
  or (_41665_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_41666_, _40579_, _41496_);
  and (_41667_, _41666_, _41665_);
  and (_41668_, _41667_, _40939_);
  or (_41669_, _41668_, _41664_);
  or (_41670_, _41669_, _40664_);
  and (_41671_, _41670_, _40890_);
  and (_41672_, _41671_, _41660_);
  or (_41673_, _41672_, _41650_);
  or (_41674_, _41673_, _40923_);
  or (_41675_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_41676_, _41675_, _41991_);
  and (_01399_, _41676_, _41674_);
  and (_41677_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_41678_, _40579_, _41147_);
  or (_41679_, _41678_, _41677_);
  and (_41680_, _41679_, _40778_);
  nor (_41681_, _40579_, _41200_);
  and (_41682_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_41683_, _41682_, _41681_);
  and (_41684_, _41683_, _40939_);
  or (_41685_, _41684_, _41680_);
  or (_41686_, _41685_, _40925_);
  and (_41687_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_41688_, _40579_, _41250_);
  or (_41689_, _41688_, _41687_);
  and (_41690_, _41689_, _40778_);
  nor (_41691_, _40579_, _41299_);
  and (_41692_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_41693_, _41692_, _41691_);
  and (_41694_, _41693_, _40939_);
  or (_41695_, _41694_, _41690_);
  or (_41696_, _41695_, _40664_);
  and (_41697_, _41696_, _40963_);
  and (_41698_, _41697_, _41686_);
  nand (_41699_, _40579_, _41324_);
  or (_41700_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_41701_, _41700_, _41699_);
  and (_41702_, _41701_, _40778_);
  or (_41703_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_41704_, _40579_, _41373_);
  and (_41705_, _41704_, _41703_);
  and (_41706_, _41705_, _40939_);
  or (_41707_, _41706_, _41702_);
  or (_41708_, _41707_, _40925_);
  nand (_41709_, _40579_, _41450_);
  or (_41710_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_41711_, _41710_, _41709_);
  and (_41712_, _41711_, _40778_);
  or (_41713_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_41714_, _40579_, _41499_);
  and (_41715_, _41714_, _41713_);
  and (_41716_, _41715_, _40939_);
  or (_41717_, _41716_, _41712_);
  or (_41718_, _41717_, _40664_);
  and (_41719_, _41718_, _40890_);
  and (_41720_, _41719_, _41708_);
  or (_41721_, _41720_, _41698_);
  or (_41722_, _41721_, _40923_);
  or (_41723_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_41724_, _41723_, _41991_);
  and (_01401_, _41724_, _41722_);
  and (_41725_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_41726_, _40579_, _41151_);
  or (_41727_, _41726_, _41725_);
  and (_41728_, _41727_, _40778_);
  nor (_41729_, _40579_, _41203_);
  and (_41730_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_41731_, _41730_, _41729_);
  and (_41732_, _41731_, _40939_);
  or (_41733_, _41732_, _41728_);
  or (_41734_, _41733_, _40925_);
  and (_41735_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_41736_, _40579_, _41253_);
  or (_41737_, _41736_, _41735_);
  and (_41738_, _41737_, _40778_);
  nor (_41739_, _40579_, _41302_);
  and (_41740_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_41741_, _41740_, _41739_);
  and (_41742_, _41741_, _40939_);
  or (_41743_, _41742_, _41738_);
  or (_41744_, _41743_, _40664_);
  and (_41745_, _41744_, _40963_);
  and (_41746_, _41745_, _41734_);
  nand (_41747_, _40579_, _41327_);
  or (_41748_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_41749_, _41748_, _41747_);
  and (_41750_, _41749_, _40778_);
  or (_41751_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_41752_, _40579_, _41376_);
  and (_41753_, _41752_, _41751_);
  and (_41754_, _41753_, _40939_);
  or (_41755_, _41754_, _41750_);
  or (_41756_, _41755_, _40925_);
  nand (_41757_, _40579_, _41453_);
  or (_41758_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_41759_, _41758_, _41757_);
  and (_41760_, _41759_, _40778_);
  or (_41761_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_41762_, _40579_, _41502_);
  and (_41763_, _41762_, _41761_);
  and (_41764_, _41763_, _40939_);
  or (_41765_, _41764_, _41760_);
  or (_41766_, _41765_, _40664_);
  and (_41767_, _41766_, _40890_);
  and (_41768_, _41767_, _41756_);
  or (_41769_, _41768_, _41746_);
  or (_41770_, _41769_, _40923_);
  or (_41771_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_41772_, _41771_, _41991_);
  and (_01403_, _41772_, _41770_);
  and (_41773_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_41774_, _40579_, _41155_);
  or (_41775_, _41774_, _41773_);
  and (_41776_, _41775_, _40778_);
  nor (_41777_, _40579_, _41206_);
  and (_41778_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_41779_, _41778_, _41777_);
  and (_41780_, _41779_, _40939_);
  or (_41781_, _41780_, _41776_);
  or (_41782_, _41781_, _40925_);
  and (_41783_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_41784_, _40579_, _41256_);
  or (_41785_, _41784_, _41783_);
  and (_41786_, _41785_, _40778_);
  nor (_41787_, _40579_, _41305_);
  and (_41788_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_41789_, _41788_, _41787_);
  and (_41790_, _41789_, _40939_);
  or (_41791_, _41790_, _41786_);
  or (_41792_, _41791_, _40664_);
  and (_41793_, _41792_, _40963_);
  and (_41794_, _41793_, _41782_);
  nand (_41795_, _40579_, _41330_);
  or (_41796_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_41797_, _41796_, _41795_);
  and (_41798_, _41797_, _40778_);
  or (_41799_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_41800_, _40579_, _41379_);
  and (_41801_, _41800_, _41799_);
  and (_41802_, _41801_, _40939_);
  or (_41803_, _41802_, _41798_);
  or (_41804_, _41803_, _40925_);
  nand (_41805_, _40579_, _41456_);
  or (_41806_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_41807_, _41806_, _41805_);
  and (_41808_, _41807_, _40778_);
  or (_41809_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_41810_, _40579_, _41505_);
  and (_41811_, _41810_, _41809_);
  and (_41812_, _41811_, _40939_);
  or (_41813_, _41812_, _41808_);
  or (_41814_, _41813_, _40664_);
  and (_41815_, _41814_, _40890_);
  and (_41816_, _41815_, _41804_);
  or (_41817_, _41816_, _41794_);
  or (_41818_, _41817_, _40923_);
  or (_41819_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_41820_, _41819_, _41991_);
  and (_01405_, _41820_, _41818_);
  and (_41821_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_41822_, _40579_, _41159_);
  or (_41823_, _41822_, _41821_);
  and (_41824_, _41823_, _40778_);
  nor (_41825_, _40579_, _41209_);
  and (_41826_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_41827_, _41826_, _41825_);
  and (_41828_, _41827_, _40939_);
  or (_41829_, _41828_, _41824_);
  or (_41830_, _41829_, _40925_);
  and (_41831_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_41832_, _40579_, _41259_);
  or (_41833_, _41832_, _41831_);
  and (_41834_, _41833_, _40778_);
  nor (_41835_, _40579_, _41308_);
  and (_41836_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_41837_, _41836_, _41835_);
  and (_41838_, _41837_, _40939_);
  or (_41839_, _41838_, _41834_);
  or (_41840_, _41839_, _40664_);
  and (_41841_, _41840_, _40963_);
  and (_41842_, _41841_, _41830_);
  nand (_41843_, _40579_, _41333_);
  or (_41844_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_41845_, _41844_, _41843_);
  and (_41846_, _41845_, _40778_);
  or (_41847_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_41848_, _40579_, _41382_);
  and (_41849_, _41848_, _41847_);
  and (_41850_, _41849_, _40939_);
  or (_41851_, _41850_, _41846_);
  or (_41852_, _41851_, _40925_);
  nand (_41853_, _40579_, _41459_);
  or (_41854_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_41855_, _41854_, _41853_);
  and (_41856_, _41855_, _40778_);
  or (_41857_, _40579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_41858_, _40579_, _41508_);
  and (_41859_, _41858_, _41857_);
  and (_41860_, _41859_, _40939_);
  or (_41861_, _41860_, _41856_);
  or (_41862_, _41861_, _40664_);
  and (_41863_, _41862_, _40890_);
  and (_41864_, _41863_, _41852_);
  or (_41865_, _41864_, _41842_);
  or (_41866_, _41865_, _40923_);
  or (_41867_, _41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_41868_, _41867_, _41991_);
  and (_01407_, _41868_, _41866_);
  or (_41869_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_41870_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_41871_, _41870_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_41872_, _41871_, _41869_);
  nand (_41873_, _41872_, _41991_);
  or (_41874_, \oc8051_gm_cxrom_1.cell0.data [7], _41991_);
  and (_01415_, _41874_, _41873_);
  or (_41875_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41876_, \oc8051_gm_cxrom_1.cell0.data [0], _41870_);
  nand (_41877_, _41876_, _41875_);
  nand (_41878_, _41877_, _41991_);
  or (_41879_, \oc8051_gm_cxrom_1.cell0.data [0], _41991_);
  and (_01422_, _41879_, _41878_);
  or (_41880_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41881_, \oc8051_gm_cxrom_1.cell0.data [1], _41870_);
  nand (_41882_, _41881_, _41880_);
  nand (_41883_, _41882_, _41991_);
  or (_41884_, \oc8051_gm_cxrom_1.cell0.data [1], _41991_);
  and (_01426_, _41884_, _41883_);
  or (_41885_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41886_, \oc8051_gm_cxrom_1.cell0.data [2], _41870_);
  nand (_41887_, _41886_, _41885_);
  nand (_41888_, _41887_, _41991_);
  or (_41889_, \oc8051_gm_cxrom_1.cell0.data [2], _41991_);
  and (_01430_, _41889_, _41888_);
  or (_41890_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41891_, \oc8051_gm_cxrom_1.cell0.data [3], _41870_);
  nand (_41892_, _41891_, _41890_);
  nand (_41893_, _41892_, _41991_);
  or (_41894_, \oc8051_gm_cxrom_1.cell0.data [3], _41991_);
  and (_01434_, _41894_, _41893_);
  or (_41895_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41896_, \oc8051_gm_cxrom_1.cell0.data [4], _41870_);
  nand (_41897_, _41896_, _41895_);
  nand (_41898_, _41897_, _41991_);
  or (_41899_, \oc8051_gm_cxrom_1.cell0.data [4], _41991_);
  and (_01438_, _41899_, _41898_);
  or (_41900_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41901_, \oc8051_gm_cxrom_1.cell0.data [5], _41870_);
  nand (_41902_, _41901_, _41900_);
  nand (_41903_, _41902_, _41991_);
  or (_41904_, \oc8051_gm_cxrom_1.cell0.data [5], _41991_);
  and (_01442_, _41904_, _41903_);
  or (_41905_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_41906_, \oc8051_gm_cxrom_1.cell0.data [6], _41870_);
  nand (_41907_, _41906_, _41905_);
  nand (_41908_, _41907_, _41991_);
  or (_41909_, \oc8051_gm_cxrom_1.cell0.data [6], _41991_);
  and (_01446_, _41909_, _41908_);
  or (_41910_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_41911_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_41912_, _41911_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_41913_, _41912_, _41910_);
  nand (_41914_, _41913_, _41991_);
  or (_41915_, \oc8051_gm_cxrom_1.cell1.data [7], _41991_);
  and (_01467_, _41915_, _41914_);
  or (_41916_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41917_, \oc8051_gm_cxrom_1.cell1.data [0], _41911_);
  nand (_41918_, _41917_, _41916_);
  nand (_41919_, _41918_, _41991_);
  or (_41920_, \oc8051_gm_cxrom_1.cell1.data [0], _41991_);
  and (_01474_, _41920_, _41919_);
  or (_41921_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41922_, \oc8051_gm_cxrom_1.cell1.data [1], _41911_);
  nand (_41923_, _41922_, _41921_);
  nand (_41924_, _41923_, _41991_);
  or (_41925_, \oc8051_gm_cxrom_1.cell1.data [1], _41991_);
  and (_01478_, _41925_, _41924_);
  or (_41926_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41927_, \oc8051_gm_cxrom_1.cell1.data [2], _41911_);
  nand (_41928_, _41927_, _41926_);
  nand (_41929_, _41928_, _41991_);
  or (_41930_, \oc8051_gm_cxrom_1.cell1.data [2], _41991_);
  and (_01482_, _41930_, _41929_);
  or (_41931_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41932_, \oc8051_gm_cxrom_1.cell1.data [3], _41911_);
  nand (_41934_, _41932_, _41931_);
  nand (_41935_, _41934_, _41991_);
  or (_41937_, \oc8051_gm_cxrom_1.cell1.data [3], _41991_);
  and (_01485_, _41937_, _41935_);
  or (_41939_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41941_, \oc8051_gm_cxrom_1.cell1.data [4], _41911_);
  nand (_41943_, _41941_, _41939_);
  nand (_41945_, _41943_, _41991_);
  or (_41947_, \oc8051_gm_cxrom_1.cell1.data [4], _41991_);
  and (_01489_, _41947_, _41945_);
  or (_41948_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41949_, \oc8051_gm_cxrom_1.cell1.data [5], _41911_);
  nand (_41950_, _41949_, _41948_);
  nand (_41951_, _41950_, _41991_);
  or (_41952_, \oc8051_gm_cxrom_1.cell1.data [5], _41991_);
  and (_01493_, _41952_, _41951_);
  or (_41953_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_41954_, \oc8051_gm_cxrom_1.cell1.data [6], _41911_);
  nand (_41955_, _41954_, _41953_);
  nand (_41956_, _41955_, _41991_);
  or (_41957_, \oc8051_gm_cxrom_1.cell1.data [6], _41991_);
  and (_01497_, _41957_, _41956_);
  or (_41958_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_41959_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_41960_, _41959_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_41961_, _41960_, _41958_);
  nand (_41962_, _41961_, _41991_);
  or (_41963_, \oc8051_gm_cxrom_1.cell2.data [7], _41991_);
  and (_01518_, _41963_, _41962_);
  or (_41964_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41965_, \oc8051_gm_cxrom_1.cell2.data [0], _41959_);
  nand (_41966_, _41965_, _41964_);
  nand (_41967_, _41966_, _41991_);
  or (_41968_, \oc8051_gm_cxrom_1.cell2.data [0], _41991_);
  and (_01525_, _41968_, _41967_);
  or (_41969_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41970_, \oc8051_gm_cxrom_1.cell2.data [1], _41959_);
  nand (_41971_, _41970_, _41969_);
  nand (_41972_, _41971_, _41991_);
  or (_41973_, \oc8051_gm_cxrom_1.cell2.data [1], _41991_);
  and (_01529_, _41973_, _41972_);
  or (_41974_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41975_, \oc8051_gm_cxrom_1.cell2.data [2], _41959_);
  nand (_41976_, _41975_, _41974_);
  nand (_41977_, _41976_, _41991_);
  or (_41979_, \oc8051_gm_cxrom_1.cell2.data [2], _41991_);
  and (_01533_, _41979_, _41977_);
  or (_41982_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41984_, \oc8051_gm_cxrom_1.cell2.data [3], _41959_);
  nand (_41986_, _41984_, _41982_);
  nand (_41988_, _41986_, _41991_);
  or (_41990_, \oc8051_gm_cxrom_1.cell2.data [3], _41991_);
  and (_01537_, _41990_, _41988_);
  or (_41992_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41993_, \oc8051_gm_cxrom_1.cell2.data [4], _41959_);
  nand (_41994_, _41993_, _41992_);
  nand (_41995_, _41994_, _41991_);
  or (_41996_, \oc8051_gm_cxrom_1.cell2.data [4], _41991_);
  and (_01541_, _41996_, _41995_);
  or (_41997_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_41998_, \oc8051_gm_cxrom_1.cell2.data [5], _41959_);
  nand (_41999_, _41998_, _41997_);
  nand (_42000_, _41999_, _41991_);
  or (_42001_, \oc8051_gm_cxrom_1.cell2.data [5], _41991_);
  and (_01545_, _42001_, _42000_);
  or (_42002_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_42003_, \oc8051_gm_cxrom_1.cell2.data [6], _41959_);
  nand (_42004_, _42003_, _42002_);
  nand (_42005_, _42004_, _41991_);
  or (_42006_, \oc8051_gm_cxrom_1.cell2.data [6], _41991_);
  and (_01549_, _42006_, _42005_);
  or (_42007_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_42008_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_42009_, _42008_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_42010_, _42009_, _42007_);
  nand (_42011_, _42010_, _41991_);
  or (_42012_, \oc8051_gm_cxrom_1.cell3.data [7], _41991_);
  and (_01570_, _42012_, _42011_);
  or (_42013_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42014_, \oc8051_gm_cxrom_1.cell3.data [0], _42008_);
  nand (_42015_, _42014_, _42013_);
  nand (_42016_, _42015_, _41991_);
  or (_42017_, \oc8051_gm_cxrom_1.cell3.data [0], _41991_);
  and (_01577_, _42017_, _42016_);
  or (_42018_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42019_, \oc8051_gm_cxrom_1.cell3.data [1], _42008_);
  nand (_42020_, _42019_, _42018_);
  nand (_42021_, _42020_, _41991_);
  or (_42022_, \oc8051_gm_cxrom_1.cell3.data [1], _41991_);
  and (_01581_, _42022_, _42021_);
  or (_42023_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42024_, \oc8051_gm_cxrom_1.cell3.data [2], _42008_);
  nand (_42025_, _42024_, _42023_);
  nand (_42026_, _42025_, _41991_);
  or (_42027_, \oc8051_gm_cxrom_1.cell3.data [2], _41991_);
  and (_01585_, _42027_, _42026_);
  or (_42028_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42029_, \oc8051_gm_cxrom_1.cell3.data [3], _42008_);
  nand (_42030_, _42029_, _42028_);
  nand (_42031_, _42030_, _41991_);
  or (_42032_, \oc8051_gm_cxrom_1.cell3.data [3], _41991_);
  and (_01589_, _42032_, _42031_);
  or (_42033_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42034_, \oc8051_gm_cxrom_1.cell3.data [4], _42008_);
  nand (_42035_, _42034_, _42033_);
  nand (_42036_, _42035_, _41991_);
  or (_42037_, \oc8051_gm_cxrom_1.cell3.data [4], _41991_);
  and (_01593_, _42037_, _42036_);
  or (_42038_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42039_, \oc8051_gm_cxrom_1.cell3.data [5], _42008_);
  nand (_42040_, _42039_, _42038_);
  nand (_42041_, _42040_, _41991_);
  or (_42042_, \oc8051_gm_cxrom_1.cell3.data [5], _41991_);
  and (_01596_, _42042_, _42041_);
  or (_42043_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_42044_, \oc8051_gm_cxrom_1.cell3.data [6], _42008_);
  nand (_42045_, _42044_, _42043_);
  nand (_42046_, _42045_, _41991_);
  or (_42047_, \oc8051_gm_cxrom_1.cell3.data [6], _41991_);
  and (_01600_, _42047_, _42046_);
  or (_42048_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_42049_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_42050_, _42049_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_42051_, _42050_, _42048_);
  nand (_42052_, _42051_, _41991_);
  or (_42053_, \oc8051_gm_cxrom_1.cell4.data [7], _41991_);
  and (_01622_, _42053_, _42052_);
  or (_42054_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42055_, \oc8051_gm_cxrom_1.cell4.data [0], _42049_);
  nand (_42056_, _42055_, _42054_);
  nand (_42057_, _42056_, _41991_);
  or (_42058_, \oc8051_gm_cxrom_1.cell4.data [0], _41991_);
  and (_01629_, _42058_, _42057_);
  or (_42059_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42060_, \oc8051_gm_cxrom_1.cell4.data [1], _42049_);
  nand (_42061_, _42060_, _42059_);
  nand (_42062_, _42061_, _41991_);
  or (_42063_, \oc8051_gm_cxrom_1.cell4.data [1], _41991_);
  and (_01632_, _42063_, _42062_);
  or (_42064_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42065_, \oc8051_gm_cxrom_1.cell4.data [2], _42049_);
  nand (_42066_, _42065_, _42064_);
  nand (_42067_, _42066_, _41991_);
  or (_42068_, \oc8051_gm_cxrom_1.cell4.data [2], _41991_);
  and (_01636_, _42068_, _42067_);
  or (_42069_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42070_, \oc8051_gm_cxrom_1.cell4.data [3], _42049_);
  nand (_42071_, _42070_, _42069_);
  nand (_42072_, _42071_, _41991_);
  or (_42073_, \oc8051_gm_cxrom_1.cell4.data [3], _41991_);
  and (_01640_, _42073_, _42072_);
  or (_42074_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42075_, \oc8051_gm_cxrom_1.cell4.data [4], _42049_);
  nand (_42076_, _42075_, _42074_);
  nand (_42077_, _42076_, _41991_);
  or (_42078_, \oc8051_gm_cxrom_1.cell4.data [4], _41991_);
  and (_01644_, _42078_, _42077_);
  or (_42079_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42080_, \oc8051_gm_cxrom_1.cell4.data [5], _42049_);
  nand (_42081_, _42080_, _42079_);
  nand (_42082_, _42081_, _41991_);
  or (_42083_, \oc8051_gm_cxrom_1.cell4.data [5], _41991_);
  and (_01648_, _42083_, _42082_);
  or (_42084_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_42085_, \oc8051_gm_cxrom_1.cell4.data [6], _42049_);
  nand (_42086_, _42085_, _42084_);
  nand (_42087_, _42086_, _41991_);
  or (_42088_, \oc8051_gm_cxrom_1.cell4.data [6], _41991_);
  and (_01652_, _42088_, _42087_);
  or (_42089_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_42090_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_42091_, _42090_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_42092_, _42091_, _42089_);
  nand (_42093_, _42092_, _41991_);
  or (_42094_, \oc8051_gm_cxrom_1.cell5.data [7], _41991_);
  and (_01669_, _42094_, _42093_);
  or (_42095_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42096_, \oc8051_gm_cxrom_1.cell5.data [0], _42090_);
  nand (_42097_, _42096_, _42095_);
  nand (_42098_, _42097_, _41991_);
  or (_42099_, \oc8051_gm_cxrom_1.cell5.data [0], _41991_);
  and (_01671_, _42099_, _42098_);
  or (_42100_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42101_, \oc8051_gm_cxrom_1.cell5.data [1], _42090_);
  nand (_42102_, _42101_, _42100_);
  nand (_42103_, _42102_, _41991_);
  or (_42104_, \oc8051_gm_cxrom_1.cell5.data [1], _41991_);
  and (_01672_, _42104_, _42103_);
  or (_42105_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42106_, \oc8051_gm_cxrom_1.cell5.data [2], _42090_);
  nand (_42107_, _42106_, _42105_);
  nand (_42108_, _42107_, _41991_);
  or (_42109_, \oc8051_gm_cxrom_1.cell5.data [2], _41991_);
  and (_01675_, _42109_, _42108_);
  or (_42110_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42111_, \oc8051_gm_cxrom_1.cell5.data [3], _42090_);
  nand (_42112_, _42111_, _42110_);
  nand (_42113_, _42112_, _41991_);
  or (_42114_, \oc8051_gm_cxrom_1.cell5.data [3], _41991_);
  and (_01679_, _42114_, _42113_);
  or (_42115_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42116_, \oc8051_gm_cxrom_1.cell5.data [4], _42090_);
  nand (_42117_, _42116_, _42115_);
  nand (_42118_, _42117_, _41991_);
  or (_42119_, \oc8051_gm_cxrom_1.cell5.data [4], _41991_);
  and (_01683_, _42119_, _42118_);
  or (_42120_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42121_, \oc8051_gm_cxrom_1.cell5.data [5], _42090_);
  nand (_42122_, _42121_, _42120_);
  nand (_42123_, _42122_, _41991_);
  or (_42124_, \oc8051_gm_cxrom_1.cell5.data [5], _41991_);
  and (_01687_, _42124_, _42123_);
  or (_42125_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_42126_, \oc8051_gm_cxrom_1.cell5.data [6], _42090_);
  nand (_42127_, _42126_, _42125_);
  nand (_42128_, _42127_, _41991_);
  or (_42129_, \oc8051_gm_cxrom_1.cell5.data [6], _41991_);
  and (_01691_, _42129_, _42128_);
  or (_42130_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_42131_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_42132_, _42131_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_42133_, _42132_, _42130_);
  nand (_42134_, _42133_, _41991_);
  or (_42135_, \oc8051_gm_cxrom_1.cell6.data [7], _41991_);
  and (_01713_, _42135_, _42134_);
  or (_42136_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42137_, \oc8051_gm_cxrom_1.cell6.data [0], _42131_);
  nand (_42138_, _42137_, _42136_);
  nand (_42139_, _42138_, _41991_);
  or (_42140_, \oc8051_gm_cxrom_1.cell6.data [0], _41991_);
  and (_01720_, _42140_, _42139_);
  or (_42141_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42142_, \oc8051_gm_cxrom_1.cell6.data [1], _42131_);
  nand (_42143_, _42142_, _42141_);
  nand (_42144_, _42143_, _41991_);
  or (_42145_, \oc8051_gm_cxrom_1.cell6.data [1], _41991_);
  and (_01724_, _42145_, _42144_);
  or (_42146_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42147_, \oc8051_gm_cxrom_1.cell6.data [2], _42131_);
  nand (_42148_, _42147_, _42146_);
  nand (_42149_, _42148_, _41991_);
  or (_42150_, \oc8051_gm_cxrom_1.cell6.data [2], _41991_);
  and (_01728_, _42150_, _42149_);
  or (_42151_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42152_, \oc8051_gm_cxrom_1.cell6.data [3], _42131_);
  nand (_42153_, _42152_, _42151_);
  nand (_42154_, _42153_, _41991_);
  or (_42155_, \oc8051_gm_cxrom_1.cell6.data [3], _41991_);
  and (_01732_, _42155_, _42154_);
  or (_42156_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42157_, \oc8051_gm_cxrom_1.cell6.data [4], _42131_);
  nand (_42158_, _42157_, _42156_);
  nand (_42159_, _42158_, _41991_);
  or (_42160_, \oc8051_gm_cxrom_1.cell6.data [4], _41991_);
  and (_01736_, _42160_, _42159_);
  or (_42161_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42162_, \oc8051_gm_cxrom_1.cell6.data [5], _42131_);
  nand (_42163_, _42162_, _42161_);
  nand (_42164_, _42163_, _41991_);
  or (_42165_, \oc8051_gm_cxrom_1.cell6.data [5], _41991_);
  and (_01740_, _42165_, _42164_);
  or (_42166_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_42167_, \oc8051_gm_cxrom_1.cell6.data [6], _42131_);
  nand (_42168_, _42167_, _42166_);
  nand (_42169_, _42168_, _41991_);
  or (_42170_, \oc8051_gm_cxrom_1.cell6.data [6], _41991_);
  and (_01744_, _42170_, _42169_);
  or (_42171_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_42172_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_42173_, _42172_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_42174_, _42173_, _42171_);
  nand (_42175_, _42174_, _41991_);
  or (_42176_, \oc8051_gm_cxrom_1.cell7.data [7], _41991_);
  and (_01766_, _42176_, _42175_);
  or (_42177_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42178_, \oc8051_gm_cxrom_1.cell7.data [0], _42172_);
  nand (_42179_, _42178_, _42177_);
  nand (_42180_, _42179_, _41991_);
  or (_42181_, \oc8051_gm_cxrom_1.cell7.data [0], _41991_);
  and (_01773_, _42181_, _42180_);
  or (_42182_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42183_, \oc8051_gm_cxrom_1.cell7.data [1], _42172_);
  nand (_42184_, _42183_, _42182_);
  nand (_42185_, _42184_, _41991_);
  or (_42186_, \oc8051_gm_cxrom_1.cell7.data [1], _41991_);
  and (_01777_, _42186_, _42185_);
  or (_42187_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42188_, \oc8051_gm_cxrom_1.cell7.data [2], _42172_);
  nand (_42189_, _42188_, _42187_);
  nand (_42190_, _42189_, _41991_);
  or (_42191_, \oc8051_gm_cxrom_1.cell7.data [2], _41991_);
  and (_01781_, _42191_, _42190_);
  or (_42192_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42193_, \oc8051_gm_cxrom_1.cell7.data [3], _42172_);
  nand (_42194_, _42193_, _42192_);
  nand (_42195_, _42194_, _41991_);
  or (_42196_, \oc8051_gm_cxrom_1.cell7.data [3], _41991_);
  and (_01785_, _42196_, _42195_);
  or (_42197_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42198_, \oc8051_gm_cxrom_1.cell7.data [4], _42172_);
  nand (_42199_, _42198_, _42197_);
  nand (_42200_, _42199_, _41991_);
  or (_42201_, \oc8051_gm_cxrom_1.cell7.data [4], _41991_);
  and (_01788_, _42201_, _42200_);
  or (_42202_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42203_, \oc8051_gm_cxrom_1.cell7.data [5], _42172_);
  nand (_42204_, _42203_, _42202_);
  nand (_42205_, _42204_, _41991_);
  or (_42206_, \oc8051_gm_cxrom_1.cell7.data [5], _41991_);
  and (_01792_, _42206_, _42205_);
  or (_42207_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_42208_, \oc8051_gm_cxrom_1.cell7.data [6], _42172_);
  nand (_42209_, _42208_, _42207_);
  nand (_42210_, _42209_, _41991_);
  or (_42211_, \oc8051_gm_cxrom_1.cell7.data [6], _41991_);
  and (_01796_, _42211_, _42210_);
  or (_42212_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_42213_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_42214_, _42213_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_42215_, _42214_, _42212_);
  nand (_42216_, _42215_, _41991_);
  or (_42217_, \oc8051_gm_cxrom_1.cell8.data [7], _41991_);
  and (_01818_, _42217_, _42216_);
  or (_42218_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42219_, \oc8051_gm_cxrom_1.cell8.data [0], _42213_);
  nand (_42220_, _42219_, _42218_);
  nand (_42221_, _42220_, _41991_);
  or (_42222_, \oc8051_gm_cxrom_1.cell8.data [0], _41991_);
  and (_01824_, _42222_, _42221_);
  or (_42223_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42224_, \oc8051_gm_cxrom_1.cell8.data [1], _42213_);
  nand (_42225_, _42224_, _42223_);
  nand (_42226_, _42225_, _41991_);
  or (_42227_, \oc8051_gm_cxrom_1.cell8.data [1], _41991_);
  and (_01828_, _42227_, _42226_);
  or (_42228_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42229_, \oc8051_gm_cxrom_1.cell8.data [2], _42213_);
  nand (_42230_, _42229_, _42228_);
  nand (_42231_, _42230_, _41991_);
  or (_42232_, \oc8051_gm_cxrom_1.cell8.data [2], _41991_);
  and (_01832_, _42232_, _42231_);
  or (_42233_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42234_, \oc8051_gm_cxrom_1.cell8.data [3], _42213_);
  nand (_42235_, _42234_, _42233_);
  nand (_42236_, _42235_, _41991_);
  or (_42237_, \oc8051_gm_cxrom_1.cell8.data [3], _41991_);
  and (_01836_, _42237_, _42236_);
  or (_42238_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42239_, \oc8051_gm_cxrom_1.cell8.data [4], _42213_);
  nand (_42240_, _42239_, _42238_);
  nand (_42241_, _42240_, _41991_);
  or (_42242_, \oc8051_gm_cxrom_1.cell8.data [4], _41991_);
  and (_01840_, _42242_, _42241_);
  or (_42243_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42244_, \oc8051_gm_cxrom_1.cell8.data [5], _42213_);
  nand (_42245_, _42244_, _42243_);
  nand (_42246_, _42245_, _41991_);
  or (_42247_, \oc8051_gm_cxrom_1.cell8.data [5], _41991_);
  and (_01844_, _42247_, _42246_);
  or (_42248_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_42249_, \oc8051_gm_cxrom_1.cell8.data [6], _42213_);
  nand (_42250_, _42249_, _42248_);
  nand (_42251_, _42250_, _41991_);
  or (_42252_, \oc8051_gm_cxrom_1.cell8.data [6], _41991_);
  and (_01848_, _42252_, _42251_);
  or (_42253_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_42254_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_42255_, _42254_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_42256_, _42255_, _42253_);
  nand (_42257_, _42256_, _41991_);
  or (_42258_, \oc8051_gm_cxrom_1.cell9.data [7], _41991_);
  and (_01869_, _42258_, _42257_);
  or (_42259_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42260_, \oc8051_gm_cxrom_1.cell9.data [0], _42254_);
  nand (_42261_, _42260_, _42259_);
  nand (_42262_, _42261_, _41991_);
  or (_42263_, \oc8051_gm_cxrom_1.cell9.data [0], _41991_);
  and (_01876_, _42263_, _42262_);
  or (_42264_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42265_, \oc8051_gm_cxrom_1.cell9.data [1], _42254_);
  nand (_42266_, _42265_, _42264_);
  nand (_42267_, _42266_, _41991_);
  or (_42268_, \oc8051_gm_cxrom_1.cell9.data [1], _41991_);
  and (_01880_, _42268_, _42267_);
  or (_42269_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42270_, \oc8051_gm_cxrom_1.cell9.data [2], _42254_);
  nand (_42271_, _42270_, _42269_);
  nand (_42272_, _42271_, _41991_);
  or (_42273_, \oc8051_gm_cxrom_1.cell9.data [2], _41991_);
  and (_01884_, _42273_, _42272_);
  or (_42274_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42275_, \oc8051_gm_cxrom_1.cell9.data [3], _42254_);
  nand (_42276_, _42275_, _42274_);
  nand (_42277_, _42276_, _41991_);
  or (_42278_, \oc8051_gm_cxrom_1.cell9.data [3], _41991_);
  and (_01888_, _42278_, _42277_);
  or (_42279_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42280_, \oc8051_gm_cxrom_1.cell9.data [4], _42254_);
  nand (_42281_, _42280_, _42279_);
  nand (_42282_, _42281_, _41991_);
  or (_42283_, \oc8051_gm_cxrom_1.cell9.data [4], _41991_);
  and (_01892_, _42283_, _42282_);
  or (_42284_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42285_, \oc8051_gm_cxrom_1.cell9.data [5], _42254_);
  nand (_42286_, _42285_, _42284_);
  nand (_42287_, _42286_, _41991_);
  or (_42288_, \oc8051_gm_cxrom_1.cell9.data [5], _41991_);
  and (_01895_, _42288_, _42287_);
  or (_42289_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_42290_, \oc8051_gm_cxrom_1.cell9.data [6], _42254_);
  nand (_42291_, _42290_, _42289_);
  nand (_42292_, _42291_, _41991_);
  or (_42293_, \oc8051_gm_cxrom_1.cell9.data [6], _41991_);
  and (_01899_, _42293_, _42292_);
  or (_42294_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_42295_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_42296_, _42295_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_42297_, _42296_, _42294_);
  nand (_42298_, _42297_, _41991_);
  or (_42299_, \oc8051_gm_cxrom_1.cell10.data [7], _41991_);
  and (_01921_, _42299_, _42298_);
  or (_42300_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42301_, \oc8051_gm_cxrom_1.cell10.data [0], _42295_);
  nand (_42302_, _42301_, _42300_);
  nand (_42303_, _42302_, _41991_);
  or (_42304_, \oc8051_gm_cxrom_1.cell10.data [0], _41991_);
  and (_01928_, _42304_, _42303_);
  or (_42305_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42306_, \oc8051_gm_cxrom_1.cell10.data [1], _42295_);
  nand (_42307_, _42306_, _42305_);
  nand (_42308_, _42307_, _41991_);
  or (_42309_, \oc8051_gm_cxrom_1.cell10.data [1], _41991_);
  and (_01932_, _42309_, _42308_);
  or (_42310_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42311_, \oc8051_gm_cxrom_1.cell10.data [2], _42295_);
  nand (_42312_, _42311_, _42310_);
  nand (_42313_, _42312_, _41991_);
  or (_42314_, \oc8051_gm_cxrom_1.cell10.data [2], _41991_);
  and (_01936_, _42314_, _42313_);
  or (_42315_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42316_, \oc8051_gm_cxrom_1.cell10.data [3], _42295_);
  nand (_42317_, _42316_, _42315_);
  nand (_42318_, _42317_, _41991_);
  or (_42319_, \oc8051_gm_cxrom_1.cell10.data [3], _41991_);
  and (_01940_, _42319_, _42318_);
  or (_42320_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42321_, \oc8051_gm_cxrom_1.cell10.data [4], _42295_);
  nand (_42322_, _42321_, _42320_);
  nand (_42323_, _42322_, _41991_);
  or (_42324_, \oc8051_gm_cxrom_1.cell10.data [4], _41991_);
  and (_01944_, _42324_, _42323_);
  or (_42325_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42326_, \oc8051_gm_cxrom_1.cell10.data [5], _42295_);
  nand (_42327_, _42326_, _42325_);
  nand (_42328_, _42327_, _41991_);
  or (_42329_, \oc8051_gm_cxrom_1.cell10.data [5], _41991_);
  and (_01948_, _42329_, _42328_);
  or (_42330_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_42331_, \oc8051_gm_cxrom_1.cell10.data [6], _42295_);
  nand (_42332_, _42331_, _42330_);
  nand (_42333_, _42332_, _41991_);
  or (_42334_, \oc8051_gm_cxrom_1.cell10.data [6], _41991_);
  and (_01951_, _42334_, _42333_);
  or (_42335_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_42336_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_42337_, _42336_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_42338_, _42337_, _42335_);
  nand (_42339_, _42338_, _41991_);
  or (_42340_, \oc8051_gm_cxrom_1.cell11.data [7], _41991_);
  and (_01973_, _42340_, _42339_);
  or (_42341_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42342_, \oc8051_gm_cxrom_1.cell11.data [0], _42336_);
  nand (_42343_, _42342_, _42341_);
  nand (_42344_, _42343_, _41991_);
  or (_42345_, \oc8051_gm_cxrom_1.cell11.data [0], _41991_);
  and (_01980_, _42345_, _42344_);
  or (_42346_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42347_, \oc8051_gm_cxrom_1.cell11.data [1], _42336_);
  nand (_42348_, _42347_, _42346_);
  nand (_42349_, _42348_, _41991_);
  or (_42350_, \oc8051_gm_cxrom_1.cell11.data [1], _41991_);
  and (_01984_, _42350_, _42349_);
  or (_42351_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42352_, \oc8051_gm_cxrom_1.cell11.data [2], _42336_);
  nand (_42353_, _42352_, _42351_);
  nand (_42354_, _42353_, _41991_);
  or (_42355_, \oc8051_gm_cxrom_1.cell11.data [2], _41991_);
  and (_01988_, _42355_, _42354_);
  or (_42356_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42357_, \oc8051_gm_cxrom_1.cell11.data [3], _42336_);
  nand (_42358_, _42357_, _42356_);
  nand (_42359_, _42358_, _41991_);
  or (_42360_, \oc8051_gm_cxrom_1.cell11.data [3], _41991_);
  and (_01992_, _42360_, _42359_);
  or (_42361_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42362_, \oc8051_gm_cxrom_1.cell11.data [4], _42336_);
  nand (_42363_, _42362_, _42361_);
  nand (_42364_, _42363_, _41991_);
  or (_42365_, \oc8051_gm_cxrom_1.cell11.data [4], _41991_);
  and (_01996_, _42365_, _42364_);
  or (_42366_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42367_, \oc8051_gm_cxrom_1.cell11.data [5], _42336_);
  nand (_42368_, _42367_, _42366_);
  nand (_42369_, _42368_, _41991_);
  or (_42370_, \oc8051_gm_cxrom_1.cell11.data [5], _41991_);
  and (_02000_, _42370_, _42369_);
  or (_42371_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_42372_, \oc8051_gm_cxrom_1.cell11.data [6], _42336_);
  nand (_42373_, _42372_, _42371_);
  nand (_42374_, _42373_, _41991_);
  or (_42375_, \oc8051_gm_cxrom_1.cell11.data [6], _41991_);
  and (_02004_, _42375_, _42374_);
  or (_42376_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_42377_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_42378_, _42377_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_42379_, _42378_, _42376_);
  nand (_42380_, _42379_, _41991_);
  or (_42381_, \oc8051_gm_cxrom_1.cell12.data [7], _41991_);
  and (_02025_, _42381_, _42380_);
  or (_42382_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42383_, \oc8051_gm_cxrom_1.cell12.data [0], _42377_);
  nand (_42384_, _42383_, _42382_);
  nand (_42385_, _42384_, _41991_);
  or (_42386_, \oc8051_gm_cxrom_1.cell12.data [0], _41991_);
  and (_02032_, _42386_, _42385_);
  or (_42387_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42388_, \oc8051_gm_cxrom_1.cell12.data [1], _42377_);
  nand (_42389_, _42388_, _42387_);
  nand (_42390_, _42389_, _41991_);
  or (_42391_, \oc8051_gm_cxrom_1.cell12.data [1], _41991_);
  and (_02036_, _42391_, _42390_);
  or (_42392_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42393_, \oc8051_gm_cxrom_1.cell12.data [2], _42377_);
  nand (_42394_, _42393_, _42392_);
  nand (_42395_, _42394_, _41991_);
  or (_42396_, \oc8051_gm_cxrom_1.cell12.data [2], _41991_);
  and (_02040_, _42396_, _42395_);
  or (_42397_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42398_, \oc8051_gm_cxrom_1.cell12.data [3], _42377_);
  nand (_42399_, _42398_, _42397_);
  nand (_42400_, _42399_, _41991_);
  or (_42401_, \oc8051_gm_cxrom_1.cell12.data [3], _41991_);
  and (_02044_, _42401_, _42400_);
  or (_42402_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42403_, \oc8051_gm_cxrom_1.cell12.data [4], _42377_);
  nand (_42404_, _42403_, _42402_);
  nand (_42405_, _42404_, _41991_);
  or (_42406_, \oc8051_gm_cxrom_1.cell12.data [4], _41991_);
  and (_02048_, _42406_, _42405_);
  or (_42407_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42408_, \oc8051_gm_cxrom_1.cell12.data [5], _42377_);
  nand (_42409_, _42408_, _42407_);
  nand (_42410_, _42409_, _41991_);
  or (_42411_, \oc8051_gm_cxrom_1.cell12.data [5], _41991_);
  and (_02052_, _42411_, _42410_);
  or (_42412_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_42413_, \oc8051_gm_cxrom_1.cell12.data [6], _42377_);
  nand (_42414_, _42413_, _42412_);
  nand (_42415_, _42414_, _41991_);
  or (_42416_, \oc8051_gm_cxrom_1.cell12.data [6], _41991_);
  and (_02056_, _42416_, _42415_);
  or (_42417_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_42418_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_42419_, _42418_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_42420_, _42419_, _42417_);
  nand (_42421_, _42420_, _41991_);
  or (_42422_, \oc8051_gm_cxrom_1.cell13.data [7], _41991_);
  and (_02077_, _42422_, _42421_);
  or (_42423_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42424_, \oc8051_gm_cxrom_1.cell13.data [0], _42418_);
  nand (_42425_, _42424_, _42423_);
  nand (_42426_, _42425_, _41991_);
  or (_42427_, \oc8051_gm_cxrom_1.cell13.data [0], _41991_);
  and (_02084_, _42427_, _42426_);
  or (_42428_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42429_, \oc8051_gm_cxrom_1.cell13.data [1], _42418_);
  nand (_42430_, _42429_, _42428_);
  nand (_42431_, _42430_, _41991_);
  or (_42432_, \oc8051_gm_cxrom_1.cell13.data [1], _41991_);
  and (_02088_, _42432_, _42431_);
  or (_42433_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42434_, \oc8051_gm_cxrom_1.cell13.data [2], _42418_);
  nand (_42435_, _42434_, _42433_);
  nand (_42436_, _42435_, _41991_);
  or (_42437_, \oc8051_gm_cxrom_1.cell13.data [2], _41991_);
  and (_02092_, _42437_, _42436_);
  or (_42438_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42439_, \oc8051_gm_cxrom_1.cell13.data [3], _42418_);
  nand (_42440_, _42439_, _42438_);
  nand (_42441_, _42440_, _41991_);
  or (_42442_, \oc8051_gm_cxrom_1.cell13.data [3], _41991_);
  and (_02096_, _42442_, _42441_);
  or (_42443_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42444_, \oc8051_gm_cxrom_1.cell13.data [4], _42418_);
  nand (_42445_, _42444_, _42443_);
  nand (_42446_, _42445_, _41991_);
  or (_42447_, \oc8051_gm_cxrom_1.cell13.data [4], _41991_);
  and (_02100_, _42447_, _42446_);
  or (_42448_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42449_, \oc8051_gm_cxrom_1.cell13.data [5], _42418_);
  nand (_42450_, _42449_, _42448_);
  nand (_42451_, _42450_, _41991_);
  or (_42452_, \oc8051_gm_cxrom_1.cell13.data [5], _41991_);
  and (_02104_, _42452_, _42451_);
  or (_42453_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_42454_, \oc8051_gm_cxrom_1.cell13.data [6], _42418_);
  nand (_42455_, _42454_, _42453_);
  nand (_42456_, _42455_, _41991_);
  or (_42457_, \oc8051_gm_cxrom_1.cell13.data [6], _41991_);
  and (_02108_, _42457_, _42456_);
  or (_42458_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_42459_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_42460_, _42459_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_42461_, _42460_, _42458_);
  nand (_42462_, _42461_, _41991_);
  or (_42463_, \oc8051_gm_cxrom_1.cell14.data [7], _41991_);
  and (_02129_, _42463_, _42462_);
  or (_42464_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42465_, \oc8051_gm_cxrom_1.cell14.data [0], _42459_);
  nand (_42466_, _42465_, _42464_);
  nand (_42467_, _42466_, _41991_);
  or (_42468_, \oc8051_gm_cxrom_1.cell14.data [0], _41991_);
  and (_02136_, _42468_, _42467_);
  or (_42469_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42470_, \oc8051_gm_cxrom_1.cell14.data [1], _42459_);
  nand (_42471_, _42470_, _42469_);
  nand (_42472_, _42471_, _41991_);
  or (_42473_, \oc8051_gm_cxrom_1.cell14.data [1], _41991_);
  and (_02140_, _42473_, _42472_);
  or (_42474_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42475_, \oc8051_gm_cxrom_1.cell14.data [2], _42459_);
  nand (_42476_, _42475_, _42474_);
  nand (_42477_, _42476_, _41991_);
  or (_42478_, \oc8051_gm_cxrom_1.cell14.data [2], _41991_);
  and (_02144_, _42478_, _42477_);
  or (_42479_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42480_, \oc8051_gm_cxrom_1.cell14.data [3], _42459_);
  nand (_42481_, _42480_, _42479_);
  nand (_42482_, _42481_, _41991_);
  or (_42483_, \oc8051_gm_cxrom_1.cell14.data [3], _41991_);
  and (_02148_, _42483_, _42482_);
  or (_42484_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42485_, \oc8051_gm_cxrom_1.cell14.data [4], _42459_);
  nand (_42486_, _42485_, _42484_);
  nand (_42487_, _42486_, _41991_);
  or (_42488_, \oc8051_gm_cxrom_1.cell14.data [4], _41991_);
  and (_02152_, _42488_, _42487_);
  or (_42489_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42490_, \oc8051_gm_cxrom_1.cell14.data [5], _42459_);
  nand (_42491_, _42490_, _42489_);
  nand (_42492_, _42491_, _41991_);
  or (_42493_, \oc8051_gm_cxrom_1.cell14.data [5], _41991_);
  and (_02156_, _42493_, _42492_);
  or (_42494_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_42495_, \oc8051_gm_cxrom_1.cell14.data [6], _42459_);
  nand (_42496_, _42495_, _42494_);
  nand (_42497_, _42496_, _41991_);
  or (_42498_, \oc8051_gm_cxrom_1.cell14.data [6], _41991_);
  and (_02160_, _42498_, _42497_);
  or (_42499_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_42500_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_42501_, _42500_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_42502_, _42501_, _42499_);
  nand (_42503_, _42502_, _41991_);
  or (_42504_, \oc8051_gm_cxrom_1.cell15.data [7], _41991_);
  and (_02181_, _42504_, _42503_);
  or (_42505_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42506_, \oc8051_gm_cxrom_1.cell15.data [0], _42500_);
  nand (_42507_, _42506_, _42505_);
  nand (_42508_, _42507_, _41991_);
  or (_42509_, \oc8051_gm_cxrom_1.cell15.data [0], _41991_);
  and (_02188_, _42509_, _42508_);
  or (_42510_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42511_, \oc8051_gm_cxrom_1.cell15.data [1], _42500_);
  nand (_42512_, _42511_, _42510_);
  nand (_42513_, _42512_, _41991_);
  or (_42514_, \oc8051_gm_cxrom_1.cell15.data [1], _41991_);
  and (_02192_, _42514_, _42513_);
  or (_42515_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42516_, \oc8051_gm_cxrom_1.cell15.data [2], _42500_);
  nand (_42517_, _42516_, _42515_);
  nand (_42518_, _42517_, _41991_);
  or (_42519_, \oc8051_gm_cxrom_1.cell15.data [2], _41991_);
  and (_02196_, _42519_, _42518_);
  or (_42520_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42521_, \oc8051_gm_cxrom_1.cell15.data [3], _42500_);
  nand (_42522_, _42521_, _42520_);
  nand (_42523_, _42522_, _41991_);
  or (_42524_, \oc8051_gm_cxrom_1.cell15.data [3], _41991_);
  and (_02200_, _42524_, _42523_);
  or (_42525_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42526_, \oc8051_gm_cxrom_1.cell15.data [4], _42500_);
  nand (_42527_, _42526_, _42525_);
  nand (_42528_, _42527_, _41991_);
  or (_42529_, \oc8051_gm_cxrom_1.cell15.data [4], _41991_);
  and (_02204_, _42529_, _42528_);
  or (_42530_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42531_, \oc8051_gm_cxrom_1.cell15.data [5], _42500_);
  nand (_42532_, _42531_, _42530_);
  nand (_42533_, _42532_, _41991_);
  or (_42534_, \oc8051_gm_cxrom_1.cell15.data [5], _41991_);
  and (_02208_, _42534_, _42533_);
  or (_42535_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_42536_, \oc8051_gm_cxrom_1.cell15.data [6], _42500_);
  nand (_42537_, _42536_, _42535_);
  nand (_42538_, _42537_, _41991_);
  or (_42539_, \oc8051_gm_cxrom_1.cell15.data [6], _41991_);
  and (_02212_, _42539_, _42538_);
  nor (_05984_, _36430_, rst);
  and (_42540_, _33838_, _41991_);
  nand (_42541_, _42540_, _36496_);
  nor (_42542_, _35530_, _36134_);
  or (_05987_, _42542_, _42541_);
  and (_42543_, _34957_, _34726_);
  and (_42544_, _42543_, _35220_);
  not (_42545_, _36013_);
  nor (_42546_, _34463_, _34222_);
  and (_42547_, _42546_, _42545_);
  and (_42548_, _42547_, _42544_);
  and (_42549_, _34463_, _34222_);
  and (_42550_, _42544_, _35461_);
  and (_42551_, _42550_, _42549_);
  and (_42552_, _42551_, _36013_);
  or (_42553_, _42552_, _42548_);
  and (_42554_, _42553_, _35772_);
  not (_42555_, _34463_);
  and (_42556_, _42555_, _34222_);
  not (_42557_, _35220_);
  and (_42558_, _42543_, _42557_);
  and (_42559_, _42558_, _35461_);
  and (_42560_, _42559_, _35772_);
  and (_42561_, _42560_, _42556_);
  not (_42562_, _34726_);
  and (_42563_, _36013_, _35772_);
  and (_42564_, _42563_, _42546_);
  and (_42565_, _42564_, _42562_);
  not (_42566_, _35461_);
  not (_42567_, _34957_);
  and (_42568_, _42567_, _34726_);
  and (_42569_, _42568_, _42557_);
  and (_42570_, _42569_, _42566_);
  and (_42571_, _42570_, _42564_);
  or (_42572_, _42571_, _42565_);
  and (_42573_, _42545_, _35772_);
  not (_42574_, _34222_);
  and (_42575_, _34463_, _42574_);
  and (_42576_, _42575_, _42573_);
  and (_42577_, _42576_, _42569_);
  and (_42578_, _35220_, _42567_);
  nor (_42579_, _42578_, _42562_);
  not (_42580_, _42579_);
  and (_42581_, _42580_, _42576_);
  or (_42582_, _42581_, _42577_);
  or (_42583_, _42582_, _42572_);
  or (_42584_, _42583_, _42561_);
  nor (_42585_, _36013_, _35772_);
  and (_42586_, _42585_, _42556_);
  nor (_42587_, _42586_, _42566_);
  and (_42588_, _42573_, _42549_);
  not (_42589_, _35772_);
  and (_42590_, _36013_, _42589_);
  and (_42591_, _42556_, _42590_);
  nor (_42592_, _42591_, _42588_);
  nand (_42593_, _42592_, _42587_);
  and (_42594_, _42593_, _42558_);
  not (_42595_, _42563_);
  and (_42596_, _42595_, _42551_);
  or (_42597_, _42596_, _42594_);
  or (_42598_, _42597_, _42584_);
  and (_42599_, _42575_, _42590_);
  and (_42600_, _42599_, _42559_);
  and (_42601_, _42569_, _35461_);
  and (_42602_, _42601_, _42589_);
  and (_42603_, _42602_, _42575_);
  nor (_42604_, _42573_, _42590_);
  and (_42605_, _42604_, _42549_);
  and (_42606_, _42605_, _42559_);
  or (_42607_, _42606_, _42603_);
  or (_42608_, _42607_, _42600_);
  and (_42609_, _42573_, _42556_);
  and (_42610_, _42544_, _42566_);
  and (_42611_, _42610_, _42609_);
  and (_42612_, _42548_, _42589_);
  or (_42613_, _42612_, _42611_);
  and (_42614_, _42575_, _36013_);
  and (_42615_, _42610_, _42614_);
  and (_42616_, _42559_, _42547_);
  or (_42617_, _42616_, _42615_);
  or (_42618_, _42617_, _42613_);
  or (_42619_, _42618_, _42608_);
  or (_42620_, _42619_, _42598_);
  or (_42621_, _42620_, _42554_);
  and (_42622_, _42621_, _33849_);
  not (_42623_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_42624_, _33816_, _15624_);
  and (_42625_, _42624_, _33761_);
  nor (_42626_, _42625_, _42623_);
  or (_42627_, _42626_, rst);
  or (_05990_, _42627_, _42622_);
  nand (_42628_, _34222_, _33827_);
  or (_42629_, _33827_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_42630_, _42629_, _41991_);
  and (_05993_, _42630_, _42628_);
  and (_42631_, \oc8051_top_1.oc8051_sfr1.wait_data , _41991_);
  and (_42632_, _42631_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_42633_, _36145_, _36299_);
  and (_42634_, _36331_, _36507_);
  or (_42635_, _42634_, _42633_);
  and (_42636_, _35530_, _36299_);
  or (_42637_, _42636_, _35552_);
  or (_42638_, _42637_, _37209_);
  and (_42639_, _36145_, _37198_);
  and (_42640_, _37110_, _36134_);
  or (_42641_, _42640_, _42639_);
  nor (_42642_, _42641_, _42638_);
  nand (_42643_, _42642_, _36934_);
  or (_42644_, _42643_, _42635_);
  and (_42645_, _42644_, _42540_);
  or (_05996_, _42645_, _42632_);
  and (_42646_, _35530_, _36200_);
  or (_42647_, _42646_, _36156_);
  and (_42648_, _37099_, _36726_);
  or (_42649_, _42648_, _37712_);
  and (_42650_, _35264_, _36320_);
  and (_42651_, _42650_, _37198_);
  or (_42652_, _42651_, _42649_);
  or (_42653_, _42652_, _42647_);
  and (_42654_, _42653_, _33838_);
  and (_42655_, \oc8051_top_1.oc8051_decoder1.state [0], _15624_);
  and (_42656_, _42655_, _42623_);
  not (_42657_, _36364_);
  and (_42658_, _42657_, _42656_);
  and (_42659_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42660_, _42659_, _42658_);
  or (_42661_, _42660_, _42654_);
  and (_05999_, _42661_, _41991_);
  and (_42662_, _42631_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_42663_, _36331_, _36759_);
  nor (_42664_, _37110_, _36759_);
  nor (_42665_, _42664_, _37245_);
  or (_42666_, _42665_, _42663_);
  and (_42667_, _42650_, _36902_);
  or (_42668_, _42667_, _42666_);
  nor (_42669_, _42664_, _34770_);
  and (_42670_, _36902_, _36715_);
  or (_42671_, _42670_, _42669_);
  or (_42672_, _42671_, _37680_);
  nor (_42673_, _35816_, _34770_);
  and (_42674_, _42673_, _36090_);
  and (_42675_, _36331_, _36584_);
  or (_42676_, _42675_, _42674_);
  or (_42677_, _42676_, _42647_);
  or (_42678_, _42677_, _42672_);
  or (_42679_, _42678_, _42668_);
  and (_42680_, _42679_, _42540_);
  or (_06002_, _42680_, _42662_);
  and (_42681_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42682_, _36649_, _33838_);
  or (_42683_, _42682_, _42681_);
  or (_42684_, _42683_, _42658_);
  and (_06005_, _42684_, _41991_);
  and (_42685_, _36145_, _36189_);
  not (_42686_, _36507_);
  nor (_42687_, _42542_, _42686_);
  nor (_42688_, _42687_, _42685_);
  not (_42689_, _42688_);
  and (_42690_, _42689_, _42656_);
  and (_42691_, _36902_, _36627_);
  and (_42692_, _35012_, _36474_);
  and (_42693_, _42692_, _36167_);
  or (_42694_, _42693_, _42691_);
  or (_42695_, _42694_, _42633_);
  and (_42696_, _42695_, _36408_);
  or (_42697_, _42696_, _42690_);
  and (_42698_, _42694_, _33783_);
  or (_42699_, _42698_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42700_, _42699_, _42697_);
  or (_42701_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _15624_);
  and (_42702_, _42701_, _41991_);
  and (_06008_, _42702_, _42700_);
  and (_42703_, _42631_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_42704_, _37198_, _36902_);
  and (_42705_, _42704_, _36551_);
  and (_42706_, _37110_, _36715_);
  or (_42707_, _42706_, _42670_);
  or (_42708_, _42707_, _42705_);
  and (_42709_, _36627_, _36090_);
  or (_42710_, _42667_, _42640_);
  or (_42711_, _42710_, _42709_);
  or (_42712_, _36156_, _37121_);
  or (_42713_, _42648_, _37306_);
  or (_42714_, _42713_, _42712_);
  or (_42715_, _42714_, _42711_);
  or (_42716_, _42715_, _42708_);
  and (_42717_, _42716_, _42540_);
  or (_06011_, _42717_, _42703_);
  and (_42718_, _42631_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_42719_, _42651_, _37055_);
  and (_42720_, _36145_, _36671_);
  and (_42721_, _42650_, _37275_);
  or (_42722_, _42721_, _42720_);
  or (_42723_, _42722_, _42719_);
  or (_42724_, _42723_, _42671_);
  and (_42725_, _36331_, _37000_);
  or (_42726_, _37088_, _37011_);
  or (_42727_, _42726_, _42725_);
  and (_42728_, _37595_, _37099_);
  and (_42729_, _36978_, _36562_);
  or (_42730_, _42729_, _37821_);
  or (_42731_, _42730_, _42728_);
  or (_42732_, _42731_, _42727_);
  or (_42733_, _42732_, _42724_);
  nor (_42734_, _37648_, _37283_);
  not (_42735_, _42734_);
  not (_42736_, _37176_);
  and (_42737_, _36978_, _36726_);
  and (_42738_, _36233_, _36726_);
  or (_42739_, _42738_, _42737_);
  or (_42740_, _42739_, _42736_);
  or (_42741_, _42740_, _42735_);
  or (_42742_, _42741_, _42668_);
  or (_42743_, _42742_, _42733_);
  and (_42744_, _42743_, _42540_);
  or (_06014_, _42744_, _42718_);
  and (_42745_, _42673_, _36189_);
  and (_42746_, _42650_, _36682_);
  or (_42747_, _42746_, _42745_);
  or (_42748_, _42747_, _37616_);
  and (_42749_, _37595_, _36189_);
  and (_42750_, _36682_, _36715_);
  or (_42751_, _42750_, _42749_);
  or (_42752_, _42751_, _42748_);
  and (_42753_, _36200_, _36485_);
  and (_42754_, _36331_, _36200_);
  or (_42755_, _42754_, _42753_);
  or (_42756_, _42755_, _42752_);
  and (_42757_, _42756_, _33838_);
  nor (_42758_, _36364_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42759_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_42760_, _42759_, _42758_);
  or (_42761_, _42760_, _42757_);
  and (_06017_, _42761_, _41991_);
  or (_42762_, _37339_, _37306_);
  or (_42763_, _42665_, _37292_);
  or (_42764_, _42763_, _42762_);
  and (_42765_, _36222_, _36167_);
  and (_42766_, _42765_, _36485_);
  or (_42767_, _42766_, _37033_);
  or (_42768_, _42767_, _37011_);
  or (_42769_, _42768_, _42691_);
  nand (_42770_, _37220_, _36660_);
  or (_42771_, _42770_, _42769_);
  or (_42772_, _42771_, _42764_);
  or (_42773_, _37691_, _36737_);
  or (_42774_, _42773_, _36847_);
  or (_42775_, _42774_, _42649_);
  and (_42776_, _37595_, _36222_);
  or (_42777_, _42776_, _37648_);
  or (_42778_, _42777_, _36573_);
  and (_42779_, _42673_, _36222_);
  and (_42780_, _36299_, _36715_);
  or (_42781_, _42780_, _42693_);
  or (_42782_, _42781_, _42779_);
  or (_42783_, _42782_, _42778_);
  or (_42784_, _42783_, _42775_);
  or (_42785_, _42784_, _42671_);
  or (_42786_, _42785_, _42772_);
  and (_42787_, _42786_, _33838_);
  or (_42788_, _42698_, _42658_);
  and (_42789_, _33783_, _37471_);
  or (_42790_, _42789_, _42788_);
  and (_42791_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42792_, _42791_, _42790_);
  or (_42793_, _42792_, _42787_);
  and (_06020_, _42793_, _41991_);
  nor (_06079_, _37942_, rst);
  nor (_06081_, _37547_, rst);
  not (_42794_, _42540_);
  or (_06084_, _42688_, _42794_);
  and (_42795_, _35530_, _36496_);
  nor (_42796_, _42795_, _42685_);
  or (_06087_, _42796_, _42794_);
  and (_42797_, _42549_, _42545_);
  and (_42798_, _42797_, _42550_);
  or (_42799_, _42615_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_42800_, _42799_, _42603_);
  or (_42801_, _42800_, _42798_);
  and (_42802_, _42801_, _42625_);
  nor (_42803_, _42624_, _33761_);
  or (_42804_, _42803_, rst);
  or (_06090_, _42804_, _42802_);
  nand (_42805_, _35461_, _33827_);
  or (_42806_, _33827_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_42807_, _42806_, _41991_);
  and (_06093_, _42807_, _42805_);
  not (_42808_, _33827_);
  or (_42809_, _35220_, _42808_);
  or (_42810_, _33827_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_42811_, _42810_, _41991_);
  and (_06096_, _42811_, _42809_);
  nand (_42812_, _34957_, _33827_);
  or (_42813_, _33827_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_42814_, _42813_, _41991_);
  and (_06099_, _42814_, _42812_);
  nand (_42815_, _34726_, _33827_);
  or (_42816_, _33827_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_42817_, _42816_, _41991_);
  and (_06102_, _42817_, _42815_);
  or (_42818_, _35772_, _42808_);
  or (_42819_, _33827_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_42820_, _42819_, _41991_);
  and (_06105_, _42820_, _42818_);
  nand (_42821_, _36013_, _33827_);
  or (_42822_, _33827_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_42823_, _42822_, _41991_);
  and (_06108_, _42823_, _42821_);
  nand (_42824_, _34463_, _33827_);
  or (_42825_, _33827_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_42826_, _42825_, _41991_);
  and (_06111_, _42826_, _42824_);
  and (_42827_, _42739_, _34266_);
  and (_42828_, _36331_, _36244_);
  and (_42829_, _36496_, _36167_);
  and (_42830_, _42829_, _36331_);
  or (_42831_, _42830_, _42828_);
  or (_42832_, _42831_, _37605_);
  and (_42833_, _36726_, _36496_);
  and (_42834_, _42650_, _36836_);
  or (_42835_, _42834_, _42833_);
  or (_42836_, _42835_, _42722_);
  or (_42837_, _42836_, _42832_);
  or (_42838_, _42837_, _42827_);
  and (_42839_, _42650_, _37000_);
  or (_42840_, _42839_, _42646_);
  nor (_42841_, _37252_, _34770_);
  or (_42842_, _42841_, _42840_);
  and (_42843_, _36331_, _36902_);
  and (_42844_, _36331_, _37110_);
  or (_42845_, _42844_, _42843_);
  or (_42846_, _42845_, _42663_);
  or (_42847_, _42846_, _42842_);
  nor (_42848_, _42634_, _36518_);
  nand (_42849_, _42848_, _37832_);
  and (_42850_, _42650_, _36200_);
  or (_42851_, _42850_, _37723_);
  or (_42852_, _42851_, _36156_);
  or (_42853_, _42852_, _42748_);
  or (_42854_, _42853_, _42849_);
  or (_42855_, _42854_, _42847_);
  or (_42856_, _42855_, _42838_);
  and (_42857_, _42856_, _33838_);
  and (_42858_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42859_, _42858_, _42690_);
  or (_42860_, _42859_, _42857_);
  and (_30457_, _42860_, _41991_);
  and (_42861_, _42631_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_42862_, _37275_, _37000_);
  and (_42863_, _42862_, _36627_);
  or (_42864_, _42840_, _42739_);
  or (_42865_, _42864_, _42863_);
  nor (_42866_, _42674_, _37659_);
  not (_42867_, _42866_);
  nor (_42868_, _42867_, _42675_);
  nand (_42869_, _42868_, _37317_);
  or (_42870_, _42869_, _42635_);
  not (_42871_, _37275_);
  nand (_42872_, _42871_, _37252_);
  and (_42873_, _42872_, _36331_);
  or (_42874_, _42873_, _42731_);
  or (_42875_, _42874_, _42870_);
  or (_42876_, _42875_, _42865_);
  and (_42877_, _42876_, _42540_);
  or (_30460_, _42877_, _42861_);
  or (_42878_, _42693_, _37691_);
  or (_42879_, _42878_, _42780_);
  or (_42880_, _42879_, _36847_);
  or (_42881_, _42880_, _42772_);
  and (_42882_, _42881_, _33838_);
  and (_42883_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42884_, _42883_, _42790_);
  or (_42885_, _42884_, _42882_);
  and (_30462_, _42885_, _41991_);
  and (_42886_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42887_, _37268_, _35816_);
  or (_42888_, _42887_, _37712_);
  or (_42889_, _42888_, _42778_);
  or (_42890_, _42889_, _42694_);
  and (_42891_, _42890_, _33838_);
  or (_42892_, _42891_, _42886_);
  or (_42893_, _42892_, _42788_);
  and (_30464_, _42893_, _41991_);
  or (_42894_, _42725_, _42694_);
  or (_42895_, _42841_, _42720_);
  and (_42896_, _42829_, _36485_);
  or (_42897_, _42828_, _42896_);
  and (_42898_, _36331_, _37275_);
  or (_42899_, _42776_, _42898_);
  or (_42900_, _42899_, _42897_);
  or (_42901_, _42900_, _42895_);
  or (_42902_, _42901_, _42894_);
  and (_42903_, _42650_, _36891_);
  or (_42904_, _42903_, _42685_);
  or (_42905_, _42834_, _36353_);
  or (_42906_, _42905_, _42904_);
  and (_42907_, _36331_, _37198_);
  or (_42908_, _42755_, _42907_);
  or (_42910_, _42830_, _36342_);
  and (_42912_, _42650_, _37044_);
  or (_42914_, _42912_, _42634_);
  or (_42916_, _42914_, _42910_);
  or (_42918_, _42916_, _42846_);
  or (_42920_, _42918_, _42908_);
  and (_42922_, _42650_, _37449_);
  and (_42924_, _36836_, _36627_);
  or (_42926_, _42779_, _42924_);
  or (_42928_, _42745_, _37627_);
  or (_42930_, _42749_, _36255_);
  or (_42932_, _42930_, _42928_);
  or (_42934_, _42932_, _42926_);
  or (_42936_, _42934_, _42922_);
  or (_42938_, _42936_, _42920_);
  or (_42940_, _42938_, _42906_);
  or (_42942_, _42940_, _42902_);
  and (_42944_, _42942_, _33838_);
  and (_42946_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42948_, _42690_, _36419_);
  or (_42950_, _42948_, _42946_);
  or (_42952_, _42950_, _42944_);
  and (_30466_, _42952_, _41991_);
  or (_42955_, _42766_, _36847_);
  and (_42957_, _36145_, _37000_);
  and (_42959_, _37275_, _36145_);
  nor (_42961_, _42959_, _42957_);
  nand (_42963_, _42961_, _36266_);
  or (_42965_, _42963_, _42955_);
  and (_42967_, _42776_, _34277_);
  and (_42969_, _42673_, _36496_);
  or (_42970_, _42969_, _42646_);
  or (_42971_, _42970_, _42967_);
  or (_42972_, _36353_, _42749_);
  or (_42973_, _42972_, _42928_);
  or (_42974_, _42973_, _42971_);
  or (_42975_, _42974_, _42965_);
  or (_42976_, _42895_, _37260_);
  or (_42977_, _42976_, _42920_);
  or (_42978_, _42977_, _42975_);
  and (_42979_, _42978_, _33838_);
  and (_42980_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42981_, _42980_, _42948_);
  or (_42982_, _42981_, _42979_);
  and (_30468_, _42982_, _41991_);
  and (_42983_, _42631_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_42984_, _36145_, _36748_);
  and (_42985_, _42984_, _36167_);
  and (_42986_, _42640_, _36112_);
  or (_42987_, _42986_, _42985_);
  not (_42988_, _40490_);
  or (_42989_, _42850_, _42988_);
  or (_42990_, _42989_, _42708_);
  or (_42991_, _42990_, _42987_);
  or (_42992_, _42844_, _42667_);
  or (_42993_, _42762_, _42712_);
  or (_42994_, _42993_, _42992_);
  and (_42995_, _36145_, _37044_);
  or (_42996_, _42995_, _36638_);
  and (_42997_, _36145_, _36891_);
  or (_42998_, _42745_, _42648_);
  or (_42999_, _42998_, _42997_);
  or (_43000_, _42999_, _42996_);
  and (_43001_, _36891_, _36320_);
  and (_43002_, _36891_, _36715_);
  or (_43003_, _43002_, _37723_);
  nor (_43004_, _43003_, _43001_);
  nand (_43005_, _43004_, _40489_);
  or (_43006_, _43005_, _43000_);
  or (_43007_, _43006_, _42994_);
  or (_43008_, _43007_, _42991_);
  and (_43009_, _43008_, _42540_);
  or (_30470_, _43009_, _42983_);
  or (_43010_, _42651_, _37165_);
  and (_43011_, _37110_, _36551_);
  or (_43012_, _43011_, _42729_);
  or (_43013_, _43012_, _43010_);
  or (_43014_, _43013_, _42727_);
  or (_43015_, _43014_, _42906_);
  or (_43016_, _42844_, _42997_);
  and (_43017_, _42746_, _35816_);
  or (_43018_, _43017_, _36255_);
  or (_43019_, _42985_, _43018_);
  or (_43020_, _43019_, _43016_);
  or (_43021_, _42737_, _40465_);
  or (_43022_, _43021_, _36156_);
  or (_43023_, _43022_, _37627_);
  not (_43024_, _36858_);
  or (_43025_, _42841_, _43024_);
  or (_43026_, _43025_, _43023_);
  or (_43027_, _43026_, _43020_);
  or (_43028_, _43027_, _43015_);
  or (_43029_, _36353_, _36408_);
  or (_43030_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15624_);
  and (_43031_, _43030_, _41991_);
  and (_43032_, _43031_, _43029_);
  and (_30472_, _43032_, _43028_);
  or (_43033_, _42830_, _37187_);
  or (_43034_, _43033_, _42995_);
  not (_43035_, _36814_);
  nor (_43036_, _42834_, _36847_);
  and (_43037_, _43036_, _43035_);
  not (_43038_, _37733_);
  or (_43039_, _42651_, _43038_);
  and (_43040_, _36145_, _36682_);
  or (_43041_, _42998_, _43040_);
  nor (_43042_, _43041_, _43039_);
  nand (_43043_, _43042_, _43037_);
  or (_43044_, _43043_, _43034_);
  and (_43045_, _42673_, _36989_);
  or (_43046_, _43045_, _37605_);
  or (_43048_, _42912_, _42850_);
  or (_43049_, _43048_, _42634_);
  or (_43050_, _36353_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_43051_, _42674_, _37154_);
  or (_43052_, _43051_, _43050_);
  or (_43053_, _43052_, _43049_);
  or (_43054_, _43053_, _43046_);
  or (_43055_, _43054_, _42672_);
  or (_43056_, _43055_, _42668_);
  or (_43057_, _43056_, _43044_);
  or (_43058_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15624_);
  and (_43060_, _43058_, _41991_);
  and (_43061_, _43060_, _43029_);
  and (_30474_, _43061_, _43057_);
  or (_43062_, _42992_, _42713_);
  not (_43063_, _43036_);
  or (_43064_, _43046_, _43063_);
  or (_43065_, _43064_, _43062_);
  or (_43066_, _37712_, _37648_);
  nor (_43067_, _43066_, _42984_);
  nand (_43068_, _43067_, _40490_);
  or (_43069_, _43068_, _42671_);
  or (_43070_, _43034_, _42666_);
  or (_43071_, _43070_, _43069_);
  or (_43072_, _43071_, _43065_);
  and (_43073_, _43072_, _33838_);
  and (_43074_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_43075_, _36342_, _15624_);
  or (_43076_, _43075_, _43074_);
  or (_43077_, _43076_, _43073_);
  and (_30476_, _43077_, _41991_);
  and (_43078_, _42631_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_43079_, _35012_);
  and (_43080_, _43079_, _37044_);
  or (_43081_, _43080_, _37328_);
  or (_43082_, _42995_, _42639_);
  or (_43083_, _43082_, _43081_);
  not (_43084_, _40489_);
  or (_43085_, _43016_, _43084_);
  or (_43086_, _43085_, _43083_);
  or (_43087_, _42989_, _42752_);
  or (_43088_, _43087_, _42987_);
  or (_43089_, _43088_, _43086_);
  and (_43090_, _43089_, _42540_);
  or (_30478_, _43090_, _43078_);
  nor (_38991_, _34222_, rst);
  nor (_38992_, _40481_, rst);
  and (_43091_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_43092_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_43093_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_43094_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_43095_, _43094_, _43093_);
  and (_43096_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_43097_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_43098_, _43097_, _43096_);
  and (_43099_, _43098_, _43095_);
  and (_43100_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_43101_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_43102_, _43101_, _43100_);
  and (_43103_, _43102_, _43099_);
  nor (_43104_, _43103_, _33904_);
  nor (_43105_, _43104_, _43092_);
  nor (_43106_, _43105_, _40465_);
  nor (_43107_, _43106_, _43091_);
  nor (_38993_, _43107_, rst);
  nor (_39004_, _35461_, rst);
  and (_39005_, _35220_, _41991_);
  nor (_39006_, _34957_, rst);
  nor (_39007_, _34726_, rst);
  and (_39008_, _35772_, _41991_);
  nor (_39009_, _36013_, rst);
  nor (_39010_, _34463_, rst);
  nor (_39011_, _40556_, rst);
  nor (_39013_, _40727_, rst);
  nor (_39014_, _40641_, rst);
  nor (_39015_, _40518_, rst);
  nor (_39016_, _40686_, rst);
  nor (_39017_, _40621_, rst);
  nor (_39019_, _40828_, rst);
  and (_43108_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_43109_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_43110_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_43111_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_43112_, _43111_, _43110_);
  and (_43113_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_43114_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_43115_, _43114_, _43113_);
  and (_43116_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_43117_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_43118_, _43117_, _43116_);
  and (_43119_, _43118_, _43115_);
  and (_43120_, _43119_, _43112_);
  nor (_43121_, _43120_, _33904_);
  nor (_43122_, _43121_, _43109_);
  nor (_43123_, _43122_, _40465_);
  nor (_43124_, _43123_, _43108_);
  nor (_39020_, _43124_, rst);
  and (_43125_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_43126_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_43127_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_43128_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_43129_, _43128_, _43127_);
  and (_43130_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_43131_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_43132_, _43131_, _43130_);
  and (_43133_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_43134_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_43135_, _43134_, _43133_);
  and (_43136_, _43135_, _43132_);
  and (_43137_, _43136_, _43129_);
  nor (_43138_, _43137_, _33904_);
  nor (_43139_, _43138_, _43126_);
  nor (_43140_, _43139_, _40465_);
  nor (_43141_, _43140_, _43125_);
  nor (_39021_, _43141_, rst);
  and (_43142_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_43143_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_43144_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_43145_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_43146_, _43145_, _43144_);
  and (_43147_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_43148_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_43149_, _43148_, _43147_);
  and (_43150_, _43149_, _43146_);
  and (_43151_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_43152_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_43153_, _43152_, _43151_);
  and (_43154_, _43153_, _43150_);
  nor (_43155_, _43154_, _33904_);
  nor (_43156_, _43155_, _43143_);
  nor (_43157_, _43156_, _40465_);
  nor (_43158_, _43157_, _43142_);
  nor (_39022_, _43158_, rst);
  and (_43159_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_43160_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_43161_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_43162_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_43163_, _43162_, _43161_);
  and (_43164_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_43165_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_43166_, _43165_, _43164_);
  and (_43167_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_43168_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_43169_, _43168_, _43167_);
  and (_43170_, _43169_, _43166_);
  and (_43171_, _43170_, _43163_);
  nor (_43172_, _43171_, _33904_);
  nor (_43173_, _43172_, _43160_);
  nor (_43174_, _43173_, _40465_);
  nor (_43175_, _43174_, _43159_);
  nor (_39023_, _43175_, rst);
  and (_43176_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_43177_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_43178_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_43179_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_43180_, _43179_, _43178_);
  and (_43181_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_43182_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_43183_, _43182_, _43181_);
  and (_43184_, _43183_, _43180_);
  and (_43185_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_43186_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_43187_, _43186_, _43185_);
  and (_43188_, _43187_, _43184_);
  nor (_43189_, _43188_, _33904_);
  nor (_43190_, _43189_, _43177_);
  nor (_43191_, _43190_, _40465_);
  nor (_43192_, _43191_, _43176_);
  nor (_39025_, _43192_, rst);
  and (_43193_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_43194_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_43195_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_43196_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_43197_, _43196_, _43195_);
  and (_43198_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_43199_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_43200_, _43199_, _43198_);
  and (_43201_, _43200_, _43197_);
  and (_43202_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_43203_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_43204_, _43203_, _43202_);
  and (_43205_, _43204_, _43201_);
  nor (_43206_, _43205_, _33904_);
  nor (_43207_, _43206_, _43194_);
  nor (_43208_, _43207_, _40465_);
  nor (_43209_, _43208_, _43193_);
  nor (_39026_, _43209_, rst);
  and (_43210_, _40465_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_43211_, _33904_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_43212_, _34123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_43213_, _33992_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_43214_, _43213_, _43212_);
  and (_43215_, _34035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_43216_, _34145_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_43217_, _43216_, _43215_);
  and (_43218_, _33937_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_43219_, _34079_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_43220_, _43219_, _43218_);
  and (_43221_, _43220_, _43217_);
  and (_43222_, _43221_, _43214_);
  nor (_43223_, _43222_, _33904_);
  nor (_43224_, _43223_, _43211_);
  nor (_43225_, _43224_, _40465_);
  nor (_43226_, _43225_, _43210_);
  nor (_39027_, _43226_, rst);
  and (_43227_, _33849_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_43228_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_43229_, _43227_, _38749_);
  and (_43230_, _43229_, _41991_);
  and (_39052_, _43230_, _43228_);
  not (_43231_, _43227_);
  or (_43232_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _43227_, _41991_);
  and (_43233_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _41991_);
  or (_43234_, _43233_, _00000_);
  and (_39054_, _43234_, _43232_);
  nor (_39091_, _40486_, rst);
  nor (_39092_, _39134_, rst);
  nor (_39093_, _40459_, rst);
  nor (_43235_, _40625_, _39202_);
  and (_43236_, _40625_, _39202_);
  nor (_43237_, _43236_, _43235_);
  nor (_43238_, _40885_, _38997_);
  and (_43239_, _40885_, _38997_);
  nor (_43240_, _43239_, _43238_);
  nand (_43241_, _43240_, _43237_);
  and (_43242_, _40486_, _24960_);
  nor (_43243_, _40486_, _24960_);
  nor (_43244_, _40540_, _25113_);
  and (_43245_, _40540_, _25113_);
  nor (_43246_, _43245_, _43244_);
  nor (_43247_, _40710_, _40779_);
  and (_43248_, _40710_, _40779_);
  nor (_43249_, _43248_, _43247_);
  nand (_43250_, _43249_, _43246_);
  or (_43251_, _43250_, _43243_);
  or (_43252_, _43251_, _43242_);
  nor (_43253_, _43252_, _43241_);
  and (_43254_, _40776_, _30698_);
  nor (_43255_, _40776_, _30698_);
  or (_43256_, _43255_, _43254_);
  nor (_43257_, _40577_, _24433_);
  and (_43258_, _40577_, _24433_);
  nor (_43259_, _43258_, _43257_);
  nor (_43260_, _43259_, _43256_);
  nor (_43261_, _40662_, _24197_);
  and (_43262_, _40662_, _24197_);
  nor (_43263_, _43262_, _43261_);
  nor (_43264_, _43263_, _28076_);
  and (_43265_, _43264_, _43260_);
  and (_43266_, _43265_, _43253_);
  nor (_43267_, _24949_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_43268_, _43267_, _43266_);
  not (_43269_, _43268_);
  nor (_43270_, _36934_, _42655_);
  and (_43271_, _39003_, _28087_);
  and (_43272_, _43271_, _43270_);
  and (_43273_, _43272_, _43253_);
  nor (_43274_, _42636_, _36255_);
  and (_43275_, _30252_, _26028_);
  nand (_43276_, _43275_, _30882_);
  nor (_43277_, _43276_, _31642_);
  and (_43278_, _43277_, _32381_);
  and (_43279_, _43278_, _33126_);
  not (_43280_, _37460_);
  and (_43281_, _40497_, _43280_);
  nor (_43282_, _43281_, _42655_);
  or (_43283_, _43282_, _35553_);
  nor (_43284_, _43283_, _28872_);
  and (_43285_, _43284_, _43279_);
  and (_43286_, _43285_, _26637_);
  and (_43287_, _43270_, _26387_);
  not (_43288_, _35553_);
  nor (_43289_, _43270_, _36057_);
  nor (_43290_, _43289_, _43288_);
  and (_43291_, _43290_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_43292_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_43293_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_43294_, _43293_, _43292_);
  nor (_43295_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_43296_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_43297_, _43296_, _43295_);
  and (_43298_, _43297_, _43294_);
  and (_43299_, _43298_, _37920_);
  or (_43300_, _43299_, _43291_);
  or (_43301_, _43300_, _43287_);
  nor (_43302_, _43301_, _43286_);
  or (_43303_, _36244_, _36891_);
  or (_43304_, _43303_, _36836_);
  and (_43305_, _43304_, _35530_);
  not (_43306_, _43305_);
  not (_43307_, _42706_);
  nor (_43308_, _42912_, _37121_);
  and (_43309_, _43308_, _43307_);
  and (_43310_, _43309_, _42866_);
  and (_43311_, _43310_, _43306_);
  not (_43312_, _43311_);
  and (_43313_, _43312_, _43302_);
  and (_43314_, _35552_, _35816_);
  not (_43316_, _43314_);
  and (_43317_, _43316_, _37482_);
  nor (_43318_, _43317_, _43302_);
  nor (_43319_, _43318_, _43313_);
  and (_43320_, _43319_, _43274_);
  nor (_43322_, _43320_, _37493_);
  and (_43323_, _36748_, _36627_);
  nor (_43324_, _43323_, _42692_);
  nor (_43325_, _43324_, _35564_);
  nor (_43326_, _43325_, _37887_);
  not (_43328_, _43326_);
  nor (_43329_, _43328_, _43322_);
  not (_43330_, _39254_);
  and (_43331_, _43330_, _37920_);
  nor (_43332_, _39002_, _39035_);
  and (_43334_, _43332_, _39045_);
  not (_43335_, _43334_);
  and (_43336_, _43335_, _43290_);
  nor (_43337_, _43336_, _43331_);
  not (_43338_, _43337_);
  nor (_43340_, _43338_, _43329_);
  not (_43341_, _43340_);
  nor (_43342_, _43341_, _43273_);
  and (_43343_, _43342_, _43269_);
  and (_43344_, _43343_, _37438_);
  and (_39097_, _43344_, _41991_);
  and (_39098_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _41991_);
  and (_39099_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _41991_);
  and (_43346_, _37898_, _28022_);
  and (_43347_, _36255_, _33783_);
  not (_43349_, _43347_);
  nor (_43350_, _43349_, _38760_);
  and (_43352_, _42866_, _43281_);
  and (_43353_, _43352_, _43308_);
  nor (_43354_, _43353_, _37493_);
  not (_43355_, _43354_);
  and (_43356_, _43323_, _36408_);
  and (_43357_, _36869_, _36408_);
  nor (_43358_, _43357_, _43356_);
  and (_43360_, _43358_, _37438_);
  and (_43361_, _43360_, _43355_);
  and (_43362_, _43361_, _43325_);
  and (_43364_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_43365_, _43364_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_43366_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43368_, _43366_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_43369_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43370_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_43372_, _43370_, _43369_);
  and (_43373_, _43372_, _43368_);
  and (_43374_, _43373_, _43365_);
  and (_43376_, _43374_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43377_, _43376_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43378_, _43377_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_43380_, _43378_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_43381_, _43380_, _38749_);
  or (_43382_, _43380_, _38749_);
  and (_43384_, _43382_, _43381_);
  and (_43385_, _43384_, _43362_);
  and (_43387_, _43356_, _40482_);
  and (_43388_, _43274_, _43309_);
  nand (_43389_, _43388_, _43352_);
  and (_43390_, _43389_, _33783_);
  or (_43391_, _43357_, _35553_);
  nor (_43392_, _43391_, _43390_);
  nor (_43393_, _43347_, _43325_);
  and (_43395_, _43393_, _43361_);
  and (_43396_, _43395_, _43392_);
  and (_43397_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_43399_, _43397_, _43387_);
  or (_43400_, _43399_, _43385_);
  nor (_43401_, _43400_, _43350_);
  nand (_43403_, _43401_, _43343_);
  or (_43404_, _43403_, _43346_);
  and (_43405_, _43361_, _40482_);
  nor (_43407_, _43361_, _43107_);
  nor (_43408_, _43407_, _43405_);
  not (_43409_, _43408_);
  not (_43411_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_43412_, _43408_, _43411_);
  and (_43413_, _43408_, _43411_);
  nor (_43415_, _43413_, _43412_);
  not (_43416_, _43415_);
  not (_43417_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_43419_, _43361_, _40830_);
  nor (_43420_, _43361_, _43226_);
  nor (_43422_, _43420_, _43419_);
  nor (_43423_, _43422_, _43417_);
  and (_43427_, _43422_, _43417_);
  nor (_43432_, _43427_, _43423_);
  not (_43445_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_43450_, _43361_, _40622_);
  nor (_43451_, _43361_, _43209_);
  nor (_43465_, _43451_, _43450_);
  nor (_43470_, _43465_, _43445_);
  and (_43471_, _43465_, _43445_);
  not (_43483_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_43490_, _43361_, _40687_);
  nor (_43491_, _43361_, _43192_);
  nor (_43501_, _43491_, _43490_);
  or (_43510_, _43501_, _43483_);
  not (_43511_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_43519_, _43361_, _40519_);
  nor (_43528_, _43361_, _43175_);
  nor (_43529_, _43528_, _43519_);
  nor (_43538_, _43529_, _43511_);
  and (_43546_, _43529_, _43511_);
  not (_43547_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_43558_, _43361_, _40642_);
  nor (_43564_, _43361_, _43158_);
  nor (_43565_, _43564_, _43558_);
  nor (_43579_, _43565_, _43547_);
  and (_43580_, _43361_, _40728_);
  nor (_43584_, _43361_, _43141_);
  or (_43591_, _43584_, _43580_);
  and (_43599_, _43591_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_43603_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_43609_, _43361_, _40557_);
  nor (_43621_, _43361_, _43124_);
  nor (_43622_, _43621_, _43609_);
  nor (_43634_, _43622_, _43603_);
  nor (_43641_, _43591_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_43642_, _43641_, _43599_);
  and (_43652_, _43642_, _43634_);
  nor (_43661_, _43652_, _43599_);
  not (_43662_, _43661_);
  and (_43663_, _43565_, _43547_);
  nor (_43665_, _43663_, _43579_);
  and (_43666_, _43665_, _43662_);
  nor (_43667_, _43666_, _43579_);
  nor (_43669_, _43667_, _43546_);
  or (_43670_, _43669_, _43538_);
  nand (_43671_, _43501_, _43483_);
  and (_43673_, _43671_, _43510_);
  nand (_43674_, _43673_, _43670_);
  and (_43675_, _43674_, _43510_);
  nor (_43677_, _43675_, _43471_);
  or (_43678_, _43677_, _43470_);
  and (_43680_, _43678_, _43432_);
  nor (_43681_, _43680_, _43423_);
  nor (_43682_, _43681_, _43416_);
  nor (_43683_, _43682_, _43412_);
  nor (_43685_, _43683_, _38721_);
  and (_43686_, _43685_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_43687_, _43686_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_43689_, _43687_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_43690_, _43689_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_43691_, _43690_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_43693_, _43691_, _43409_);
  and (_43694_, _43683_, _38721_);
  and (_43695_, _43694_, _38727_);
  and (_43697_, _43695_, _38732_);
  and (_43698_, _43697_, _38717_);
  and (_43699_, _43698_, _38738_);
  and (_43701_, _43699_, _38713_);
  nor (_43702_, _43701_, _43408_);
  nor (_43703_, _43702_, _43693_);
  or (_43705_, _43408_, _38744_);
  nand (_43706_, _43408_, _38744_);
  and (_43707_, _43706_, _43705_);
  and (_43709_, _43707_, _43703_);
  or (_43710_, _43709_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_43712_, _43709_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_43713_, _43712_, _43710_);
  not (_43714_, _43361_);
  nor (_43715_, _43393_, _43714_);
  and (_43717_, _35530_, _36408_);
  and (_43718_, _43717_, _36682_);
  and (_43719_, _42673_, _37099_);
  not (_43721_, _43719_);
  and (_43722_, _43308_, _43721_);
  not (_43723_, _35552_);
  and (_43725_, _43274_, _43723_);
  and (_43726_, _43725_, _43722_);
  and (_43727_, _43726_, _43352_);
  nor (_43729_, _43727_, _37493_);
  nor (_43730_, _43729_, _43718_);
  nor (_43731_, _43730_, _43715_);
  and (_43733_, _43731_, _43713_);
  or (_43734_, _43733_, _43404_);
  not (_43735_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_43737_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_43738_, _43737_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_43739_, _43738_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_43741_, _43739_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_43742_, _43741_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_43744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_43745_, _43744_, _43742_);
  and (_43746_, _43745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_43747_, _43746_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_43749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_43750_, _34024_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43751_, _43750_, _40465_);
  nor (_43753_, _43751_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_43754_, _43753_);
  and (_43755_, _43754_, _43749_);
  and (_43757_, _43755_, _43747_);
  nand (_43758_, _43757_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_43759_, _43758_, _43735_);
  or (_43761_, _43758_, _43735_);
  and (_43762_, _43761_, _43759_);
  or (_43763_, _43762_, _43343_);
  and (_43765_, _43763_, _41991_);
  and (_39101_, _43765_, _43734_);
  and (_43766_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _41991_);
  and (_43768_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_43769_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_43770_, _33838_, _43769_);
  not (_43772_, _43770_);
  not (_43773_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_43775_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_43776_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_43777_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_43778_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_43779_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_43780_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_43781_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_43783_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_43784_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43785_, _43784_, _43783_);
  and (_43787_, _43785_, _43781_);
  and (_43788_, _43787_, _43780_);
  and (_43789_, _43788_, _43779_);
  and (_43791_, _43789_, _43778_);
  and (_43792_, _43791_, _43777_);
  and (_43793_, _43792_, _43776_);
  and (_43795_, _43793_, _43775_);
  and (_43796_, _43795_, _43773_);
  nor (_43797_, _43796_, _43735_);
  and (_43799_, _43796_, _43735_);
  nor (_43800_, _43799_, _43797_);
  nor (_43801_, _43795_, _43773_);
  nor (_43803_, _43801_, _43796_);
  not (_43804_, _43803_);
  not (_43805_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_43807_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_43808_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_43810_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_43811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_43812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_43813_, _43812_, _43810_);
  and (_43815_, _43813_, _43811_);
  nor (_43816_, _43815_, _43810_);
  nor (_43817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_43819_, _43817_, _43808_);
  not (_43820_, _43819_);
  nor (_43821_, _43820_, _43816_);
  nor (_43823_, _43821_, _43808_);
  not (_43824_, _43823_);
  and (_43825_, _43824_, _43793_);
  and (_43827_, _43825_, _43807_);
  and (_43828_, _43827_, _43805_);
  and (_43829_, _43828_, _43804_);
  nor (_43831_, _43828_, _43804_);
  or (_43832_, _43831_, _43829_);
  not (_43833_, _43832_);
  and (_43835_, _43823_, _43795_);
  and (_43836_, _43823_, _43793_);
  and (_43837_, _43836_, _43807_);
  nor (_43839_, _43837_, _43805_);
  or (_43840_, _43839_, _43835_);
  nor (_43842_, _43836_, _43807_);
  nor (_43843_, _43842_, _43837_);
  not (_43844_, _43843_);
  and (_43845_, _43823_, _43792_);
  nor (_43847_, _43845_, _43776_);
  nor (_43848_, _43847_, _43836_);
  not (_43849_, _43848_);
  and (_43851_, _43823_, _43789_);
  and (_43852_, _43851_, _43778_);
  nor (_43853_, _43852_, _43777_);
  nor (_43855_, _43853_, _43845_);
  not (_43856_, _43855_);
  nor (_43857_, _43851_, _43778_);
  nor (_43859_, _43857_, _43852_);
  and (_43860_, _43823_, _43787_);
  and (_43861_, _43860_, _43780_);
  nor (_43863_, _43860_, _43780_);
  nor (_43864_, _43863_, _43861_);
  not (_43865_, _43864_);
  and (_43867_, _43823_, _43785_);
  nor (_43868_, _43867_, _43781_);
  nor (_43869_, _43868_, _43860_);
  not (_43871_, _43869_);
  and (_43872_, _43823_, _43784_);
  nor (_43874_, _43872_, _43783_);
  nor (_43875_, _43874_, _43867_);
  not (_43876_, _43875_);
  not (_43877_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_43879_, _43823_, _43877_);
  nor (_43880_, _43823_, _43877_);
  nor (_43881_, _43880_, _43879_);
  not (_43883_, _43881_);
  and (_43884_, _42585_, _42575_);
  nor (_43885_, _43884_, _42609_);
  nor (_43887_, _43885_, _34726_);
  not (_43888_, _43887_);
  and (_43889_, _42578_, _34726_);
  and (_43891_, _42575_, _42589_);
  and (_43892_, _43891_, _43889_);
  nor (_43893_, _43892_, _42565_);
  and (_43895_, _43893_, _43888_);
  not (_43896_, _42570_);
  nor (_43897_, _42599_, _42609_);
  nor (_43899_, _43897_, _43896_);
  not (_43900_, _42559_);
  and (_43901_, _42546_, _36013_);
  nor (_43903_, _43884_, _43901_);
  nor (_43904_, _43903_, _43900_);
  nor (_43906_, _43904_, _43899_);
  and (_43907_, _43906_, _43895_);
  and (_43908_, _42585_, _42546_);
  and (_43909_, _43908_, _42570_);
  and (_43910_, _42588_, _42601_);
  nor (_43912_, _43910_, _43909_);
  and (_43913_, _42601_, _42609_);
  and (_43914_, _42599_, _42562_);
  nor (_43916_, _43914_, _43913_);
  and (_43917_, _43916_, _43912_);
  and (_43918_, _43889_, _42609_);
  nor (_43920_, _43918_, _42581_);
  and (_43921_, _42586_, _42544_);
  and (_43922_, _42570_, _42549_);
  nor (_43924_, _43922_, _43921_);
  and (_43925_, _43924_, _43920_);
  and (_43926_, _43925_, _43917_);
  and (_43928_, _43926_, _43907_);
  not (_43929_, _42550_);
  and (_43930_, _42590_, _42546_);
  not (_43932_, _43930_);
  nor (_43933_, _42591_, _42576_);
  and (_43934_, _43933_, _43932_);
  and (_43936_, _42575_, _42563_);
  or (_43937_, _43936_, _43884_);
  not (_43939_, _43937_);
  nor (_43940_, _42564_, _42609_);
  and (_43941_, _43940_, _43939_);
  and (_43942_, _43941_, _43934_);
  nor (_43944_, _43942_, _43929_);
  and (_43945_, _42576_, _42559_);
  not (_43946_, _43945_);
  and (_43948_, _42610_, _42591_);
  and (_43949_, _42602_, _42797_);
  nor (_43950_, _43949_, _43948_);
  and (_43952_, _43950_, _43946_);
  not (_43953_, _43952_);
  nor (_43954_, _43953_, _43944_);
  and (_43956_, _43954_, _43928_);
  and (_43957_, _43936_, _42559_);
  not (_43958_, _43957_);
  and (_43960_, _42601_, _42576_);
  not (_43961_, _43960_);
  nor (_43962_, _42606_, _42571_);
  and (_43964_, _43962_, _43961_);
  and (_43965_, _43964_, _43958_);
  not (_43966_, _42569_);
  nor (_43968_, _43936_, _42586_);
  and (_43969_, _42591_, _35461_);
  not (_43971_, _43969_);
  and (_43972_, _43971_, _43968_);
  nor (_43973_, _43972_, _43966_);
  and (_43974_, _42573_, _42546_);
  nor (_43976_, _43974_, _42591_);
  and (_43977_, _43976_, _43932_);
  nor (_43978_, _43977_, _43896_);
  nor (_43980_, _43978_, _43973_);
  and (_43981_, _42576_, _42570_);
  and (_43982_, _42556_, _42563_);
  and (_43984_, _42610_, _43982_);
  nor (_43985_, _43984_, _43981_);
  not (_43986_, _43985_);
  not (_43988_, _42599_);
  nor (_43989_, _42559_, _42550_);
  nor (_43990_, _43989_, _43988_);
  nor (_43992_, _43990_, _43986_);
  and (_43993_, _43992_, _43980_);
  nor (_43994_, _42561_, _42552_);
  not (_43996_, _43982_);
  nor (_43997_, _42569_, _42550_);
  nor (_43998_, _43997_, _43996_);
  nor (_44000_, _43998_, _42594_);
  and (_44001_, _44000_, _43994_);
  and (_44003_, _44001_, _43993_);
  and (_44004_, _44003_, _43965_);
  and (_44005_, _44004_, _43956_);
  nor (_44006_, _43813_, _43811_);
  nor (_44008_, _44006_, _43815_);
  not (_44009_, _44008_);
  nor (_44010_, _44009_, _44005_);
  not (_44012_, _44010_);
  and (_44013_, _42610_, _42586_);
  and (_44014_, _42588_, _42559_);
  or (_44016_, _43948_, _44014_);
  nor (_44017_, _44016_, _44013_);
  or (_44018_, _42581_, _42552_);
  or (_44020_, _44018_, _43899_);
  nor (_44021_, _44020_, _43986_);
  and (_44022_, _44021_, _44017_);
  nand (_44024_, _44022_, _43965_);
  nor (_44025_, _44024_, _44005_);
  not (_44026_, _44025_);
  nor (_44028_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_44029_, _44028_, _43811_);
  and (_44030_, _44029_, _44026_);
  and (_44032_, _44009_, _44005_);
  nor (_44033_, _44032_, _44010_);
  nand (_44034_, _44033_, _44030_);
  and (_44035_, _44034_, _44012_);
  not (_44036_, _44035_);
  and (_44037_, _43820_, _43816_);
  nor (_44038_, _44037_, _43821_);
  and (_44039_, _44038_, _44036_);
  and (_44040_, _44039_, _43883_);
  not (_44041_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_44042_, _43879_, _44041_);
  or (_44043_, _44042_, _43872_);
  and (_44044_, _44043_, _44040_);
  and (_44045_, _44044_, _43876_);
  and (_44046_, _44045_, _43871_);
  and (_44047_, _44046_, _43865_);
  nor (_44048_, _43861_, _43779_);
  or (_44049_, _44048_, _43851_);
  nand (_44050_, _44049_, _44047_);
  nor (_44051_, _44050_, _43859_);
  and (_44052_, _44051_, _43856_);
  and (_44053_, _44052_, _43849_);
  and (_44054_, _44053_, _43844_);
  and (_44055_, _44054_, _43840_);
  and (_44056_, _44055_, _43833_);
  nor (_44057_, _44056_, _43829_);
  not (_44058_, _44057_);
  nor (_44059_, _44058_, _43800_);
  and (_44060_, _44058_, _43800_);
  or (_44061_, _44060_, _44059_);
  or (_44062_, _44061_, _43772_);
  or (_44063_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_44064_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_44065_, _44064_, _44063_);
  and (_44066_, _44065_, _44062_);
  or (_39102_, _44066_, _43768_);
  nor (_44067_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_39103_, _44067_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_39104_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _41991_);
  nor (_44068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_44069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_44070_, _44069_, _44068_);
  nor (_44071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_44072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_44073_, _44072_, _44071_);
  and (_44074_, _44073_, _44070_);
  nor (_44075_, _44074_, rst);
  and (_44076_, \oc8051_top_1.oc8051_rom1.ea_int , _33794_);
  nand (_44077_, _44076_, _33838_);
  and (_44078_, _44077_, _39104_);
  or (_39106_, _44078_, _44075_);
  and (_44079_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_44080_, _44079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_39107_, _44080_, _41991_);
  nor (_44081_, _43753_, _40465_);
  nor (_44082_, _44005_, _33970_);
  not (_44083_, _44082_);
  nor (_44084_, _44025_, _34057_);
  and (_44085_, _44005_, _33970_);
  nor (_44086_, _44085_, _44082_);
  nand (_44087_, _44086_, _44084_);
  and (_44088_, _44087_, _44083_);
  nor (_44089_, _44088_, _40465_);
  and (_44090_, _44089_, _33959_);
  nor (_44091_, _44089_, _33959_);
  nor (_44092_, _44091_, _44090_);
  nor (_44093_, _44092_, _44081_);
  and (_44094_, _33981_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_44095_, _44094_, _44081_);
  and (_44096_, _44095_, _44024_);
  or (_44097_, _44096_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_44098_, _44097_, _44093_);
  and (_39108_, _44098_, _41991_);
  not (_44099_, _35154_);
  and (_44100_, _34419_, _44099_);
  not (_44101_, _35706_);
  and (_44102_, _34178_, _44101_);
  and (_44103_, _44102_, _44100_);
  and (_44104_, _33849_, _41991_);
  nand (_44105_, _44104_, _34913_);
  nor (_44106_, _44105_, _34683_);
  not (_44107_, _35970_);
  nor (_44108_, _44107_, _35417_);
  and (_44109_, _44108_, _44106_);
  and (_39111_, _44109_, _44103_);
  nor (_44110_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_44111_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_44112_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_39114_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _41991_);
  and (_44113_, _39114_, _44112_);
  or (_39113_, _44113_, _44111_);
  not (_44114_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_44115_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44116_, _44115_, _44114_);
  and (_44117_, _44115_, _44114_);
  nor (_44118_, _44117_, _44116_);
  not (_44119_, _44118_);
  and (_44120_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_44121_, _44120_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44122_, _44120_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_44123_, _44122_, _44121_);
  or (_44124_, _44123_, _44115_);
  and (_44125_, _44124_, _44119_);
  nor (_44126_, _44116_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_44127_, _44116_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_44128_, _44127_, _44126_);
  or (_44129_, _44121_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_39116_, _44129_, _41991_);
  and (_44130_, _39116_, _44128_);
  and (_39115_, _44130_, _44125_);
  not (_44131_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_44132_, _43753_, _44131_);
  and (_44133_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_44134_, _44132_);
  and (_44135_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_44136_, _44135_, _44133_);
  and (_39117_, _44136_, _41991_);
  and (_44137_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_44138_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_44139_, _44138_, _44137_);
  and (_39118_, _44139_, _41991_);
  and (_44140_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_44141_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_44142_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _44141_);
  and (_44143_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_44144_, _44143_, _44140_);
  and (_39120_, _44144_, _41991_);
  and (_44145_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_44146_, _44145_, _44142_);
  and (_39121_, _44146_, _41991_);
  or (_44147_, _44141_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_39122_, _44147_, _41991_);
  not (_44148_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_44149_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_44150_, _44149_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_44151_, _44141_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_44152_, _44151_, _41991_);
  and (_39123_, _44152_, _44150_);
  or (_44153_, _44141_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_39124_, _44153_, _41991_);
  nor (_44154_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_44155_, _44154_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_44156_, _44155_, _41991_);
  and (_44157_, _39114_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_39125_, _44157_, _44156_);
  and (_44158_, _44131_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_44159_, _44158_, _44155_);
  and (_39126_, _44159_, _41991_);
  nand (_44160_, _44155_, _38760_);
  or (_44161_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_44162_, _44161_, _41991_);
  and (_39127_, _44162_, _44160_);
  nand (_44163_, _36452_, _41991_);
  nor (_39128_, _44163_, _37964_);
  or (_44164_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_44165_, _43227_, _43603_);
  and (_44166_, _44165_, _41991_);
  and (_39164_, _44166_, _44164_);
  or (_44167_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_44168_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_44169_, _43227_, _44168_);
  and (_44170_, _44169_, _41991_);
  and (_39165_, _44170_, _44167_);
  or (_44171_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_44172_, _43227_, _43547_);
  and (_44173_, _44172_, _41991_);
  and (_39166_, _44173_, _44171_);
  or (_44174_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_44175_, _43227_, _43511_);
  and (_44176_, _44175_, _41991_);
  and (_39168_, _44176_, _44174_);
  or (_44177_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_44178_, _43227_, _43483_);
  and (_44179_, _44178_, _41991_);
  and (_39169_, _44179_, _44177_);
  or (_44180_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_44181_, _43227_, _43445_);
  and (_44182_, _44181_, _41991_);
  and (_39170_, _44182_, _44180_);
  or (_44183_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_44184_, _43227_, _43417_);
  and (_44185_, _44184_, _41991_);
  and (_39171_, _44185_, _44183_);
  or (_44186_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_44187_, _43227_, _43411_);
  and (_44188_, _44187_, _41991_);
  and (_39172_, _44188_, _44186_);
  or (_44189_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_44190_, _43227_, _38721_);
  and (_44191_, _44190_, _41991_);
  and (_39173_, _44191_, _44189_);
  or (_44192_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_44193_, _43227_, _38727_);
  and (_44194_, _44193_, _41991_);
  and (_39174_, _44194_, _44192_);
  or (_44195_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_44196_, _43227_, _38732_);
  and (_44197_, _44196_, _41991_);
  and (_39175_, _44197_, _44195_);
  or (_44198_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_44199_, _43227_, _38717_);
  and (_44200_, _44199_, _41991_);
  and (_39176_, _44200_, _44198_);
  or (_44201_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_44202_, _43227_, _38738_);
  and (_44203_, _44202_, _41991_);
  and (_39177_, _44203_, _44201_);
  or (_44204_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_44205_, _43227_, _38713_);
  and (_44206_, _44205_, _41991_);
  and (_39179_, _44206_, _44204_);
  or (_44207_, _43227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_44208_, _43227_, _38744_);
  and (_44209_, _44208_, _41991_);
  and (_39180_, _44209_, _44207_);
  or (_44210_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_44211_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _41991_);
  or (_44212_, _44211_, _00000_);
  and (_39183_, _44212_, _44210_);
  or (_44213_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_44214_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _41991_);
  or (_44215_, _44214_, _00000_);
  and (_39184_, _44215_, _44213_);
  or (_44216_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_44217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _41991_);
  or (_44218_, _44217_, _00000_);
  and (_39185_, _44218_, _44216_);
  or (_44219_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_44220_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _41991_);
  or (_44221_, _44220_, _00000_);
  and (_39186_, _44221_, _44219_);
  or (_44222_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_44223_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _41991_);
  or (_44224_, _44223_, _00000_);
  and (_39187_, _44224_, _44222_);
  or (_44225_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_44226_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _41991_);
  or (_44227_, _44226_, _00000_);
  and (_39188_, _44227_, _44225_);
  or (_44228_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_44229_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _41991_);
  or (_44230_, _44229_, _00000_);
  and (_39189_, _44230_, _44228_);
  or (_44231_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_44232_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _41991_);
  or (_44233_, _44232_, _00000_);
  and (_39190_, _44233_, _44231_);
  or (_44234_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_44235_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _41991_);
  or (_44236_, _44235_, _00000_);
  and (_39192_, _44236_, _44234_);
  or (_44237_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_44238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _41991_);
  or (_44239_, _44238_, _00000_);
  and (_39193_, _44239_, _44237_);
  or (_44240_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_44241_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _41991_);
  or (_44242_, _44241_, _00000_);
  and (_39194_, _44242_, _44240_);
  or (_44243_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_44244_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _41991_);
  or (_44245_, _44244_, _00000_);
  and (_39195_, _44245_, _44243_);
  or (_44246_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_44247_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _41991_);
  or (_44248_, _44247_, _00000_);
  and (_39196_, _44248_, _44246_);
  or (_44249_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_44250_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _41991_);
  or (_44251_, _44250_, _00000_);
  and (_39197_, _44251_, _44249_);
  or (_00008_, _43231_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_00009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _41991_);
  or (_00010_, _00009_, _00000_);
  and (_39198_, _00010_, _00008_);
  and (_00011_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00012_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_00013_, _00012_, _00011_);
  and (_39376_, _00013_, _41991_);
  and (_00014_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00015_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_00016_, _00015_, _00014_);
  and (_39377_, _00016_, _41991_);
  and (_00017_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00018_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00019_, _00018_, _44132_);
  or (_00020_, _00019_, _00017_);
  and (_39378_, _00020_, _41991_);
  and (_00021_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00022_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_00023_, _00022_, _00021_);
  and (_39379_, _00023_, _41991_);
  and (_00024_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00025_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_00026_, _00025_, _00024_);
  and (_39380_, _00026_, _41991_);
  and (_00027_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00028_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00029_, _00028_, _44132_);
  or (_00030_, _00029_, _00027_);
  and (_39381_, _00030_, _41991_);
  and (_00031_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00032_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_00033_, _00032_, _00031_);
  and (_39383_, _00033_, _41991_);
  and (_00034_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00035_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_00036_, _00035_, _00034_);
  and (_39384_, _00036_, _41991_);
  and (_00037_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_00038_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_00039_, _00038_, _00037_);
  and (_39385_, _00039_, _41991_);
  and (_00040_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_00041_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_00042_, _00041_, _00040_);
  and (_39386_, _00042_, _41991_);
  and (_00043_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_00044_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_00045_, _00044_, _00043_);
  and (_39387_, _00045_, _41991_);
  and (_00046_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_00047_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_00048_, _00047_, _00046_);
  and (_39388_, _00048_, _41991_);
  and (_00049_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_00050_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_00051_, _00050_, _00049_);
  and (_39389_, _00051_, _41991_);
  and (_00052_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_00053_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_00054_, _00053_, _00052_);
  and (_39390_, _00054_, _41991_);
  and (_00055_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_00056_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_00057_, _00056_, _00055_);
  and (_39391_, _00057_, _41991_);
  and (_00058_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_00059_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_00060_, _00059_, _00058_);
  and (_39392_, _00060_, _41991_);
  and (_00061_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_00062_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_00063_, _00062_, _00061_);
  and (_39394_, _00063_, _41991_);
  and (_00064_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_00065_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_00066_, _00065_, _00064_);
  and (_39395_, _00066_, _41991_);
  and (_00067_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_00068_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_00069_, _00068_, _00067_);
  and (_39396_, _00069_, _41991_);
  and (_00070_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_00071_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_00072_, _00071_, _00070_);
  and (_39397_, _00072_, _41991_);
  and (_00073_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_00074_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_00075_, _00074_, _00073_);
  and (_39398_, _00075_, _41991_);
  and (_00076_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_00077_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_00078_, _00077_, _00076_);
  and (_39399_, _00078_, _41991_);
  and (_00079_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_00080_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_00081_, _00080_, _00079_);
  and (_39400_, _00081_, _41991_);
  and (_00082_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_00083_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_00084_, _00083_, _00082_);
  and (_39401_, _00084_, _41991_);
  and (_00085_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_00086_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_00087_, _00086_, _00085_);
  and (_39402_, _00087_, _41991_);
  and (_00088_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_00089_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_00090_, _00089_, _00088_);
  and (_39403_, _00090_, _41991_);
  and (_00091_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_00092_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_00093_, _00092_, _00091_);
  and (_39405_, _00093_, _41991_);
  and (_00094_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_00095_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_00096_, _00095_, _00094_);
  and (_39406_, _00096_, _41991_);
  and (_00097_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_00098_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_00099_, _00098_, _00097_);
  and (_39407_, _00099_, _41991_);
  and (_00100_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_00101_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_00102_, _00101_, _00100_);
  and (_39408_, _00102_, _41991_);
  and (_00103_, _44132_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_00104_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_00105_, _00104_, _00103_);
  and (_39409_, _00105_, _41991_);
  nor (_39410_, _35507_, rst);
  nor (_39411_, _35264_, rst);
  nor (_39412_, _35001_, rst);
  nor (_39413_, _40433_, rst);
  nor (_39414_, _40569_, rst);
  nor (_39415_, _40743_, rst);
  nor (_39416_, _40654_, rst);
  nor (_39417_, _40536_, rst);
  nor (_39418_, _40702_, rst);
  nor (_39420_, _40597_, rst);
  nor (_39421_, _40874_, rst);
  and (_39437_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _41991_);
  and (_39438_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _41991_);
  and (_39439_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _41991_);
  and (_39441_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _41991_);
  and (_39442_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _41991_);
  and (_39443_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _41991_);
  and (_39444_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _41991_);
  nor (_00106_, _43396_, _43347_);
  nor (_00107_, _00106_, _29221_);
  not (_00108_, _43356_);
  nor (_00109_, _00108_, _43124_);
  and (_00110_, _43362_, _40557_);
  or (_00111_, _00110_, _00109_);
  and (_00112_, _37427_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00113_, _00112_, _00111_);
  and (_00114_, _43622_, _43603_);
  nor (_00115_, _00114_, _43634_);
  and (_00116_, _00115_, _43731_);
  nor (_00117_, _00116_, _00113_);
  nand (_00118_, _00117_, _43343_);
  or (_00119_, _00118_, _00107_);
  or (_00120_, _43343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00121_, _00120_, _41991_);
  and (_39445_, _00121_, _00119_);
  not (_00122_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_00123_, _43344_, _00122_);
  and (_00124_, _43591_, _43325_);
  or (_00125_, _43642_, _43634_);
  not (_00126_, _43731_);
  nor (_00127_, _00126_, _43652_);
  and (_00128_, _00127_, _00125_);
  or (_00129_, _00128_, _00124_);
  nor (_00130_, _00106_, _29894_);
  or (_00131_, _00130_, _00129_);
  and (_00132_, _00131_, _43343_);
  or (_00133_, _00132_, _00123_);
  and (_39446_, _00133_, _41991_);
  nor (_00134_, _00106_, _30578_);
  nor (_00135_, _00108_, _43158_);
  and (_00136_, _43362_, _40642_);
  or (_00137_, _00136_, _00135_);
  and (_00138_, _37427_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_00139_, _00138_, _00137_);
  or (_00140_, _00139_, _00134_);
  nor (_00141_, _43665_, _43662_);
  nor (_00142_, _00141_, _43666_);
  nand (_00143_, _00142_, _43731_);
  nand (_00144_, _00143_, _43343_);
  or (_00145_, _00144_, _00140_);
  not (_00146_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00147_, _43753_, _00146_);
  and (_00148_, _43753_, _00146_);
  nor (_00149_, _00148_, _00147_);
  or (_00150_, _00149_, _43343_);
  and (_00151_, _00150_, _41991_);
  and (_39447_, _00151_, _00145_);
  nor (_00152_, _00106_, _31327_);
  or (_00153_, _43546_, _43538_);
  or (_00154_, _00153_, _43667_);
  nor (_00155_, _43392_, _43715_);
  nand (_00156_, _00153_, _43667_);
  and (_00157_, _00156_, _00155_);
  nand (_00158_, _00157_, _00154_);
  nor (_00159_, _00108_, _43175_);
  and (_00160_, _37898_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_00161_, _43519_, _43325_);
  or (_00162_, _00161_, _00160_);
  nor (_00163_, _00162_, _00159_);
  and (_00164_, _00163_, _00158_);
  nand (_00165_, _00164_, _43343_);
  or (_00166_, _00165_, _00152_);
  and (_00167_, _00147_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00168_, _00147_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00169_, _00168_, _00167_);
  or (_00170_, _00169_, _43343_);
  and (_00171_, _00170_, _41991_);
  and (_39448_, _00171_, _00166_);
  nor (_00172_, _00106_, _32022_);
  nor (_00173_, _00108_, _43192_);
  and (_00174_, _43362_, _40687_);
  or (_00175_, _00174_, _00173_);
  and (_00176_, _37427_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00177_, _00176_, _00175_);
  or (_00178_, _43673_, _43670_);
  and (_00179_, _43731_, _43674_);
  and (_00180_, _00179_, _00178_);
  nor (_00181_, _00180_, _00177_);
  nand (_00182_, _00181_, _43343_);
  or (_00183_, _00182_, _00172_);
  and (_00184_, _43738_, _43754_);
  nor (_00185_, _00167_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00186_, _00185_, _00184_);
  or (_00187_, _00186_, _43343_);
  and (_00188_, _00187_, _41991_);
  and (_39449_, _00188_, _00183_);
  nor (_00189_, _00106_, _32842_);
  nor (_00190_, _00108_, _43209_);
  and (_00191_, _43362_, _40622_);
  or (_00192_, _00191_, _00190_);
  and (_00193_, _37427_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00194_, _00193_, _00192_);
  or (_00195_, _43470_, _43471_);
  nand (_00196_, _00195_, _43675_);
  or (_00197_, _00195_, _43675_);
  and (_00198_, _00197_, _00155_);
  and (_00199_, _00198_, _00196_);
  nor (_00200_, _00199_, _00194_);
  nand (_00201_, _00200_, _43343_);
  or (_00202_, _00201_, _00189_);
  and (_00203_, _43739_, _43754_);
  nor (_00204_, _00184_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00205_, _00204_, _00203_);
  or (_00206_, _00205_, _43343_);
  and (_00207_, _00206_, _41991_);
  and (_39450_, _00207_, _00202_);
  nor (_00208_, _00106_, _33554_);
  nor (_00209_, _00108_, _43226_);
  and (_00210_, _43362_, _40830_);
  or (_00211_, _00210_, _00209_);
  or (_00212_, _43678_, _43432_);
  nor (_00213_, _00126_, _43680_);
  and (_00214_, _00213_, _00212_);
  or (_00215_, _00214_, _00211_);
  and (_00216_, _37427_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00217_, _00216_, _00215_);
  nand (_00218_, _00217_, _43343_);
  or (_00219_, _00218_, _00208_);
  and (_00220_, _00203_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00221_, _00203_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00222_, _00221_, _00220_);
  or (_00223_, _00222_, _43343_);
  and (_00224_, _00223_, _41991_);
  and (_39452_, _00224_, _00219_);
  nand (_00225_, _37427_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_00226_, _00106_, _28011_);
  or (_00227_, _00108_, _43107_);
  nand (_00228_, _43362_, _40482_);
  and (_00229_, _00228_, _00227_);
  and (_00230_, _43681_, _43416_);
  or (_00231_, _00126_, _43682_);
  or (_00232_, _00231_, _00230_);
  and (_00233_, _00232_, _00229_);
  and (_00234_, _00233_, _00226_);
  and (_00235_, _00234_, _00225_);
  nand (_00236_, _00235_, _43343_);
  and (_00237_, _00220_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00238_, _00220_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00239_, _00238_, _00237_);
  or (_00240_, _00239_, _43343_);
  and (_00241_, _00240_, _41991_);
  and (_39453_, _00241_, _00236_);
  and (_00242_, _37898_, _29232_);
  nor (_00243_, _43349_, _38795_);
  nor (_00244_, _43683_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00245_, _43683_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00246_, _00245_, _00244_);
  or (_00247_, _00246_, _43408_);
  nand (_00248_, _00246_, _43408_);
  and (_00249_, _00248_, _00155_);
  and (_00250_, _00249_, _00247_);
  and (_00251_, _43356_, _40557_);
  and (_00252_, _43362_, _42545_);
  and (_00253_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00254_, _00253_, _00252_);
  nor (_00255_, _00254_, _00251_);
  nand (_00256_, _00255_, _43343_);
  or (_00257_, _00256_, _00250_);
  or (_00258_, _00257_, _00243_);
  or (_00259_, _00258_, _00242_);
  and (_00260_, _00237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00261_, _00237_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00262_, _00261_, _00260_);
  or (_00263_, _00262_, _43343_);
  and (_00264_, _00263_, _41991_);
  and (_39454_, _00264_, _00259_);
  nor (_00265_, _43349_, _38823_);
  and (_00266_, _43362_, _42555_);
  and (_00267_, _43356_, _40728_);
  and (_00268_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_00269_, _00268_, _00267_);
  or (_00270_, _00269_, _00266_);
  or (_00271_, _00270_, _00265_);
  nor (_00272_, _37438_, _29894_);
  or (_00273_, _00272_, _00271_);
  nor (_00274_, _43694_, _43408_);
  nor (_00275_, _43685_, _43409_);
  nor (_00276_, _00275_, _00274_);
  nor (_00277_, _00276_, _38727_);
  and (_00278_, _00276_, _38727_);
  or (_00279_, _00278_, _00277_);
  nand (_00280_, _00279_, _43731_);
  nand (_00281_, _00280_, _43343_);
  or (_00282_, _00281_, _00273_);
  and (_00283_, _43745_, _43754_);
  nor (_00284_, _00260_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00285_, _00284_, _00283_);
  or (_00286_, _00285_, _43343_);
  and (_00287_, _00286_, _41991_);
  and (_39455_, _00287_, _00282_);
  or (_00288_, _37438_, _30578_);
  or (_00289_, _43349_, _38851_);
  nand (_00290_, _43356_, _40642_);
  nand (_00291_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00292_, _00291_, _00290_);
  and (_00293_, _00292_, _00289_);
  nand (_00294_, _43362_, _42574_);
  and (_00295_, _43686_, _43408_);
  and (_00296_, _43695_, _43409_);
  or (_00297_, _00296_, _00295_);
  and (_00298_, _00297_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_00299_, _00297_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_00300_, _00299_, _00126_);
  or (_00301_, _00300_, _00298_);
  and (_00302_, _00301_, _00294_);
  and (_00303_, _00302_, _00293_);
  and (_00304_, _00303_, _00288_);
  nand (_00305_, _00304_, _43343_);
  and (_00306_, _00283_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00307_, _00283_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00308_, _00307_, _00306_);
  or (_00309_, _00308_, _43343_);
  and (_00310_, _00309_, _41991_);
  and (_39456_, _00310_, _00305_);
  and (_00311_, _37898_, _31338_);
  and (_00312_, _43687_, _43408_);
  and (_00313_, _43697_, _43409_);
  nor (_00314_, _00313_, _00312_);
  and (_00315_, _00314_, _38717_);
  or (_00316_, _00314_, _38717_);
  nand (_00317_, _00316_, _00155_);
  nor (_00318_, _00317_, _00315_);
  or (_00319_, _43349_, _38880_);
  nand (_00320_, _43356_, _40519_);
  nor (_00321_, _43374_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00322_, _00321_, _43376_);
  nand (_00323_, _00322_, _43362_);
  nand (_00324_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_00325_, _00324_, _00323_);
  and (_00326_, _00325_, _00320_);
  and (_00327_, _00326_, _00319_);
  nand (_00328_, _00327_, _43343_);
  or (_00329_, _00328_, _00318_);
  or (_00330_, _00329_, _00311_);
  and (_00331_, _00306_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00332_, _00306_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00333_, _00332_, _00331_);
  or (_00334_, _00333_, _43343_);
  and (_00335_, _00334_, _41991_);
  and (_39457_, _00335_, _00330_);
  and (_00336_, _43689_, _43408_);
  and (_00337_, _43698_, _43409_);
  nor (_00338_, _00337_, _00336_);
  and (_00339_, _00338_, _38738_);
  or (_00340_, _00338_, _38738_);
  nand (_00341_, _00340_, _00155_);
  nor (_00342_, _00341_, _00339_);
  and (_00343_, _37898_, _32033_);
  or (_00344_, _43349_, _38910_);
  nand (_00345_, _43356_, _40687_);
  nor (_00346_, _43376_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00347_, _00346_, _43377_);
  nand (_00348_, _00347_, _43362_);
  nand (_00349_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_00350_, _00349_, _00348_);
  and (_00351_, _00350_, _00345_);
  and (_00352_, _00351_, _00344_);
  nand (_00353_, _00352_, _43343_);
  or (_00354_, _00353_, _00343_);
  or (_00355_, _00354_, _00342_);
  and (_00356_, _00331_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00357_, _00331_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00358_, _00357_, _00356_);
  or (_00359_, _00358_, _43343_);
  and (_00360_, _00359_, _41991_);
  and (_39458_, _00360_, _00355_);
  and (_00361_, _43690_, _43408_);
  and (_00362_, _43699_, _43409_);
  nor (_00363_, _00362_, _00361_);
  nand (_00364_, _00363_, _38713_);
  or (_00365_, _00363_, _38713_);
  and (_00366_, _00365_, _00155_);
  and (_00367_, _00366_, _00364_);
  and (_00368_, _37898_, _32853_);
  nor (_00369_, _43349_, _38940_);
  nor (_00370_, _43377_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00371_, _00370_, _43378_);
  and (_00372_, _00371_, _43362_);
  and (_00373_, _43356_, _40622_);
  and (_00374_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00375_, _00374_, _00373_);
  or (_00376_, _00375_, _00372_);
  nor (_00377_, _00376_, _00369_);
  nand (_00378_, _00377_, _43343_);
  or (_00379_, _00378_, _00368_);
  or (_00380_, _00379_, _00367_);
  or (_00381_, _00356_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_00382_, _00356_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_00383_, _00382_, _00381_);
  or (_00384_, _00383_, _43343_);
  and (_00385_, _00384_, _41991_);
  and (_39459_, _00385_, _00380_);
  and (_00386_, _43703_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_00387_, _43703_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_00388_, _00387_, _00155_);
  nor (_00389_, _00388_, _00386_);
  and (_00390_, _37898_, _33565_);
  or (_00391_, _43349_, _38967_);
  or (_00392_, _43378_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00393_, _00392_, _43380_);
  nand (_00394_, _00393_, _43362_);
  nand (_00395_, _43356_, _40830_);
  nand (_00396_, _43396_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00397_, _00396_, _00395_);
  and (_00398_, _00397_, _00394_);
  and (_00399_, _00398_, _00391_);
  nand (_00400_, _00399_, _43343_);
  or (_00401_, _00400_, _00390_);
  or (_00402_, _00401_, _00389_);
  or (_00403_, _43757_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00404_, _00403_, _43758_);
  or (_00405_, _00404_, _43343_);
  and (_00406_, _00405_, _41991_);
  and (_39460_, _00406_, _00402_);
  and (_00407_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_00408_, _44029_, _44026_);
  nor (_00409_, _00408_, _44030_);
  or (_00410_, _00409_, _43772_);
  or (_00411_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00412_, _00411_, _44064_);
  and (_00413_, _00412_, _00410_);
  or (_39461_, _00413_, _00407_);
  or (_00414_, _44033_, _44030_);
  and (_00415_, _00414_, _44034_);
  or (_00416_, _00415_, _43772_);
  or (_00417_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00418_, _00417_, _44064_);
  and (_00419_, _00418_, _00416_);
  and (_00420_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_39463_, _00420_, _00419_);
  and (_00421_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00422_, _44038_, _44036_);
  nor (_00423_, _00422_, _44039_);
  or (_00424_, _00423_, _43772_);
  or (_00425_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00426_, _00425_, _44064_);
  and (_00427_, _00426_, _00424_);
  or (_39464_, _00427_, _00421_);
  and (_00428_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00429_, _44039_, _43883_);
  nor (_00430_, _00429_, _44040_);
  or (_00431_, _00430_, _43772_);
  or (_00432_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00433_, _00432_, _44064_);
  and (_00434_, _00433_, _00431_);
  or (_39465_, _00434_, _00428_);
  nor (_00435_, _44043_, _44040_);
  nor (_00436_, _00435_, _44044_);
  or (_00437_, _00436_, _43772_);
  or (_00438_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00439_, _00438_, _44064_);
  and (_00440_, _00439_, _00437_);
  and (_00441_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_39466_, _00441_, _00440_);
  and (_00442_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00443_, _44044_, _43876_);
  nor (_00444_, _00443_, _44045_);
  or (_00445_, _00444_, _43772_);
  or (_00446_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00447_, _00446_, _44064_);
  and (_00448_, _00447_, _00445_);
  or (_39467_, _00448_, _00442_);
  nor (_00449_, _44045_, _43871_);
  nor (_00450_, _00449_, _44046_);
  or (_00451_, _00450_, _43772_);
  or (_00452_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00453_, _00452_, _44064_);
  and (_00454_, _00453_, _00451_);
  and (_00455_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_39468_, _00455_, _00454_);
  and (_00456_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00457_, _44046_, _43865_);
  nor (_00458_, _00457_, _44047_);
  or (_00459_, _00458_, _43772_);
  or (_00460_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00461_, _00460_, _44064_);
  and (_00462_, _00461_, _00459_);
  or (_39469_, _00462_, _00456_);
  or (_00463_, _44049_, _44047_);
  and (_00464_, _00463_, _44050_);
  or (_00465_, _00464_, _43772_);
  or (_00466_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00467_, _00466_, _44064_);
  and (_00468_, _00467_, _00465_);
  and (_00469_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_39470_, _00469_, _00468_);
  and (_00470_, _44050_, _43859_);
  nor (_00471_, _00470_, _44051_);
  or (_00472_, _00471_, _43772_);
  or (_00473_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00474_, _00473_, _44064_);
  and (_00475_, _00474_, _00472_);
  and (_00476_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_39471_, _00476_, _00475_);
  nor (_00477_, _44051_, _43856_);
  nor (_00478_, _00477_, _44052_);
  or (_00479_, _00478_, _43772_);
  or (_00480_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00481_, _00480_, _44064_);
  and (_00482_, _00481_, _00479_);
  and (_00483_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_39472_, _00483_, _00482_);
  nor (_00484_, _44052_, _43849_);
  nor (_00485_, _00484_, _44053_);
  or (_00486_, _00485_, _43772_);
  or (_00487_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00488_, _00487_, _44064_);
  and (_00489_, _00488_, _00486_);
  and (_00490_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_39474_, _00490_, _00489_);
  nor (_00491_, _44053_, _43844_);
  nor (_00492_, _00491_, _44054_);
  or (_00493_, _00492_, _43772_);
  or (_00494_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00495_, _00494_, _44064_);
  and (_00496_, _00495_, _00493_);
  and (_00497_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_39475_, _00497_, _00496_);
  and (_00498_, _43766_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_00499_, _44054_, _43840_);
  nor (_00500_, _00499_, _44055_);
  or (_00501_, _00500_, _43772_);
  or (_00502_, _43770_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00503_, _00502_, _44064_);
  and (_00504_, _00503_, _00501_);
  or (_39476_, _00504_, _00498_);
  or (_00505_, _44055_, _43833_);
  nor (_00506_, _43772_, _44056_);
  and (_00507_, _00506_, _00505_);
  nor (_00508_, _43770_, _38744_);
  or (_00509_, _00508_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00510_, _00509_, _00507_);
  or (_00511_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _33794_);
  and (_00512_, _00511_, _41991_);
  and (_39477_, _00512_, _00510_);
  and (_00513_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_00514_, _00513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_39478_, _00514_, _41991_);
  and (_00515_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_00516_, _00515_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_39479_, _00516_, _41991_);
  and (_00517_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_00518_, _00517_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_39480_, _00518_, _41991_);
  and (_00519_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_00520_, _00519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_39481_, _00520_, _41991_);
  and (_00521_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_00522_, _00521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_39482_, _00522_, _41991_);
  and (_00523_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_00524_, _00523_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_39483_, _00524_, _41991_);
  and (_00525_, _44074_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_00526_, _00525_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_39485_, _00526_, _41991_);
  nor (_00527_, _44025_, _40465_);
  nand (_00528_, _00527_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00529_, _00527_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00530_, _00529_, _44064_);
  and (_39486_, _00530_, _00528_);
  or (_00531_, _44086_, _44084_);
  and (_00532_, _00531_, _44087_);
  or (_00533_, _00532_, _40465_);
  or (_00534_, _33838_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00535_, _00534_, _44064_);
  and (_39487_, _00535_, _00533_);
  and (_00536_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00537_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_00538_, _00537_, _39114_);
  or (_39503_, _00538_, _00536_);
  and (_00539_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00540_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00541_, _00540_, _39114_);
  or (_39504_, _00541_, _00539_);
  and (_00542_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00543_, _00018_, _39114_);
  or (_39505_, _00543_, _00542_);
  and (_00544_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00545_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00546_, _00545_, _39114_);
  or (_39507_, _00546_, _00544_);
  and (_00547_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00548_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_00549_, _00548_, _39114_);
  or (_39508_, _00549_, _00547_);
  and (_00550_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00551_, _00028_, _39114_);
  or (_39509_, _00551_, _00550_);
  and (_00552_, _44110_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00553_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00554_, _00553_, _39114_);
  or (_39510_, _00554_, _00552_);
  and (_39511_, _44118_, _41991_);
  nor (_39512_, _44128_, rst);
  and (_39513_, _44124_, _41991_);
  and (_00555_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00556_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00557_, _00556_, _00555_);
  and (_39514_, _00557_, _41991_);
  and (_00558_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00559_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00560_, _00559_, _00558_);
  and (_39515_, _00560_, _41991_);
  and (_00561_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00562_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00563_, _00562_, _00561_);
  and (_39516_, _00563_, _41991_);
  and (_00564_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00565_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00566_, _00565_, _00564_);
  and (_39518_, _00566_, _41991_);
  and (_00567_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00568_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00569_, _00568_, _00567_);
  and (_39519_, _00569_, _41991_);
  and (_00570_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00571_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00572_, _00571_, _00570_);
  and (_39520_, _00572_, _41991_);
  and (_00573_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00574_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00575_, _00574_, _00573_);
  and (_39521_, _00575_, _41991_);
  and (_00576_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00577_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00578_, _00577_, _00576_);
  and (_39522_, _00578_, _41991_);
  and (_00579_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00580_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00581_, _00580_, _00579_);
  and (_39523_, _00581_, _41991_);
  and (_00582_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00583_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00584_, _00583_, _00582_);
  and (_39524_, _00584_, _41991_);
  and (_00585_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00586_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00587_, _00586_, _00585_);
  and (_39525_, _00587_, _41991_);
  and (_00588_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00589_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00590_, _00589_, _00588_);
  and (_39526_, _00590_, _41991_);
  and (_00591_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00592_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00593_, _00592_, _00591_);
  and (_39527_, _00593_, _41991_);
  and (_00594_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00595_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00596_, _00595_, _00594_);
  and (_39529_, _00596_, _41991_);
  and (_00597_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00598_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00599_, _00598_, _00597_);
  and (_39530_, _00599_, _41991_);
  and (_00600_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00601_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00602_, _00601_, _00600_);
  and (_39531_, _00602_, _41991_);
  and (_00603_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00604_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00605_, _00604_, _00603_);
  and (_39532_, _00605_, _41991_);
  and (_00606_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00607_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00608_, _00607_, _00606_);
  and (_39533_, _00608_, _41991_);
  and (_00609_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00610_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00611_, _00610_, _00609_);
  and (_39534_, _00611_, _41991_);
  and (_00612_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00613_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00614_, _00613_, _00612_);
  and (_39535_, _00614_, _41991_);
  and (_00615_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00616_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00617_, _00616_, _00615_);
  and (_39536_, _00617_, _41991_);
  and (_00618_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00619_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00620_, _00619_, _00618_);
  and (_39537_, _00620_, _41991_);
  and (_00621_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00622_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00623_, _00622_, _00621_);
  and (_39538_, _00623_, _41991_);
  and (_00624_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00625_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00626_, _00625_, _00624_);
  and (_39540_, _00626_, _41991_);
  and (_00627_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00628_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00629_, _00628_, _00627_);
  and (_39541_, _00629_, _41991_);
  and (_00630_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00631_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00632_, _00631_, _00630_);
  and (_39542_, _00632_, _41991_);
  and (_00633_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00634_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00635_, _00634_, _00633_);
  and (_39543_, _00635_, _41991_);
  and (_00636_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00637_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00638_, _00637_, _00636_);
  and (_39544_, _00638_, _41991_);
  and (_00639_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00640_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00641_, _00640_, _00639_);
  and (_39545_, _00641_, _41991_);
  and (_00642_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00643_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00644_, _00643_, _00642_);
  and (_39546_, _00644_, _41991_);
  and (_00645_, _44132_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00646_, _44134_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00647_, _00646_, _00645_);
  and (_39547_, _00647_, _41991_);
  and (_00648_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00649_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00650_, _00649_, _00648_);
  and (_39548_, _00650_, _41991_);
  and (_00651_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00652_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00653_, _00652_, _00651_);
  and (_39549_, _00653_, _41991_);
  and (_00654_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00655_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00656_, _00655_, _00654_);
  and (_39550_, _00656_, _41991_);
  and (_00657_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00658_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00659_, _00658_, _00657_);
  and (_39551_, _00659_, _41991_);
  and (_00660_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00661_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00662_, _00661_, _00660_);
  and (_39552_, _00662_, _41991_);
  and (_00663_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00664_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00665_, _00664_, _00663_);
  and (_39553_, _00665_, _41991_);
  and (_00666_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00667_, _44142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00668_, _00667_, _00666_);
  and (_39554_, _00668_, _41991_);
  and (_00669_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00670_, _40569_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00671_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00672_, _00671_, _44141_);
  and (_00673_, _00672_, _00670_);
  or (_00674_, _00673_, _00669_);
  and (_39555_, _00674_, _41991_);
  and (_00675_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00676_, _40743_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00677_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00678_, _00677_, _44141_);
  and (_00679_, _00678_, _00676_);
  or (_00680_, _00679_, _00675_);
  and (_39556_, _00680_, _41991_);
  and (_00681_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00682_, _40654_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00683_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00684_, _00683_, _44141_);
  and (_00685_, _00684_, _00682_);
  or (_00686_, _00685_, _00681_);
  and (_39557_, _00686_, _41991_);
  and (_00687_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00688_, _40536_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00689_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00690_, _00689_, _44141_);
  and (_00691_, _00690_, _00688_);
  or (_00692_, _00691_, _00687_);
  and (_39558_, _00692_, _41991_);
  and (_00693_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00694_, _40702_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00695_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00696_, _00695_, _44141_);
  and (_00697_, _00696_, _00694_);
  or (_00698_, _00697_, _00693_);
  and (_39559_, _00698_, _41991_);
  and (_00699_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00700_, _40597_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00701_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00702_, _00701_, _44141_);
  and (_00703_, _00702_, _00700_);
  or (_00704_, _00703_, _00699_);
  and (_39561_, _00704_, _41991_);
  and (_00705_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00706_, _40874_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00707_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00708_, _00707_, _44141_);
  and (_00709_, _00708_, _00706_);
  or (_00710_, _00709_, _00705_);
  and (_39562_, _00710_, _41991_);
  and (_00711_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00712_, _40459_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00713_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00714_, _00713_, _44141_);
  and (_00715_, _00714_, _00712_);
  or (_00716_, _00715_, _00711_);
  and (_39563_, _00716_, _41991_);
  and (_00717_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00718_, _00717_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00719_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _44141_);
  and (_00720_, _00719_, _41991_);
  and (_39564_, _00720_, _00718_);
  and (_00721_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00722_, _00721_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00723_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _44141_);
  and (_00724_, _00723_, _41991_);
  and (_39565_, _00724_, _00722_);
  and (_00725_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00726_, _00725_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00727_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _44141_);
  and (_00728_, _00727_, _41991_);
  and (_39566_, _00728_, _00726_);
  and (_00729_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00730_, _00729_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00731_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _44141_);
  and (_00732_, _00731_, _41991_);
  and (_39567_, _00732_, _00730_);
  and (_00733_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00734_, _00733_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00735_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _44141_);
  and (_00736_, _00735_, _41991_);
  and (_39568_, _00736_, _00734_);
  and (_00737_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00738_, _00737_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00739_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _44141_);
  and (_00740_, _00739_, _41991_);
  and (_39569_, _00740_, _00738_);
  and (_00741_, _44148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00742_, _00741_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00743_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _44141_);
  and (_00744_, _00743_, _41991_);
  and (_39570_, _00744_, _00742_);
  nand (_00745_, _44155_, _29221_);
  or (_00746_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00747_, _00746_, _41991_);
  and (_39572_, _00747_, _00745_);
  nand (_00748_, _44155_, _29894_);
  or (_00749_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00750_, _00749_, _41991_);
  and (_39573_, _00750_, _00748_);
  nand (_00751_, _44155_, _30578_);
  or (_00752_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00753_, _00752_, _41991_);
  and (_39574_, _00753_, _00751_);
  nand (_00754_, _44155_, _31327_);
  or (_00755_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00756_, _00755_, _41991_);
  and (_39575_, _00756_, _00754_);
  nand (_00757_, _44155_, _32022_);
  or (_00758_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00759_, _00758_, _41991_);
  and (_39576_, _00759_, _00757_);
  nand (_00760_, _44155_, _32842_);
  or (_00761_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00762_, _00761_, _41991_);
  and (_39577_, _00762_, _00760_);
  nand (_00763_, _44155_, _33554_);
  or (_00764_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00765_, _00764_, _41991_);
  and (_39578_, _00765_, _00763_);
  nand (_00766_, _44155_, _28011_);
  or (_00767_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00768_, _00767_, _41991_);
  and (_39579_, _00768_, _00766_);
  nand (_00769_, _44155_, _38795_);
  or (_00770_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00771_, _00770_, _41991_);
  and (_39580_, _00771_, _00769_);
  nand (_00772_, _44155_, _38823_);
  or (_00773_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00774_, _00773_, _41991_);
  and (_39581_, _00774_, _00772_);
  nand (_00775_, _44155_, _38851_);
  or (_00776_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00777_, _00776_, _41991_);
  and (_39583_, _00777_, _00775_);
  nand (_00778_, _44155_, _38880_);
  or (_00779_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00780_, _00779_, _41991_);
  and (_39584_, _00780_, _00778_);
  nand (_00781_, _44155_, _38910_);
  or (_00782_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00783_, _00782_, _41991_);
  and (_39585_, _00783_, _00781_);
  nand (_00784_, _44155_, _38940_);
  or (_00785_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00786_, _00785_, _41991_);
  and (_39586_, _00786_, _00784_);
  nand (_00787_, _44155_, _38967_);
  or (_00788_, _44155_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00789_, _00788_, _41991_);
  and (_39587_, _00789_, _00787_);
  nor (_39795_, _40499_, rst);
  nor (_00790_, _40541_, _40710_);
  and (_00791_, _00790_, _40625_);
  nor (_00792_, _40885_, _40486_);
  and (_00793_, _00792_, _00791_);
  not (_00794_, _40662_);
  nor (_00795_, _39300_, _39289_);
  and (_00796_, _39300_, _39289_);
  nor (_00797_, _00796_, _00795_);
  nor (_00798_, _39311_, _39224_);
  and (_00799_, _39311_, _39224_);
  nor (_00800_, _00799_, _00798_);
  and (_00801_, _00800_, _00797_);
  nor (_00802_, _00800_, _00797_);
  or (_00803_, _00802_, _00801_);
  and (_00804_, _39247_, _39235_);
  nor (_00805_, _39247_, _39235_);
  or (_00806_, _00805_, _00804_);
  not (_00807_, _00806_);
  nor (_00808_, _39278_, _39267_);
  and (_00809_, _39278_, _39267_);
  or (_00810_, _00809_, _00808_);
  and (_00811_, _00810_, _00807_);
  nor (_00812_, _00810_, _00807_);
  nor (_00813_, _00812_, _00811_);
  or (_00814_, _00813_, _00803_);
  nand (_00815_, _00813_, _00803_);
  and (_00816_, _00815_, _00814_);
  or (_00817_, _00816_, _00794_);
  and (_00818_, _40577_, _40776_);
  or (_00819_, _40662_, _39141_);
  and (_00820_, _00819_, _00818_);
  and (_00821_, _00820_, _00817_);
  not (_00822_, _40577_);
  and (_00823_, _00822_, _40776_);
  and (_00824_, _00794_, _39148_);
  and (_00825_, _40662_, _39055_);
  or (_00826_, _00825_, _00824_);
  and (_00827_, _00826_, _00823_);
  nor (_00828_, _40577_, _40776_);
  and (_00829_, _00828_, _40662_);
  and (_00830_, _00829_, _39130_);
  and (_00831_, _00828_, _00794_);
  and (_00832_, _00831_, _39044_);
  or (_00833_, _00832_, _00830_);
  or (_00834_, _00833_, _00827_);
  or (_00835_, _00794_, _39090_);
  nor (_00836_, _00822_, _40776_);
  or (_00837_, _40662_, _39178_);
  and (_00838_, _00837_, _00836_);
  and (_00839_, _00838_, _00835_);
  or (_00840_, _00839_, _00834_);
  or (_00841_, _00840_, _00821_);
  and (_00842_, _00841_, _00793_);
  and (_00843_, _40885_, _40626_);
  nor (_00844_, _40711_, _40486_);
  and (_00845_, _00844_, _40541_);
  and (_00846_, _00845_, _00843_);
  and (_00847_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_00848_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00849_, _00848_, _00847_);
  and (_00851_, _00849_, _00836_);
  and (_00852_, _00829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_00853_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_00854_, _00853_, _00852_);
  or (_00855_, _00854_, _00851_);
  and (_00856_, _00818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_00857_, _00823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_00858_, _00857_, _00856_);
  and (_00859_, _00858_, _40662_);
  and (_00860_, _00818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_00861_, _00823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_00862_, _00861_, _00860_);
  and (_00863_, _00862_, _00794_);
  or (_00864_, _00863_, _00859_);
  or (_00865_, _00864_, _00855_);
  and (_00866_, _00865_, _00846_);
  and (_00867_, _40885_, _40625_);
  and (_00868_, _00867_, _00844_);
  and (_00869_, _00868_, _40541_);
  and (_00870_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_00871_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_00872_, _00871_, _00870_);
  and (_00873_, _00872_, _00836_);
  and (_00874_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_00875_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_00876_, _00875_, _00874_);
  and (_00877_, _00876_, _00818_);
  or (_00878_, _00877_, _00873_);
  and (_00879_, _00829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_00880_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_00882_, _00880_, _00879_);
  and (_00883_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_00884_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_00885_, _00884_, _00883_);
  and (_00886_, _00885_, _00823_);
  or (_00887_, _00886_, _00882_);
  or (_00888_, _00887_, _00878_);
  and (_00889_, _00888_, _00869_);
  not (_00890_, _40486_);
  and (_00891_, _40885_, _00890_);
  and (_00892_, _00891_, _00791_);
  and (_00893_, _36989_, _36715_);
  not (_00894_, _00893_);
  nor (_00895_, _42670_, _36770_);
  and (_00896_, _00895_, _00894_);
  nor (_00897_, _37339_, _37295_);
  and (_00898_, _00897_, _00896_);
  nor (_00899_, _42735_, _42669_);
  and (_00900_, _00899_, _00898_);
  nor (_00901_, _42738_, _37605_);
  and (_00903_, _34518_, _36562_);
  not (_00904_, _00903_);
  and (_00905_, _00904_, _00901_);
  and (_00906_, _00905_, _43037_);
  and (_00907_, _00906_, _00900_);
  and (_00908_, _00907_, _37237_);
  nor (_00909_, _00908_, _35564_);
  and (_00910_, _43231_, p1in_reg[4]);
  and (_00911_, _43227_, p1_in[4]);
  or (_00912_, _00911_, _00910_);
  or (_00913_, _00912_, _00909_);
  not (_00914_, _00909_);
  or (_00915_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_00916_, _00915_, _00913_);
  and (_00917_, _00916_, _00794_);
  and (_00918_, _43231_, p1in_reg[0]);
  and (_00919_, _43227_, p1_in[0]);
  or (_00920_, _00919_, _00918_);
  or (_00921_, _00920_, _00909_);
  nand (_00922_, _00909_, _39673_);
  and (_00923_, _00922_, _00921_);
  and (_00924_, _00923_, _40662_);
  or (_00925_, _00924_, _00917_);
  and (_00926_, _00925_, _00818_);
  and (_00927_, _43231_, p1in_reg[3]);
  and (_00928_, _43227_, p1_in[3]);
  or (_00929_, _00928_, _00927_);
  or (_00930_, _00929_, _00909_);
  or (_00931_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00932_, _00931_, _00930_);
  and (_00933_, _00932_, _00829_);
  or (_00934_, _00933_, _00926_);
  and (_00935_, _43231_, p1in_reg[1]);
  and (_00936_, _43227_, p1_in[1]);
  or (_00937_, _00936_, _00935_);
  or (_00938_, _00937_, _00909_);
  nand (_00939_, _00909_, _39686_);
  and (_00940_, _00939_, _00938_);
  and (_00941_, _00940_, _40662_);
  and (_00942_, _43231_, p1in_reg[5]);
  and (_00943_, _43227_, p1_in[5]);
  or (_00944_, _00943_, _00942_);
  or (_00945_, _00944_, _00909_);
  or (_00946_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_00947_, _00946_, _00945_);
  and (_00948_, _00947_, _00794_);
  or (_00949_, _00948_, _00941_);
  and (_00950_, _00949_, _00823_);
  and (_00951_, _43231_, p1in_reg[2]);
  and (_00952_, _43227_, p1_in[2]);
  or (_00953_, _00952_, _00951_);
  or (_00954_, _00953_, _00909_);
  nand (_00955_, _00909_, _39699_);
  and (_00956_, _00955_, _00954_);
  and (_00957_, _00956_, _40662_);
  and (_00958_, _43231_, p1in_reg[6]);
  and (_00959_, _43227_, p1_in[6]);
  or (_00960_, _00959_, _00958_);
  or (_00961_, _00960_, _00909_);
  nand (_00962_, _00909_, _39748_);
  and (_00963_, _00962_, _00961_);
  and (_00964_, _00963_, _00794_);
  or (_00965_, _00964_, _00957_);
  and (_00966_, _00965_, _00836_);
  and (_00967_, _43231_, p1in_reg[7]);
  and (_00968_, _43227_, p1_in[7]);
  or (_00969_, _00968_, _00967_);
  or (_00970_, _00969_, _00909_);
  nand (_00971_, _00909_, _39336_);
  and (_00972_, _00971_, _00970_);
  and (_00973_, _00972_, _00831_);
  or (_00974_, _00973_, _00966_);
  or (_00975_, _00974_, _00950_);
  or (_00976_, _00975_, _00934_);
  and (_00977_, _00976_, _00892_);
  or (_00978_, _00977_, _00889_);
  or (_00979_, _00978_, _00866_);
  nor (_00980_, _40885_, _40625_);
  and (_00981_, _00790_, _00890_);
  and (_00982_, _00981_, _00980_);
  nor (_00983_, _40662_, _32875_);
  and (_00984_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_00985_, _00984_, _00983_);
  and (_00986_, _00985_, _00823_);
  and (_00987_, _00818_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_00988_, _00987_, _00794_);
  and (_00989_, _00836_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00990_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00991_, _00990_, _00989_);
  or (_00992_, _00991_, _00988_);
  and (_00993_, _00818_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_00994_, _00993_, _40662_);
  and (_00995_, _00836_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00996_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_00997_, _00996_, _00995_);
  or (_00998_, _00997_, _00994_);
  and (_00999_, _00998_, _00992_);
  or (_01000_, _00999_, _00986_);
  and (_01001_, _01000_, _00982_);
  nor (_01002_, _40540_, _40486_);
  and (_01003_, _40885_, _40711_);
  and (_01004_, _01003_, _01002_);
  and (_01005_, _01004_, _40626_);
  and (_01006_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01007_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_01008_, _01007_, _01006_);
  and (_01009_, _01008_, _00823_);
  and (_01010_, _00829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_01011_, _01010_, _01009_);
  and (_01012_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_01013_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01014_, _01013_, _01012_);
  and (_01015_, _01014_, _00836_);
  and (_01016_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_01017_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_01018_, _01017_, _01016_);
  and (_01019_, _01018_, _00818_);
  or (_01020_, _01019_, _01015_);
  and (_01021_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_01022_, _01021_, _01020_);
  or (_01023_, _01022_, _01011_);
  and (_01024_, _01023_, _01005_);
  or (_01025_, _01024_, _01001_);
  and (_01026_, _00981_, _00843_);
  and (_01027_, _43231_, p3in_reg[7]);
  and (_01028_, _43227_, p3_in[7]);
  or (_01029_, _01028_, _01027_);
  or (_01030_, _01029_, _00909_);
  nand (_01031_, _00909_, _39372_);
  and (_01032_, _01031_, _01030_);
  and (_01033_, _01032_, _00831_);
  and (_01034_, _43231_, p3in_reg[4]);
  and (_01035_, _43227_, p3_in[4]);
  or (_01036_, _01035_, _01034_);
  or (_01037_, _01036_, _00909_);
  or (_01038_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_01039_, _01038_, _01037_);
  and (_01040_, _01039_, _00794_);
  and (_01041_, _43231_, p3in_reg[0]);
  and (_01042_, _43227_, p3_in[0]);
  or (_01043_, _01042_, _01041_);
  or (_01044_, _01043_, _00909_);
  nand (_01045_, _00909_, _39853_);
  and (_01046_, _01045_, _01044_);
  and (_01047_, _01046_, _40662_);
  or (_01048_, _01047_, _01040_);
  and (_01049_, _01048_, _00818_);
  and (_01050_, _43231_, p3in_reg[3]);
  and (_01051_, _43227_, p3_in[3]);
  or (_01052_, _01051_, _01050_);
  or (_01053_, _01052_, _00909_);
  or (_01054_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_01055_, _01054_, _01053_);
  and (_01056_, _01055_, _00829_);
  or (_01057_, _01056_, _01049_);
  or (_01058_, _01057_, _01033_);
  and (_01059_, _43231_, p3in_reg[2]);
  and (_01060_, _43227_, p3_in[2]);
  or (_01061_, _01060_, _01059_);
  or (_01062_, _01061_, _00909_);
  nand (_01063_, _00909_, _39879_);
  and (_01064_, _01063_, _01062_);
  and (_01065_, _01064_, _40662_);
  and (_01066_, _43231_, p3in_reg[6]);
  and (_01067_, _43227_, p3_in[6]);
  or (_01068_, _01067_, _01066_);
  or (_01069_, _01068_, _00909_);
  nand (_01070_, _00909_, _39935_);
  and (_01071_, _01070_, _01069_);
  and (_01072_, _01071_, _00794_);
  or (_01073_, _01072_, _01065_);
  and (_01074_, _01073_, _00836_);
  and (_01075_, _43231_, p3in_reg[1]);
  and (_01076_, _43227_, p3_in[1]);
  or (_01077_, _01076_, _01075_);
  or (_01078_, _01077_, _00909_);
  nand (_01079_, _00909_, _39866_);
  and (_01080_, _01079_, _01078_);
  and (_01081_, _01080_, _40662_);
  and (_01082_, _43231_, p3in_reg[5]);
  and (_01083_, _43227_, p3_in[5]);
  or (_01084_, _01083_, _01082_);
  or (_01085_, _01084_, _00909_);
  or (_01086_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01087_, _01086_, _01085_);
  and (_01088_, _01087_, _00794_);
  or (_01089_, _01088_, _01081_);
  and (_01090_, _01089_, _00823_);
  or (_01091_, _01090_, _01074_);
  or (_01092_, _01091_, _01058_);
  and (_01093_, _01092_, _01026_);
  and (_01094_, _00868_, _40540_);
  and (_01095_, _43231_, p0in_reg[3]);
  and (_01096_, _43227_, p0_in[3]);
  or (_01097_, _01096_, _01095_);
  or (_01098_, _01097_, _00909_);
  nand (_01099_, _00909_, _39614_);
  and (_01100_, _01099_, _01098_);
  and (_01101_, _01100_, _00829_);
  and (_01102_, _43231_, p0in_reg[2]);
  and (_01103_, _43227_, p0_in[2]);
  or (_01104_, _01103_, _01102_);
  or (_01105_, _01104_, _00909_);
  nand (_01106_, _00909_, _39610_);
  and (_01107_, _01106_, _01105_);
  and (_01108_, _01107_, _40662_);
  and (_01109_, _43231_, p0in_reg[6]);
  and (_01110_, _43227_, p0_in[6]);
  or (_01111_, _01110_, _01109_);
  or (_01112_, _01111_, _00909_);
  nand (_01113_, _00909_, _39664_);
  and (_01114_, _01113_, _01112_);
  and (_01115_, _01114_, _00794_);
  or (_01116_, _01115_, _01108_);
  and (_01117_, _01116_, _00836_);
  and (_01118_, _43231_, p0in_reg[7]);
  and (_01119_, _43227_, p0_in[7]);
  or (_01120_, _01119_, _01118_);
  or (_01121_, _01120_, _00909_);
  nand (_01122_, _00909_, _39322_);
  and (_01123_, _01122_, _01121_);
  and (_01124_, _01123_, _00831_);
  or (_01125_, _01124_, _01117_);
  or (_01126_, _01125_, _01101_);
  and (_01127_, _43231_, p0in_reg[0]);
  and (_01128_, _43227_, p0_in[0]);
  or (_01129_, _01128_, _01127_);
  or (_01130_, _01129_, _00909_);
  nand (_01131_, _00909_, _39419_);
  and (_01132_, _01131_, _01130_);
  and (_01133_, _01132_, _00818_);
  and (_01134_, _43231_, p0in_reg[1]);
  and (_01135_, _43227_, p0_in[1]);
  or (_01136_, _01135_, _01134_);
  or (_01137_, _01136_, _00909_);
  nand (_01138_, _00909_, _39594_);
  and (_01139_, _01138_, _01137_);
  and (_01140_, _01139_, _00823_);
  or (_01141_, _01140_, _01133_);
  and (_01142_, _01141_, _40662_);
  and (_01143_, _43231_, p0in_reg[4]);
  and (_01144_, _43227_, p0_in[4]);
  or (_01145_, _01144_, _01143_);
  or (_01146_, _01145_, _00909_);
  or (_01147_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01148_, _01147_, _01146_);
  and (_01149_, _01148_, _00818_);
  and (_01150_, _43231_, p0in_reg[5]);
  and (_01151_, _43227_, p0_in[5]);
  or (_01152_, _01151_, _01150_);
  or (_01153_, _01152_, _00909_);
  or (_01154_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01155_, _01154_, _01153_);
  and (_01156_, _01155_, _00823_);
  or (_01157_, _01156_, _01149_);
  and (_01158_, _01157_, _00794_);
  or (_01159_, _01158_, _01142_);
  or (_01160_, _01159_, _01126_);
  and (_01161_, _01160_, _01094_);
  or (_01162_, _01161_, _01093_);
  or (_01163_, _01162_, _01025_);
  or (_01164_, _01163_, _00979_);
  and (_01165_, _00845_, _40885_);
  or (_01166_, _01165_, _00793_);
  nor (_01167_, _01166_, _00982_);
  and (_01168_, _00844_, _40540_);
  and (_01169_, _01168_, _00980_);
  not (_01170_, _01169_);
  nor (_01171_, _40541_, _40486_);
  and (_01172_, _01171_, _40885_);
  nor (_01173_, _01172_, _01004_);
  and (_01174_, _01173_, _01170_);
  and (_01175_, _01174_, _01167_);
  nand (_01176_, _43266_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_01177_, _01176_, _01175_);
  and (_01178_, _43231_, p2in_reg[7]);
  and (_01179_, _43227_, p2_in[7]);
  or (_01180_, _01179_, _01178_);
  or (_01181_, _01180_, _00909_);
  nand (_01182_, _00909_, _39354_);
  and (_01183_, _01182_, _01181_);
  and (_01184_, _01183_, _00831_);
  and (_01185_, _43231_, p2in_reg[4]);
  and (_01186_, _43227_, p2_in[4]);
  or (_01187_, _01186_, _01185_);
  or (_01188_, _01187_, _00909_);
  or (_01189_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_01190_, _01189_, _01188_);
  and (_01191_, _01190_, _00794_);
  and (_01192_, _43231_, p2in_reg[0]);
  and (_01193_, _43227_, p2_in[0]);
  or (_01194_, _01193_, _01192_);
  or (_01195_, _01194_, _00909_);
  nand (_01196_, _00909_, _39760_);
  and (_01197_, _01196_, _01195_);
  and (_01198_, _01197_, _40662_);
  or (_01199_, _01198_, _01191_);
  and (_01200_, _01199_, _00818_);
  and (_01201_, _43231_, p2in_reg[3]);
  and (_01202_, _43227_, p2_in[3]);
  or (_01203_, _01202_, _01201_);
  or (_01204_, _01203_, _00909_);
  or (_01205_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_01206_, _01205_, _01204_);
  and (_01207_, _01206_, _00829_);
  or (_01208_, _01207_, _01200_);
  or (_01209_, _01208_, _01184_);
  and (_01210_, _43231_, p2in_reg[2]);
  and (_01211_, _43227_, p2_in[2]);
  or (_01212_, _01211_, _01210_);
  or (_01213_, _01212_, _00909_);
  nand (_01214_, _00909_, _39786_);
  and (_01215_, _01214_, _01213_);
  and (_01216_, _01215_, _40662_);
  and (_01217_, _43231_, p2in_reg[6]);
  and (_01218_, _43227_, p2_in[6]);
  or (_01219_, _01218_, _01217_);
  or (_01220_, _01219_, _00909_);
  nand (_01221_, _00909_, _39840_);
  and (_01222_, _01221_, _01220_);
  and (_01223_, _01222_, _00794_);
  or (_01224_, _01223_, _01216_);
  and (_01225_, _01224_, _00836_);
  and (_01226_, _43231_, p2in_reg[1]);
  and (_01227_, _43227_, p2_in[1]);
  or (_01228_, _01227_, _01226_);
  or (_01229_, _01228_, _00909_);
  nand (_01230_, _00909_, _39773_);
  and (_01231_, _01230_, _01229_);
  and (_01232_, _01231_, _40662_);
  and (_01233_, _43231_, p2in_reg[5]);
  and (_01234_, _43227_, p2_in[5]);
  or (_01235_, _01234_, _01233_);
  or (_01236_, _01235_, _00909_);
  or (_01237_, _00914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01238_, _01237_, _01236_);
  and (_01239_, _01238_, _00794_);
  or (_01240_, _01239_, _01232_);
  and (_01241_, _01240_, _00823_);
  or (_01242_, _01241_, _01225_);
  or (_01243_, _01242_, _01209_);
  and (_01244_, _01243_, _00843_);
  not (_01245_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_01246_, _40662_, _01245_);
  and (_01247_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_01248_, _01247_, _01246_);
  and (_01249_, _01248_, _00836_);
  and (_01250_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01251_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01252_, _01251_, _01250_);
  and (_01253_, _01252_, _00818_);
  or (_01254_, _01253_, _01249_);
  and (_01255_, _00829_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01256_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01257_, _01256_, _01255_);
  and (_01258_, _00794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01259_, _40662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_01260_, _01259_, _01258_);
  and (_01261_, _01260_, _00823_);
  or (_01262_, _01261_, _01257_);
  or (_01263_, _01262_, _01254_);
  and (_01264_, _01263_, _00980_);
  or (_01265_, _01264_, _01244_);
  nand (_01266_, _01265_, _01168_);
  nand (_01267_, _01266_, _01177_);
  or (_01268_, _01267_, _01164_);
  or (_01269_, _01268_, _00842_);
  and (_01270_, _01169_, _39200_);
  nor (_01271_, _01177_, _29308_);
  nor (_01272_, _01271_, _01270_);
  and (_01273_, _01272_, _01269_);
  or (_01274_, _00794_, _39235_);
  or (_01275_, _40662_, _39289_);
  and (_01276_, _01275_, _00818_);
  and (_01277_, _01276_, _01274_);
  or (_01278_, _40662_, _39311_);
  nand (_01279_, _40662_, _39267_);
  and (_01280_, _01279_, _00836_);
  and (_01281_, _01280_, _01278_);
  or (_01282_, _40662_, _39300_);
  or (_01283_, _00794_, _39247_);
  and (_01284_, _01283_, _00823_);
  and (_01285_, _01284_, _01282_);
  not (_01286_, _00829_);
  nor (_01287_, _01286_, _39278_);
  and (_01288_, _00831_, _39224_);
  or (_01289_, _01288_, _01287_);
  or (_01290_, _01289_, _01285_);
  or (_01291_, _01290_, _01281_);
  or (_01292_, _01291_, _01277_);
  and (_01293_, _01292_, _01270_);
  not (_01294_, _39030_);
  and (_01295_, _01172_, _00914_);
  nor (_01296_, _01295_, _01294_);
  and (_01297_, _01296_, _43253_);
  not (_01298_, _01297_);
  nor (_01299_, _01298_, _01175_);
  or (_01300_, _01299_, _01293_);
  or (_01301_, _01300_, _01273_);
  not (_01302_, _38194_);
  and (_01303_, _00831_, _01302_);
  nor (_01304_, _40662_, _38326_);
  nor (_01305_, _00794_, _38592_);
  or (_01306_, _01305_, _01304_);
  and (_01307_, _01306_, _00836_);
  nor (_01308_, _40662_, _38477_);
  and (_01309_, _40662_, _38608_);
  or (_01310_, _01309_, _01308_);
  and (_01311_, _01310_, _00818_);
  or (_01312_, _01311_, _01307_);
  nor (_01313_, _01286_, _38552_);
  nor (_01314_, _40662_, _38402_);
  and (_01315_, _40662_, _40741_);
  or (_01316_, _01315_, _01314_);
  and (_01317_, _01316_, _00823_);
  or (_01318_, _01317_, _01313_);
  or (_01319_, _01318_, _01312_);
  nor (_01320_, _01319_, _01303_);
  nand (_01321_, _01320_, _01299_);
  and (_01322_, _01321_, _41991_);
  and (_39826_, _01322_, _01301_);
  and (_01323_, _01094_, _00829_);
  and (_01324_, _01323_, _38674_);
  and (_01325_, _00818_, _40662_);
  and (_01326_, _01325_, _00793_);
  and (_01327_, _01326_, _39035_);
  nor (_01328_, _01327_, _01324_);
  nor (_01329_, _01328_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_01330_, _01329_);
  not (_01331_, _39001_);
  nor (_01332_, _00831_, _01331_);
  and (_01333_, _01332_, _43253_);
  and (_01334_, _01325_, _01169_);
  and (_01335_, _01334_, _39215_);
  nor (_01336_, _01335_, _01333_);
  and (_01337_, _01336_, _43269_);
  and (_01338_, _01337_, _01330_);
  and (_01339_, _40540_, _40662_);
  and (_01340_, _01339_, _00836_);
  and (_01341_, _01340_, _00868_);
  and (_01342_, _01341_, _38674_);
  or (_01343_, _01342_, rst);
  nor (_39827_, _01343_, _01338_);
  not (_01344_, _01342_);
  and (_01345_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_01346_, _40710_, _40625_);
  and (_01347_, _01346_, _00891_);
  and (_01348_, _01325_, _40541_);
  and (_01349_, _01348_, _01347_);
  and (_01350_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_01351_, _01350_, _01345_);
  and (_01352_, _01348_, _00868_);
  and (_01353_, _01352_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_01354_, _00843_, _00844_);
  and (_01355_, _01348_, _01354_);
  and (_01356_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_01357_, _01356_, _01353_);
  or (_01358_, _01357_, _01351_);
  and (_01359_, _01339_, _00818_);
  and (_01360_, _01346_, _00792_);
  and (_01361_, _01360_, _01359_);
  and (_01362_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01363_, _01339_, _00828_);
  and (_01364_, _01363_, _00868_);
  and (_01365_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01366_, _01365_, _01362_);
  and (_01367_, _01339_, _00823_);
  and (_01368_, _01367_, _00868_);
  and (_01369_, _01368_, _40425_);
  and (_01370_, _01347_, _01359_);
  and (_01371_, _01370_, _01032_);
  or (_01372_, _01371_, _01369_);
  or (_01373_, _01372_, _01366_);
  or (_01374_, _01373_, _01358_);
  and (_01375_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01376_, _01359_, _01354_);
  and (_01377_, _01376_, _01183_);
  and (_01378_, _40711_, _40625_);
  and (_01379_, _00891_, _01378_);
  and (_01380_, _01379_, _01359_);
  and (_01381_, _01380_, _00972_);
  or (_01382_, _01381_, _01377_);
  and (_01383_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01384_, _01359_, _00868_);
  and (_01385_, _01384_, _01123_);
  or (_01386_, _01385_, _01383_);
  or (_01387_, _01386_, _01382_);
  or (_01388_, _01387_, _01375_);
  or (_01389_, _01388_, _01374_);
  and (_01390_, _01389_, _01338_);
  nor (_01391_, _01338_, _17486_);
  or (_01392_, _01391_, _01390_);
  and (_01393_, _01392_, _01344_);
  nor (_01394_, _01344_, _28011_);
  or (_01395_, _01394_, _01393_);
  and (_39828_, _01395_, _41991_);
  and (_01398_, _01326_, _00816_);
  and (_01400_, _01325_, _00846_);
  and (_01402_, _01400_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01404_, _01325_, _00869_);
  and (_01406_, _01404_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01408_, _01325_, _01094_);
  and (_01409_, _01408_, _01132_);
  or (_01410_, _01409_, _01406_);
  or (_01411_, _01410_, _01402_);
  and (_01412_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_01413_, _01376_, _01197_);
  and (_01414_, _01325_, _00892_);
  and (_01416_, _01414_, _00923_);
  or (_01417_, _01416_, _01413_);
  or (_01419_, _01417_, _01412_);
  and (_01420_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01421_, _01370_, _01046_);
  or (_01423_, _01421_, _01420_);
  and (_01424_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01425_, _01368_, _40573_);
  or (_01427_, _01425_, _01424_);
  or (_01428_, _01427_, _01423_);
  and (_01429_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_01431_, _01323_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_01432_, _01431_, _01429_);
  or (_01433_, _01432_, _01428_);
  or (_01435_, _01433_, _01419_);
  nor (_01436_, _01435_, _01411_);
  nand (_01437_, _01436_, _01338_);
  or (_01439_, _01437_, _01398_);
  or (_01440_, _01338_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_01441_, _01440_, _01439_);
  or (_01443_, _01441_, _01342_);
  nand (_01444_, _01342_, _29221_);
  and (_01445_, _01444_, _41991_);
  and (_39891_, _01445_, _01443_);
  and (_01447_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_01448_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_01449_, _01448_, _01447_);
  and (_01450_, _01352_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_01451_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_01452_, _01451_, _01450_);
  or (_01453_, _01452_, _01449_);
  and (_01454_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01455_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_01456_, _01455_, _01454_);
  and (_01457_, _01370_, _01080_);
  and (_01458_, _01368_, _40731_);
  or (_01459_, _01458_, _01457_);
  or (_01460_, _01459_, _01456_);
  or (_01461_, _01460_, _01453_);
  and (_01462_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01463_, _01376_, _01231_);
  and (_01464_, _01380_, _00940_);
  or (_01465_, _01464_, _01463_);
  and (_01466_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_01468_, _01384_, _01139_);
  or (_01469_, _01468_, _01466_);
  or (_01471_, _01469_, _01465_);
  or (_01472_, _01471_, _01462_);
  or (_01473_, _01472_, _01461_);
  and (_01475_, _01473_, _01338_);
  nor (_01476_, _01338_, _17312_);
  or (_01477_, _01476_, _01475_);
  and (_01479_, _01477_, _01344_);
  nor (_01480_, _01344_, _29894_);
  or (_01481_, _01480_, _01479_);
  and (_39892_, _01481_, _41991_);
  and (_01483_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_01484_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01486_, _01484_, _01483_);
  and (_01487_, _01352_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_01488_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01490_, _01488_, _01487_);
  or (_01491_, _01490_, _01486_);
  and (_01492_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01494_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_01495_, _01494_, _01492_);
  and (_01496_, _01368_, _40658_);
  and (_01498_, _01370_, _01064_);
  or (_01499_, _01498_, _01496_);
  or (_01500_, _01499_, _01495_);
  or (_01501_, _01500_, _01491_);
  and (_01502_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01503_, _01376_, _01215_);
  and (_01504_, _01380_, _00956_);
  or (_01505_, _01504_, _01503_);
  and (_01506_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_01507_, _01384_, _01107_);
  or (_01508_, _01507_, _01506_);
  or (_01509_, _01508_, _01505_);
  or (_01510_, _01509_, _01502_);
  or (_01511_, _01510_, _01501_);
  and (_01512_, _01511_, _01338_);
  nor (_01513_, _01338_, _15963_);
  or (_01514_, _01513_, _01512_);
  and (_01515_, _01514_, _01344_);
  nor (_01516_, _01344_, _30578_);
  or (_01517_, _01516_, _01515_);
  and (_39893_, _01517_, _41991_);
  and (_01519_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_01520_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_01522_, _01520_, _01519_);
  and (_01523_, _01352_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_01524_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_01526_, _01524_, _01523_);
  or (_01527_, _01526_, _01522_);
  and (_01528_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01530_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_01531_, _01530_, _01528_);
  and (_01532_, _01370_, _01055_);
  and (_01534_, _01368_, _40502_);
  or (_01535_, _01534_, _01532_);
  or (_01536_, _01535_, _01531_);
  or (_01538_, _01536_, _01527_);
  and (_01539_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01540_, _01376_, _01206_);
  and (_01542_, _01380_, _00932_);
  or (_01543_, _01542_, _01540_);
  and (_01544_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_01546_, _01384_, _01100_);
  or (_01547_, _01546_, _01544_);
  or (_01548_, _01547_, _01543_);
  or (_01550_, _01548_, _01539_);
  or (_01551_, _01550_, _01538_);
  and (_01552_, _01551_, _01338_);
  nor (_01553_, _01338_, _16995_);
  or (_01554_, _01553_, _01552_);
  and (_01555_, _01554_, _01344_);
  nor (_01556_, _01344_, _31327_);
  or (_01557_, _01556_, _01555_);
  and (_39894_, _01557_, _41991_);
  and (_01558_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01559_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01560_, _01559_, _01558_);
  and (_01561_, _01352_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01562_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01563_, _01562_, _01561_);
  or (_01564_, _01563_, _01560_);
  and (_01565_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01566_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01567_, _01566_, _01565_);
  and (_01568_, _01368_, _40706_);
  and (_01569_, _01370_, _01039_);
  or (_01571_, _01569_, _01568_);
  or (_01572_, _01571_, _01567_);
  or (_01574_, _01572_, _01564_);
  and (_01575_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01576_, _01376_, _01190_);
  and (_01578_, _01380_, _00916_);
  or (_01579_, _01578_, _01576_);
  and (_01580_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01582_, _01384_, _01148_);
  or (_01583_, _01582_, _01580_);
  or (_01584_, _01583_, _01579_);
  or (_01586_, _01584_, _01575_);
  or (_01587_, _01586_, _01574_);
  and (_01588_, _01587_, _01338_);
  nor (_01590_, _01338_, _16161_);
  or (_01591_, _01590_, _01588_);
  and (_01592_, _01591_, _01344_);
  nor (_01594_, _01344_, _32022_);
  or (_01595_, _01594_, _01592_);
  and (_39895_, _01595_, _41991_);
  and (_01597_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01598_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_01599_, _01598_, _01597_);
  and (_01601_, _01352_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_01602_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01603_, _01602_, _01601_);
  or (_01604_, _01603_, _01599_);
  and (_01605_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01606_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_01607_, _01606_, _01605_);
  and (_01608_, _01370_, _01087_);
  and (_01609_, _01368_, _40603_);
  or (_01610_, _01609_, _01608_);
  or (_01611_, _01610_, _01607_);
  or (_01612_, _01611_, _01604_);
  and (_01613_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01614_, _01376_, _01238_);
  and (_01615_, _01380_, _00947_);
  or (_01616_, _01615_, _01614_);
  and (_01617_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01618_, _01384_, _01155_);
  or (_01619_, _01618_, _01617_);
  or (_01620_, _01619_, _01616_);
  or (_01621_, _01620_, _01613_);
  or (_01623_, _01621_, _01612_);
  and (_01624_, _01623_, _01338_);
  nor (_01626_, _01338_, _17148_);
  or (_01627_, _01626_, _01624_);
  and (_01628_, _01627_, _01344_);
  nor (_01630_, _01344_, _32842_);
  or (_01631_, _01630_, _01628_);
  and (_39896_, _01631_, _41991_);
  and (_01633_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_01634_, _01341_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_01635_, _01634_, _01633_);
  and (_01637_, _01352_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_01638_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_01639_, _01638_, _01637_);
  or (_01641_, _01639_, _01635_);
  and (_01642_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01643_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_01645_, _01643_, _01642_);
  and (_01646_, _01370_, _01071_);
  and (_01647_, _01368_, _40789_);
  or (_01649_, _01647_, _01646_);
  or (_01650_, _01649_, _01645_);
  or (_01651_, _01650_, _01641_);
  and (_01653_, _01334_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01654_, _01376_, _01222_);
  and (_01655_, _01380_, _00963_);
  or (_01656_, _01655_, _01654_);
  and (_01657_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01658_, _01384_, _01114_);
  or (_01659_, _01658_, _01657_);
  or (_01660_, _01659_, _01656_);
  or (_01661_, _01660_, _01653_);
  or (_01662_, _01661_, _01651_);
  and (_01663_, _01662_, _01338_);
  nor (_01664_, _01338_, _16500_);
  or (_01665_, _01664_, _01663_);
  and (_01666_, _01665_, _01344_);
  nor (_01667_, _01344_, _33554_);
  or (_01668_, _01667_, _01666_);
  and (_39897_, _01668_, _41991_);
  and (_39942_, _40923_, _41991_);
  and (_39943_, _41039_, _41991_);
  nor (_39945_, _40662_, rst);
  and (_39960_, _41057_, _41991_);
  and (_39961_, _41072_, _41991_);
  and (_39962_, _41083_, _41991_);
  and (_39963_, _41093_, _41991_);
  and (_39964_, _41102_, _41991_);
  and (_39965_, _41113_, _41991_);
  and (_39966_, _41124_, _41991_);
  nor (_39967_, _40577_, rst);
  nor (_39968_, _40776_, rst);
  not (_01673_, _41913_);
  nor (_01674_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01676_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01677_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01676_);
  nor (_01678_, _01677_, _01674_);
  nor (_01680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01681_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01676_);
  nor (_01682_, _01681_, _01680_);
  not (_01684_, _01682_);
  nor (_01685_, _01684_, _01678_);
  nor (_01686_, _00169_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01688_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01676_);
  nor (_01689_, _01688_, _01686_);
  nor (_01690_, _00149_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01692_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01676_);
  nor (_01693_, _01692_, _01690_);
  not (_01694_, _01693_);
  nor (_01695_, _01694_, _01689_);
  nor (_01696_, _01682_, _01678_);
  not (_01697_, _01696_);
  and (_01698_, _01693_, _01697_);
  nor (_01699_, _01689_, _01697_);
  nor (_01700_, _01699_, _01698_);
  nor (_01701_, _01700_, _01695_);
  and (_01702_, _01701_, _01685_);
  and (_01703_, _01702_, _01673_);
  not (_01704_, _41961_);
  and (_01705_, _01682_, _01678_);
  and (_01706_, _01701_, _01705_);
  and (_01707_, _01706_, _01704_);
  or (_01708_, _01707_, _01703_);
  not (_01709_, _41872_);
  and (_01710_, _01684_, _01678_);
  and (_01711_, _01710_, _01701_);
  and (_01712_, _01711_, _01709_);
  not (_01714_, _42256_);
  and (_01715_, _01695_, _01685_);
  and (_01717_, _01715_, _01714_);
  not (_01718_, _42297_);
  and (_01719_, _01695_, _01705_);
  and (_01721_, _01719_, _01718_);
  or (_01722_, _01721_, _01717_);
  not (_01723_, _42010_);
  not (_01725_, _01689_);
  nor (_01726_, _01693_, _01697_);
  and (_01727_, _01726_, _01725_);
  and (_01729_, _01727_, _01723_);
  not (_01730_, _42215_);
  and (_01731_, _01710_, _01695_);
  and (_01733_, _01731_, _01730_);
  or (_01734_, _01733_, _01729_);
  or (_01735_, _01734_, _01722_);
  or (_01737_, _01735_, _01712_);
  or (_01738_, _01737_, _01708_);
  not (_01739_, _42051_);
  nor (_01741_, _01726_, _01698_);
  and (_01742_, _01741_, _01725_);
  and (_01743_, _01742_, _01710_);
  and (_01745_, _01743_, _01739_);
  not (_01746_, _42092_);
  and (_01747_, _01742_, _01685_);
  and (_01748_, _01747_, _01746_);
  not (_01749_, _42420_);
  and (_01750_, _01741_, _01689_);
  and (_01751_, _01750_, _01685_);
  and (_01752_, _01751_, _01749_);
  or (_01753_, _01752_, _01748_);
  or (_01754_, _01753_, _01745_);
  not (_01755_, _42379_);
  and (_01756_, _01750_, _01710_);
  and (_01757_, _01756_, _01755_);
  not (_01758_, _42502_);
  and (_01759_, _01693_, _01696_);
  and (_01760_, _01759_, _01689_);
  and (_01761_, _01760_, _01758_);
  not (_01762_, _42174_);
  and (_01763_, _01695_, _01696_);
  and (_01764_, _01763_, _01762_);
  not (_01765_, _42338_);
  and (_01767_, _01726_, _01689_);
  and (_01768_, _01767_, _01765_);
  or (_01770_, _01768_, _01764_);
  or (_01771_, _01770_, _01761_);
  or (_01772_, _01771_, _01757_);
  not (_01774_, _42133_);
  and (_01775_, _01742_, _01705_);
  and (_01776_, _01775_, _01774_);
  not (_01778_, _42461_);
  and (_01779_, _01750_, _01705_);
  and (_01780_, _01779_, _01778_);
  or (_01782_, _01780_, _01776_);
  or (_01783_, _01782_, _01772_);
  or (_01784_, _01783_, _01754_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01784_, _01738_);
  and (_01786_, _01702_, _01758_);
  and (_01787_, _01719_, _01730_);
  and (_01789_, _01715_, _01762_);
  or (_01790_, _01789_, _01787_);
  and (_01791_, _01727_, _01673_);
  and (_01793_, _01731_, _01774_);
  or (_01794_, _01793_, _01791_);
  or (_01795_, _01794_, _01790_);
  or (_01797_, _01795_, _01786_);
  and (_01798_, _01711_, _01778_);
  and (_01799_, _01706_, _01709_);
  or (_01800_, _01799_, _01798_);
  or (_01801_, _01800_, _01797_);
  and (_01802_, _01779_, _01755_);
  and (_01803_, _01756_, _01718_);
  and (_01804_, _01743_, _01704_);
  or (_01805_, _01804_, _01803_);
  or (_01806_, _01805_, _01802_);
  and (_01807_, _01775_, _01739_);
  and (_01808_, _01747_, _01723_);
  or (_01809_, _01808_, _01807_);
  and (_01810_, _01751_, _01765_);
  and (_01811_, _01767_, _01714_);
  and (_01812_, _01760_, _01749_);
  and (_01813_, _01763_, _01746_);
  or (_01814_, _01813_, _01812_);
  or (_01815_, _01814_, _01811_);
  or (_01816_, _01815_, _01810_);
  or (_01817_, _01816_, _01809_);
  or (_01819_, _01817_, _01806_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01819_, _01801_);
  and (_01821_, _01702_, _01709_);
  and (_01822_, _01731_, _01762_);
  and (_01823_, _01715_, _01730_);
  or (_01825_, _01823_, _01822_);
  and (_01826_, _01727_, _01704_);
  and (_01827_, _01719_, _01714_);
  or (_01829_, _01827_, _01826_);
  or (_01830_, _01829_, _01825_);
  or (_01831_, _01830_, _01821_);
  and (_01833_, _01711_, _01758_);
  and (_01834_, _01706_, _01673_);
  or (_01835_, _01834_, _01833_);
  or (_01837_, _01835_, _01831_);
  and (_01838_, _01747_, _01739_);
  and (_01839_, _01775_, _01746_);
  and (_01841_, _01756_, _01765_);
  or (_01842_, _01841_, _01839_);
  or (_01843_, _01842_, _01838_);
  and (_01845_, _01779_, _01749_);
  and (_01846_, _01763_, _01774_);
  and (_01847_, _01767_, _01718_);
  and (_01849_, _01760_, _01778_);
  or (_01850_, _01849_, _01847_);
  or (_01851_, _01850_, _01846_);
  or (_01852_, _01851_, _01845_);
  and (_01853_, _01743_, _01723_);
  and (_01854_, _01751_, _01755_);
  or (_01855_, _01854_, _01853_);
  or (_01856_, _01855_, _01852_);
  or (_01857_, _01856_, _01843_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01857_, _01837_);
  and (_01858_, _01743_, _01673_);
  and (_01859_, _01727_, _01709_);
  and (_01860_, _01747_, _01704_);
  or (_01861_, _01860_, _01859_);
  or (_01862_, _01861_, _01858_);
  and (_01863_, _01706_, _01758_);
  and (_01864_, _01702_, _01778_);
  or (_01865_, _01864_, _01863_);
  and (_01866_, _01711_, _01749_);
  or (_01867_, _01866_, _01865_);
  or (_01868_, _01867_, _01862_);
  and (_01870_, _01760_, _01755_);
  and (_01871_, _01715_, _01774_);
  and (_01873_, _01731_, _01746_);
  or (_01874_, _01873_, _01871_);
  and (_01875_, _01775_, _01723_);
  and (_01877_, _01763_, _01739_);
  or (_01878_, _01877_, _01875_);
  or (_01879_, _01878_, _01874_);
  and (_01881_, _01756_, _01714_);
  and (_01882_, _01719_, _01762_);
  and (_01883_, _01767_, _01730_);
  or (_01885_, _01883_, _01882_);
  or (_01886_, _01885_, _01881_);
  and (_01887_, _01779_, _01765_);
  and (_01889_, _01751_, _01718_);
  or (_01890_, _01889_, _01887_);
  or (_01891_, _01890_, _01886_);
  or (_01893_, _01891_, _01879_);
  or (_01894_, _01893_, _01870_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01894_, _01868_);
  not (_01896_, _42425_);
  and (_01897_, _01711_, _01896_);
  not (_01898_, _42466_);
  and (_01900_, _01702_, _01898_);
  or (_01901_, _01900_, _01897_);
  not (_01902_, _42507_);
  and (_01903_, _01706_, _01902_);
  not (_01904_, _42179_);
  and (_01905_, _01719_, _01904_);
  not (_01906_, _42138_);
  and (_01907_, _01715_, _01906_);
  or (_01908_, _01907_, _01905_);
  not (_01909_, _42097_);
  and (_01910_, _01731_, _01909_);
  not (_01911_, _41877_);
  and (_01912_, _01727_, _01911_);
  or (_01913_, _01912_, _01910_);
  or (_01914_, _01913_, _01908_);
  or (_01915_, _01914_, _01903_);
  or (_01916_, _01915_, _01901_);
  not (_01917_, _42343_);
  and (_01918_, _01779_, _01917_);
  not (_01919_, _42261_);
  and (_01920_, _01756_, _01919_);
  not (_01922_, _41966_);
  and (_01923_, _01747_, _01922_);
  or (_01925_, _01923_, _01920_);
  or (_01926_, _01925_, _01918_);
  not (_01927_, _41918_);
  and (_01929_, _01743_, _01927_);
  not (_01930_, _42056_);
  and (_01931_, _01763_, _01930_);
  not (_01933_, _42384_);
  and (_01934_, _01760_, _01933_);
  not (_01935_, _42220_);
  and (_01937_, _01767_, _01935_);
  or (_01938_, _01937_, _01934_);
  or (_01939_, _01938_, _01931_);
  or (_01941_, _01939_, _01929_);
  not (_01942_, _42302_);
  and (_01943_, _01751_, _01942_);
  not (_01945_, _42015_);
  and (_01946_, _01775_, _01945_);
  or (_01947_, _01946_, _01943_);
  or (_01949_, _01947_, _01941_);
  or (_01950_, _01949_, _01926_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _01950_, _01916_);
  not (_01952_, _42430_);
  and (_01953_, _01711_, _01952_);
  not (_01954_, _42471_);
  and (_01955_, _01702_, _01954_);
  or (_01956_, _01955_, _01953_);
  not (_01957_, _42512_);
  and (_01958_, _01706_, _01957_);
  not (_01959_, _42102_);
  and (_01960_, _01731_, _01959_);
  not (_01961_, _42143_);
  and (_01962_, _01715_, _01961_);
  or (_01963_, _01962_, _01960_);
  not (_01964_, _41882_);
  and (_01965_, _01727_, _01964_);
  not (_01966_, _42184_);
  and (_01967_, _01719_, _01966_);
  or (_01968_, _01967_, _01965_);
  or (_01969_, _01968_, _01963_);
  or (_01970_, _01969_, _01958_);
  or (_01971_, _01970_, _01956_);
  not (_01972_, _42266_);
  and (_01974_, _01756_, _01972_);
  not (_01975_, _41923_);
  and (_01977_, _01743_, _01975_);
  not (_01978_, _42348_);
  and (_01979_, _01779_, _01978_);
  or (_01981_, _01979_, _01977_);
  or (_01982_, _01981_, _01974_);
  not (_01983_, _42307_);
  and (_01985_, _01751_, _01983_);
  not (_01986_, _42389_);
  and (_01987_, _01760_, _01986_);
  not (_01989_, _42061_);
  and (_01990_, _01763_, _01989_);
  not (_01991_, _42225_);
  and (_01993_, _01767_, _01991_);
  or (_01994_, _01993_, _01990_);
  or (_01995_, _01994_, _01987_);
  or (_01997_, _01995_, _01985_);
  not (_01998_, _41971_);
  and (_01999_, _01747_, _01998_);
  not (_02001_, _42020_);
  and (_02002_, _01775_, _02001_);
  or (_02003_, _02002_, _01999_);
  or (_02005_, _02003_, _01997_);
  or (_02006_, _02005_, _01982_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02006_, _01971_);
  not (_02007_, _42517_);
  and (_02008_, _01706_, _02007_);
  not (_02009_, _42476_);
  and (_02010_, _01702_, _02009_);
  or (_02011_, _02010_, _02008_);
  not (_02012_, _42435_);
  and (_02013_, _01711_, _02012_);
  not (_02014_, _42107_);
  and (_02015_, _01731_, _02014_);
  not (_02016_, _41887_);
  and (_02017_, _01727_, _02016_);
  or (_02018_, _02017_, _02015_);
  not (_02019_, _42148_);
  and (_02020_, _01715_, _02019_);
  not (_02021_, _42189_);
  and (_02022_, _01719_, _02021_);
  or (_02023_, _02022_, _02020_);
  or (_02024_, _02023_, _02018_);
  or (_02026_, _02024_, _02013_);
  or (_02027_, _02026_, _02011_);
  not (_02029_, _42025_);
  and (_02030_, _01775_, _02029_);
  not (_02031_, _41928_);
  and (_02033_, _01743_, _02031_);
  not (_02034_, _42312_);
  and (_02035_, _01751_, _02034_);
  or (_02037_, _02035_, _02033_);
  or (_02038_, _02037_, _02030_);
  not (_02039_, _42271_);
  and (_02041_, _01756_, _02039_);
  not (_02042_, _42394_);
  and (_02043_, _01760_, _02042_);
  not (_02045_, _42066_);
  and (_02046_, _01763_, _02045_);
  not (_02047_, _42230_);
  and (_02049_, _01767_, _02047_);
  or (_02050_, _02049_, _02046_);
  or (_02051_, _02050_, _02043_);
  or (_02053_, _02051_, _02041_);
  not (_02054_, _41976_);
  and (_02055_, _01747_, _02054_);
  not (_02057_, _42353_);
  and (_02058_, _01779_, _02057_);
  or (_02059_, _02058_, _02055_);
  or (_02060_, _02059_, _02053_);
  or (_02061_, _02060_, _02038_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02061_, _02027_);
  not (_02062_, _42440_);
  and (_02063_, _01711_, _02062_);
  not (_02064_, _42481_);
  and (_02065_, _01702_, _02064_);
  or (_02066_, _02065_, _02063_);
  not (_02067_, _42522_);
  and (_02068_, _01706_, _02067_);
  not (_02069_, _42112_);
  and (_02070_, _01731_, _02069_);
  not (_02071_, _42153_);
  and (_02072_, _01715_, _02071_);
  or (_02073_, _02072_, _02070_);
  not (_02074_, _41892_);
  and (_02075_, _01727_, _02074_);
  not (_02076_, _42194_);
  and (_02078_, _01719_, _02076_);
  or (_02079_, _02078_, _02075_);
  or (_02081_, _02079_, _02073_);
  or (_02082_, _02081_, _02068_);
  or (_02083_, _02082_, _02066_);
  not (_02085_, _41986_);
  and (_02086_, _01747_, _02085_);
  not (_02087_, _41934_);
  and (_02089_, _01743_, _02087_);
  not (_02090_, _42030_);
  and (_02091_, _01775_, _02090_);
  or (_02093_, _02091_, _02089_);
  or (_02094_, _02093_, _02086_);
  not (_02095_, _42317_);
  and (_02097_, _01751_, _02095_);
  not (_02098_, _42071_);
  and (_02099_, _01763_, _02098_);
  not (_02101_, _42235_);
  and (_02102_, _01767_, _02101_);
  not (_02103_, _42399_);
  and (_02105_, _01760_, _02103_);
  or (_02106_, _02105_, _02102_);
  or (_02107_, _02106_, _02099_);
  or (_02109_, _02107_, _02097_);
  not (_02110_, _42276_);
  and (_02111_, _01756_, _02110_);
  not (_02112_, _42358_);
  and (_02113_, _01779_, _02112_);
  or (_02114_, _02113_, _02111_);
  or (_02115_, _02114_, _02109_);
  or (_02116_, _02115_, _02094_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02116_, _02083_);
  not (_02117_, _42445_);
  and (_02118_, _01711_, _02117_);
  not (_02119_, _42486_);
  and (_02120_, _01702_, _02119_);
  or (_02121_, _02120_, _02118_);
  not (_02122_, _42527_);
  and (_02123_, _01706_, _02122_);
  not (_02124_, _42199_);
  and (_02125_, _01719_, _02124_);
  not (_02126_, _42158_);
  and (_02127_, _01715_, _02126_);
  or (_02128_, _02127_, _02125_);
  not (_02130_, _42117_);
  and (_02131_, _01731_, _02130_);
  not (_02133_, _41897_);
  and (_02134_, _01727_, _02133_);
  or (_02135_, _02134_, _02131_);
  or (_02137_, _02135_, _02128_);
  or (_02138_, _02137_, _02123_);
  or (_02139_, _02138_, _02121_);
  not (_02141_, _42363_);
  and (_02142_, _01779_, _02141_);
  not (_02143_, _42281_);
  and (_02145_, _01756_, _02143_);
  not (_02146_, _41994_);
  and (_02147_, _01747_, _02146_);
  or (_02149_, _02147_, _02145_);
  or (_02150_, _02149_, _02142_);
  not (_02151_, _41943_);
  and (_02153_, _01743_, _02151_);
  not (_02154_, _42076_);
  and (_02155_, _01763_, _02154_);
  not (_02157_, _42404_);
  and (_02158_, _01760_, _02157_);
  not (_02159_, _42240_);
  and (_02161_, _01767_, _02159_);
  or (_02162_, _02161_, _02158_);
  or (_02163_, _02162_, _02155_);
  or (_02164_, _02163_, _02153_);
  not (_02165_, _42322_);
  and (_02166_, _01751_, _02165_);
  not (_02167_, _42035_);
  and (_02168_, _01775_, _02167_);
  or (_02169_, _02168_, _02166_);
  or (_02170_, _02169_, _02164_);
  or (_02171_, _02170_, _02150_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02171_, _02139_);
  not (_02172_, _42450_);
  and (_02173_, _01711_, _02172_);
  not (_02174_, _42491_);
  and (_02175_, _01702_, _02174_);
  or (_02176_, _02175_, _02173_);
  not (_02177_, _42532_);
  and (_02178_, _01706_, _02177_);
  not (_02179_, _42204_);
  and (_02180_, _01719_, _02179_);
  not (_02182_, _42163_);
  and (_02183_, _01715_, _02182_);
  or (_02185_, _02183_, _02180_);
  not (_02186_, _42122_);
  and (_02187_, _01731_, _02186_);
  not (_02189_, _41902_);
  and (_02190_, _01727_, _02189_);
  or (_02191_, _02190_, _02187_);
  or (_02193_, _02191_, _02185_);
  or (_02194_, _02193_, _02178_);
  or (_02195_, _02194_, _02176_);
  not (_02197_, _42368_);
  and (_02198_, _01779_, _02197_);
  not (_02199_, _42286_);
  and (_02201_, _01756_, _02199_);
  not (_02202_, _41999_);
  and (_02203_, _01747_, _02202_);
  or (_02205_, _02203_, _02201_);
  or (_02206_, _02205_, _02198_);
  not (_02207_, _41950_);
  and (_02209_, _01743_, _02207_);
  not (_02210_, _42081_);
  and (_02211_, _01763_, _02210_);
  not (_02213_, _42409_);
  and (_02214_, _01760_, _02213_);
  not (_02215_, _42245_);
  and (_02216_, _01767_, _02215_);
  or (_02217_, _02216_, _02214_);
  or (_02218_, _02217_, _02211_);
  or (_02219_, _02218_, _02209_);
  not (_02220_, _42327_);
  and (_02221_, _01751_, _02220_);
  not (_02222_, _42040_);
  and (_02223_, _01775_, _02222_);
  or (_02224_, _02223_, _02221_);
  or (_02225_, _02224_, _02219_);
  or (_02226_, _02225_, _02206_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02226_, _02195_);
  not (_02227_, _42455_);
  and (_02228_, _01711_, _02227_);
  not (_02229_, _42496_);
  and (_02230_, _01702_, _02229_);
  or (_02231_, _02230_, _02228_);
  not (_02232_, _42537_);
  and (_02233_, _01706_, _02232_);
  not (_02234_, _42209_);
  and (_02235_, _01719_, _02234_);
  not (_02236_, _42127_);
  and (_02237_, _01731_, _02236_);
  or (_02238_, _02237_, _02235_);
  not (_02239_, _42168_);
  and (_02240_, _01715_, _02239_);
  not (_02241_, _41907_);
  and (_02242_, _01727_, _02241_);
  or (_02243_, _02242_, _02240_);
  or (_02244_, _02243_, _02238_);
  or (_02245_, _02244_, _02233_);
  or (_02246_, _02245_, _02231_);
  not (_02247_, _42373_);
  and (_02248_, _01779_, _02247_);
  not (_02249_, _42291_);
  and (_02250_, _01756_, _02249_);
  not (_02251_, _42004_);
  and (_02252_, _01747_, _02251_);
  or (_02253_, _02252_, _02250_);
  or (_02254_, _02253_, _02248_);
  not (_02255_, _41955_);
  and (_02256_, _01743_, _02255_);
  not (_02257_, _42086_);
  and (_02258_, _01763_, _02257_);
  not (_02259_, _42414_);
  and (_02260_, _01760_, _02259_);
  not (_02261_, _42250_);
  and (_02262_, _01767_, _02261_);
  or (_02263_, _02262_, _02260_);
  or (_02264_, _02263_, _02258_);
  or (_02265_, _02264_, _02256_);
  not (_02266_, _42332_);
  and (_02267_, _01751_, _02266_);
  not (_02268_, _42045_);
  and (_02269_, _01775_, _02268_);
  or (_02270_, _02269_, _02267_);
  or (_02271_, _02270_, _02265_);
  or (_02272_, _02271_, _02254_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02272_, _02246_);
  and (_02273_, _01702_, _01927_);
  and (_02274_, _01706_, _01922_);
  or (_02275_, _02274_, _02273_);
  and (_02276_, _01711_, _01911_);
  and (_02277_, _01715_, _01919_);
  and (_02278_, _01731_, _01935_);
  or (_02279_, _02278_, _02277_);
  and (_02280_, _01719_, _01942_);
  and (_02281_, _01727_, _01945_);
  or (_02282_, _02281_, _02280_);
  or (_02283_, _02282_, _02279_);
  or (_02284_, _02283_, _02276_);
  or (_02285_, _02284_, _02275_);
  and (_02286_, _01775_, _01906_);
  and (_02287_, _01751_, _01896_);
  and (_02288_, _01756_, _01933_);
  or (_02289_, _02288_, _02287_);
  or (_02290_, _02289_, _02286_);
  and (_02291_, _01747_, _01909_);
  and (_02292_, _01760_, _01902_);
  and (_02293_, _01767_, _01917_);
  and (_02294_, _01763_, _01904_);
  or (_02295_, _02294_, _02293_);
  or (_02296_, _02295_, _02292_);
  or (_02297_, _02296_, _02291_);
  and (_02298_, _01779_, _01898_);
  and (_02299_, _01743_, _01930_);
  or (_02300_, _02299_, _02298_);
  or (_02301_, _02300_, _02297_);
  or (_02302_, _02301_, _02290_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _02302_, _02285_);
  and (_02303_, _01711_, _01964_);
  and (_02304_, _01706_, _01998_);
  or (_02305_, _02304_, _02303_);
  and (_02306_, _01702_, _01975_);
  and (_02307_, _01715_, _01972_);
  and (_02308_, _01731_, _01991_);
  or (_02309_, _02308_, _02307_);
  and (_02310_, _01719_, _01983_);
  and (_02311_, _01727_, _02001_);
  or (_02312_, _02311_, _02310_);
  or (_02313_, _02312_, _02309_);
  or (_02314_, _02313_, _02306_);
  or (_02315_, _02314_, _02305_);
  and (_02316_, _01751_, _01952_);
  and (_02317_, _01747_, _01959_);
  and (_02318_, _01743_, _01989_);
  or (_02319_, _02318_, _02317_);
  or (_02320_, _02319_, _02316_);
  and (_02321_, _01775_, _01961_);
  and (_02322_, _01767_, _01978_);
  and (_02323_, _01760_, _01957_);
  and (_02324_, _01763_, _01966_);
  or (_02325_, _02324_, _02323_);
  or (_02326_, _02325_, _02322_);
  or (_02327_, _02326_, _02321_);
  and (_02328_, _01779_, _01954_);
  and (_02329_, _01756_, _01986_);
  or (_02330_, _02329_, _02328_);
  or (_02331_, _02330_, _02327_);
  or (_02332_, _02331_, _02320_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _02332_, _02315_);
  and (_02333_, _01706_, _02054_);
  and (_02334_, _01702_, _02031_);
  or (_02335_, _02334_, _02333_);
  and (_02336_, _01711_, _02016_);
  and (_02337_, _01715_, _02039_);
  and (_02338_, _01719_, _02034_);
  or (_02339_, _02338_, _02337_);
  and (_02340_, _01727_, _02029_);
  and (_02341_, _01731_, _02047_);
  or (_02342_, _02341_, _02340_);
  or (_02343_, _02342_, _02339_);
  or (_02344_, _02343_, _02336_);
  or (_02345_, _02344_, _02335_);
  and (_02346_, _01747_, _02014_);
  and (_02347_, _01775_, _02019_);
  or (_02348_, _02347_, _02346_);
  and (_02349_, _01751_, _02012_);
  or (_02350_, _02349_, _02348_);
  and (_02351_, _01756_, _02042_);
  and (_02352_, _01760_, _02007_);
  and (_02353_, _01763_, _02021_);
  and (_02354_, _01767_, _02057_);
  or (_02355_, _02354_, _02353_);
  or (_02356_, _02355_, _02352_);
  or (_02357_, _02356_, _02351_);
  and (_02358_, _01743_, _02045_);
  and (_02359_, _01779_, _02009_);
  or (_02360_, _02359_, _02358_);
  or (_02361_, _02360_, _02357_);
  or (_02362_, _02361_, _02350_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _02362_, _02345_);
  and (_02363_, _01711_, _02074_);
  and (_02364_, _01706_, _02085_);
  or (_02365_, _02364_, _02363_);
  and (_02366_, _01702_, _02087_);
  and (_02367_, _01727_, _02090_);
  and (_02368_, _01715_, _02110_);
  or (_02369_, _02368_, _02367_);
  and (_02370_, _01719_, _02095_);
  and (_02371_, _01731_, _02101_);
  or (_02372_, _02371_, _02370_);
  or (_02373_, _02372_, _02369_);
  or (_02374_, _02373_, _02366_);
  or (_02375_, _02374_, _02365_);
  and (_02376_, _01747_, _02069_);
  and (_02377_, _01775_, _02071_);
  or (_02378_, _02377_, _02376_);
  and (_02379_, _01779_, _02064_);
  or (_02380_, _02379_, _02378_);
  and (_02381_, _01756_, _02103_);
  and (_02382_, _01760_, _02067_);
  and (_02383_, _01763_, _02076_);
  and (_02384_, _01767_, _02112_);
  or (_02385_, _02384_, _02383_);
  or (_02386_, _02385_, _02382_);
  or (_02387_, _02386_, _02381_);
  and (_02388_, _01743_, _02098_);
  and (_02389_, _01751_, _02062_);
  or (_02390_, _02389_, _02388_);
  or (_02391_, _02390_, _02387_);
  or (_02392_, _02391_, _02380_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _02392_, _02375_);
  and (_02393_, _01702_, _02151_);
  and (_02394_, _01706_, _02146_);
  or (_02395_, _02394_, _02393_);
  and (_02396_, _01711_, _02133_);
  and (_02397_, _01719_, _02165_);
  and (_02398_, _01727_, _02167_);
  or (_02399_, _02398_, _02397_);
  and (_02400_, _01715_, _02143_);
  and (_02401_, _01731_, _02159_);
  or (_02402_, _02401_, _02400_);
  or (_02403_, _02402_, _02399_);
  or (_02404_, _02403_, _02396_);
  or (_02405_, _02404_, _02395_);
  and (_02406_, _01775_, _02126_);
  and (_02407_, _01756_, _02157_);
  and (_02408_, _01747_, _02130_);
  or (_02409_, _02408_, _02407_);
  or (_02410_, _02409_, _02406_);
  and (_02411_, _01751_, _02117_);
  and (_02412_, _01779_, _02119_);
  or (_02413_, _02412_, _02411_);
  and (_02414_, _01743_, _02154_);
  and (_02415_, _01760_, _02122_);
  and (_02416_, _01767_, _02141_);
  and (_02417_, _01763_, _02124_);
  or (_02418_, _02417_, _02416_);
  or (_02419_, _02418_, _02415_);
  or (_02420_, _02419_, _02414_);
  or (_02421_, _02420_, _02413_);
  or (_02422_, _02421_, _02410_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _02422_, _02405_);
  and (_02423_, _01706_, _02202_);
  and (_02424_, _01702_, _02207_);
  or (_02425_, _02424_, _02423_);
  and (_02426_, _01711_, _02189_);
  and (_02427_, _01719_, _02220_);
  and (_02428_, _01715_, _02199_);
  or (_02429_, _02428_, _02427_);
  and (_02430_, _01727_, _02222_);
  and (_02431_, _01731_, _02215_);
  or (_02432_, _02431_, _02430_);
  or (_02433_, _02432_, _02429_);
  or (_02434_, _02433_, _02426_);
  or (_02435_, _02434_, _02425_);
  and (_02436_, _01779_, _02174_);
  and (_02437_, _01743_, _02210_);
  and (_02438_, _01756_, _02213_);
  or (_02439_, _02438_, _02437_);
  or (_02440_, _02439_, _02436_);
  and (_02441_, _01775_, _02182_);
  and (_02442_, _01767_, _02197_);
  and (_02443_, _01760_, _02177_);
  and (_02444_, _01763_, _02179_);
  or (_02445_, _02444_, _02443_);
  or (_02446_, _02445_, _02442_);
  or (_02447_, _02446_, _02441_);
  and (_02448_, _01747_, _02186_);
  and (_02449_, _01751_, _02172_);
  or (_02450_, _02449_, _02448_);
  or (_02451_, _02450_, _02447_);
  or (_02452_, _02451_, _02440_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _02452_, _02435_);
  and (_02453_, _01711_, _02241_);
  and (_02455_, _01706_, _02251_);
  or (_02456_, _02455_, _02453_);
  and (_02457_, _01702_, _02255_);
  and (_02458_, _01727_, _02268_);
  and (_02459_, _01715_, _02249_);
  or (_02460_, _02459_, _02458_);
  and (_02461_, _01719_, _02266_);
  and (_02462_, _01731_, _02261_);
  or (_02463_, _02462_, _02461_);
  or (_02464_, _02463_, _02460_);
  or (_02465_, _02464_, _02457_);
  or (_02466_, _02465_, _02456_);
  and (_02467_, _01751_, _02227_);
  and (_02468_, _01747_, _02236_);
  and (_02469_, _01779_, _02229_);
  or (_02470_, _02469_, _02468_);
  or (_02471_, _02470_, _02467_);
  and (_02472_, _01756_, _02259_);
  and (_02473_, _01763_, _02234_);
  and (_02474_, _01760_, _02232_);
  and (_02475_, _01767_, _02247_);
  or (_02476_, _02475_, _02474_);
  or (_02477_, _02476_, _02473_);
  or (_02478_, _02477_, _02472_);
  and (_02479_, _01775_, _02239_);
  and (_02480_, _01743_, _02257_);
  or (_02481_, _02480_, _02479_);
  or (_02482_, _02481_, _02478_);
  or (_02483_, _02482_, _02471_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _02483_, _02466_);
  and (_02484_, _01706_, _01927_);
  and (_02485_, _01719_, _01919_);
  and (_02486_, _01731_, _01904_);
  or (_02487_, _02486_, _02485_);
  and (_02488_, _01715_, _01935_);
  and (_02489_, _01727_, _01922_);
  or (_02490_, _02489_, _02488_);
  or (_02491_, _02490_, _02487_);
  or (_02492_, _02491_, _02484_);
  and (_02493_, _01711_, _01902_);
  and (_02494_, _01702_, _01911_);
  or (_02495_, _02494_, _02493_);
  or (_02496_, _02495_, _02492_);
  and (_02497_, _01775_, _01909_);
  and (_02498_, _01756_, _01917_);
  and (_02499_, _01747_, _01930_);
  or (_02500_, _02499_, _02498_);
  or (_02501_, _02500_, _02497_);
  and (_02502_, _01779_, _01896_);
  and (_02503_, _01763_, _01906_);
  and (_02504_, _01760_, _01898_);
  and (_02505_, _01767_, _01942_);
  or (_02506_, _02505_, _02504_);
  or (_02507_, _02506_, _02503_);
  or (_02508_, _02507_, _02502_);
  and (_02509_, _01751_, _01933_);
  and (_02510_, _01743_, _01945_);
  or (_02511_, _02510_, _02509_);
  or (_02512_, _02511_, _02508_);
  or (_02513_, _02512_, _02501_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _02513_, _02496_);
  and (_02514_, _01706_, _01975_);
  and (_02515_, _01715_, _01991_);
  and (_02516_, _01727_, _01998_);
  or (_02517_, _02516_, _02515_);
  and (_02518_, _01719_, _01972_);
  and (_02519_, _01731_, _01966_);
  or (_02520_, _02519_, _02518_);
  or (_02521_, _02520_, _02517_);
  or (_02522_, _02521_, _02514_);
  and (_02523_, _01711_, _01957_);
  and (_02524_, _01702_, _01964_);
  or (_02525_, _02524_, _02523_);
  or (_02526_, _02525_, _02522_);
  and (_02527_, _01779_, _01952_);
  and (_02528_, _01751_, _01986_);
  and (_02529_, _01747_, _01989_);
  or (_02530_, _02529_, _02528_);
  or (_02531_, _02530_, _02527_);
  and (_02532_, _01743_, _02001_);
  and (_02533_, _01767_, _01983_);
  and (_02534_, _01760_, _01954_);
  and (_02535_, _01763_, _01961_);
  or (_02536_, _02535_, _02534_);
  or (_02537_, _02536_, _02533_);
  or (_02538_, _02537_, _02532_);
  and (_02539_, _01756_, _01978_);
  and (_02540_, _01775_, _01959_);
  or (_02541_, _02540_, _02539_);
  or (_02542_, _02541_, _02538_);
  or (_02543_, _02542_, _02531_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02543_, _02526_);
  and (_02544_, _01706_, _02031_);
  and (_02545_, _01727_, _02054_);
  and (_02546_, _01731_, _02021_);
  or (_02547_, _02546_, _02545_);
  and (_02548_, _01719_, _02039_);
  and (_02549_, _01715_, _02047_);
  or (_02550_, _02549_, _02548_);
  or (_02551_, _02550_, _02547_);
  or (_02552_, _02551_, _02544_);
  and (_02553_, _01711_, _02007_);
  and (_02554_, _01702_, _02016_);
  or (_02555_, _02554_, _02553_);
  or (_02556_, _02555_, _02552_);
  and (_02557_, _01747_, _02045_);
  and (_02558_, _01775_, _02014_);
  and (_02559_, _01756_, _02057_);
  or (_02560_, _02559_, _02558_);
  or (_02561_, _02560_, _02557_);
  and (_02562_, _01751_, _02042_);
  and (_02563_, _01767_, _02034_);
  and (_02564_, _01763_, _02019_);
  and (_02565_, _01760_, _02009_);
  or (_02566_, _02565_, _02564_);
  or (_02567_, _02566_, _02563_);
  or (_02568_, _02567_, _02562_);
  and (_02569_, _01743_, _02029_);
  and (_02570_, _01779_, _02012_);
  or (_02571_, _02570_, _02569_);
  or (_02572_, _02571_, _02568_);
  or (_02573_, _02572_, _02561_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02573_, _02556_);
  and (_02574_, _01702_, _02074_);
  and (_02575_, _01715_, _02101_);
  and (_02576_, _01731_, _02076_);
  or (_02577_, _02576_, _02575_);
  and (_02578_, _01727_, _02085_);
  and (_02579_, _01719_, _02110_);
  or (_02580_, _02579_, _02578_);
  or (_02581_, _02580_, _02577_);
  or (_02582_, _02581_, _02574_);
  and (_02583_, _01711_, _02067_);
  and (_02584_, _01706_, _02087_);
  or (_02585_, _02584_, _02583_);
  or (_02586_, _02585_, _02582_);
  and (_02587_, _01743_, _02090_);
  and (_02588_, _01747_, _02098_);
  and (_02589_, _01756_, _02112_);
  or (_02590_, _02589_, _02588_);
  or (_02591_, _02590_, _02587_);
  and (_02592_, _01751_, _02103_);
  and (_02593_, _01767_, _02095_);
  and (_02594_, _01763_, _02071_);
  and (_02595_, _01760_, _02064_);
  or (_02596_, _02595_, _02594_);
  or (_02597_, _02596_, _02593_);
  or (_02598_, _02597_, _02592_);
  and (_02599_, _01775_, _02069_);
  and (_02600_, _01779_, _02062_);
  or (_02601_, _02600_, _02599_);
  or (_02602_, _02601_, _02598_);
  or (_02603_, _02602_, _02591_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02603_, _02586_);
  and (_02604_, _01711_, _02122_);
  and (_02605_, _01727_, _02146_);
  and (_02606_, _01731_, _02124_);
  or (_02607_, _02606_, _02605_);
  and (_02608_, _01719_, _02143_);
  and (_02609_, _01715_, _02159_);
  or (_02610_, _02609_, _02608_);
  or (_02611_, _02610_, _02607_);
  or (_02612_, _02611_, _02604_);
  and (_02613_, _01702_, _02133_);
  and (_02614_, _01706_, _02151_);
  or (_02615_, _02614_, _02613_);
  or (_02616_, _02615_, _02612_);
  and (_02617_, _01779_, _02117_);
  and (_02618_, _01775_, _02130_);
  and (_02619_, _01747_, _02154_);
  or (_02620_, _02619_, _02618_);
  or (_02621_, _02620_, _02617_);
  and (_02622_, _01756_, _02141_);
  and (_02623_, _01760_, _02119_);
  and (_02624_, _01763_, _02126_);
  and (_02625_, _01767_, _02165_);
  or (_02626_, _02625_, _02624_);
  or (_02627_, _02626_, _02623_);
  or (_02628_, _02627_, _02622_);
  and (_02629_, _01743_, _02167_);
  and (_02630_, _01751_, _02157_);
  or (_02631_, _02630_, _02629_);
  or (_02632_, _02631_, _02628_);
  or (_02633_, _02632_, _02621_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _02633_, _02616_);
  and (_02634_, _01702_, _02189_);
  and (_02635_, _01719_, _02199_);
  and (_02636_, _01715_, _02215_);
  or (_02637_, _02636_, _02635_);
  and (_02638_, _01731_, _02179_);
  and (_02639_, _01727_, _02202_);
  or (_02640_, _02639_, _02638_);
  or (_02641_, _02640_, _02637_);
  or (_02642_, _02641_, _02634_);
  and (_02643_, _01711_, _02177_);
  and (_02644_, _01706_, _02207_);
  or (_02645_, _02644_, _02643_);
  or (_02646_, _02645_, _02642_);
  and (_02647_, _01779_, _02172_);
  and (_02648_, _01775_, _02186_);
  and (_02650_, _01743_, _02222_);
  or (_02651_, _02650_, _02648_);
  or (_02652_, _02651_, _02647_);
  and (_02653_, _01756_, _02197_);
  and (_02654_, _01751_, _02213_);
  or (_02655_, _02654_, _02653_);
  and (_02656_, _01747_, _02210_);
  and (_02657_, _01760_, _02174_);
  and (_02658_, _01767_, _02220_);
  and (_02659_, _01763_, _02182_);
  or (_02660_, _02659_, _02658_);
  or (_02661_, _02660_, _02657_);
  or (_02662_, _02661_, _02656_);
  or (_02663_, _02662_, _02655_);
  or (_02664_, _02663_, _02652_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _02664_, _02646_);
  and (_02665_, _01706_, _02255_);
  and (_02666_, _01715_, _02261_);
  and (_02667_, _01727_, _02251_);
  or (_02668_, _02667_, _02666_);
  and (_02669_, _01719_, _02249_);
  and (_02670_, _01731_, _02234_);
  or (_02671_, _02670_, _02669_);
  or (_02672_, _02671_, _02668_);
  or (_02673_, _02672_, _02665_);
  and (_02674_, _01711_, _02232_);
  and (_02675_, _01702_, _02241_);
  or (_02676_, _02675_, _02674_);
  or (_02677_, _02676_, _02673_);
  and (_02678_, _01779_, _02227_);
  and (_02679_, _01751_, _02259_);
  and (_02680_, _01747_, _02257_);
  or (_02681_, _02680_, _02679_);
  or (_02682_, _02681_, _02678_);
  and (_02683_, _01743_, _02268_);
  and (_02684_, _01767_, _02266_);
  and (_02685_, _01760_, _02229_);
  and (_02686_, _01763_, _02239_);
  or (_02687_, _02686_, _02685_);
  or (_02688_, _02687_, _02684_);
  or (_02689_, _02688_, _02683_);
  and (_02690_, _01756_, _02247_);
  and (_02691_, _01775_, _02236_);
  or (_02692_, _02691_, _02690_);
  or (_02693_, _02692_, _02689_);
  or (_02694_, _02693_, _02682_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02694_, _02677_);
  and (_02695_, _01702_, _01902_);
  and (_02696_, _01727_, _01927_);
  and (_02697_, _01719_, _01935_);
  or (_02698_, _02697_, _02696_);
  and (_02699_, _01731_, _01906_);
  and (_02700_, _01715_, _01904_);
  or (_02701_, _02700_, _02699_);
  or (_02702_, _02701_, _02698_);
  or (_02703_, _02702_, _02695_);
  and (_02704_, _01706_, _01911_);
  and (_02705_, _01711_, _01898_);
  or (_02706_, _02705_, _02704_);
  or (_02707_, _02706_, _02703_);
  and (_02708_, _01756_, _01942_);
  and (_02709_, _01743_, _01922_);
  and (_02710_, _01751_, _01917_);
  or (_02711_, _02710_, _02709_);
  or (_02712_, _02711_, _02708_);
  and (_02713_, _01747_, _01945_);
  and (_02714_, _01760_, _01896_);
  and (_02715_, _01763_, _01909_);
  and (_02716_, _01767_, _01919_);
  or (_02717_, _02716_, _02715_);
  or (_02718_, _02717_, _02714_);
  or (_02719_, _02718_, _02713_);
  and (_02720_, _01775_, _01930_);
  and (_02721_, _01779_, _01933_);
  or (_02722_, _02721_, _02720_);
  or (_02723_, _02722_, _02719_);
  or (_02724_, _02723_, _02712_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _02724_, _02707_);
  and (_02725_, _01702_, _01957_);
  and (_02726_, _01719_, _01991_);
  and (_02727_, _01715_, _01966_);
  or (_02728_, _02727_, _02726_);
  and (_02729_, _01727_, _01975_);
  and (_02730_, _01731_, _01961_);
  or (_02731_, _02730_, _02729_);
  or (_02732_, _02731_, _02728_);
  or (_02733_, _02732_, _02725_);
  and (_02734_, _01711_, _01954_);
  and (_02735_, _01706_, _01964_);
  or (_02736_, _02735_, _02734_);
  or (_02737_, _02736_, _02733_);
  and (_02738_, _01779_, _01986_);
  and (_02739_, _01756_, _01983_);
  and (_02740_, _01743_, _01998_);
  or (_02741_, _02740_, _02739_);
  or (_02742_, _02741_, _02738_);
  and (_02743_, _01775_, _01989_);
  and (_02744_, _01747_, _02001_);
  or (_02745_, _02744_, _02743_);
  and (_02746_, _01751_, _01978_);
  and (_02747_, _01767_, _01972_);
  and (_02748_, _01760_, _01952_);
  and (_02749_, _01763_, _01959_);
  or (_02750_, _02749_, _02748_);
  or (_02751_, _02750_, _02747_);
  or (_02752_, _02751_, _02746_);
  or (_02753_, _02752_, _02745_);
  or (_02754_, _02753_, _02742_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _02754_, _02737_);
  and (_02755_, _01702_, _02007_);
  and (_02756_, _01711_, _02009_);
  or (_02757_, _02756_, _02755_);
  and (_02758_, _01751_, _02057_);
  and (_02759_, _01756_, _02034_);
  and (_02760_, _01715_, _02021_);
  and (_02761_, _01719_, _02047_);
  or (_02762_, _02761_, _02760_);
  and (_02763_, _01767_, _02039_);
  or (_02764_, _02763_, _02762_);
  or (_02765_, _02764_, _02759_);
  or (_02766_, _02765_, _02758_);
  or (_02767_, _02766_, _02757_);
  and (_02768_, _01706_, _02016_);
  and (_02769_, _01727_, _02031_);
  and (_02770_, _01743_, _02054_);
  or (_02771_, _02770_, _02769_);
  or (_02772_, _02771_, _02768_);
  and (_02773_, _01747_, _02029_);
  and (_02774_, _01775_, _02045_);
  or (_02775_, _02774_, _02773_);
  and (_02776_, _01731_, _02019_);
  and (_02777_, _01763_, _02014_);
  or (_02778_, _02777_, _02776_);
  or (_02779_, _02778_, _02775_);
  or (_02780_, _02779_, _02772_);
  and (_02781_, _01779_, _02042_);
  and (_02782_, _01760_, _02012_);
  or (_02783_, _02782_, _02781_);
  or (_02784_, _02783_, _02780_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _02784_, _02767_);
  and (_02785_, _01702_, _02067_);
  and (_02786_, _01711_, _02064_);
  or (_02787_, _02786_, _02785_);
  and (_02788_, _01706_, _02074_);
  and (_02789_, _01727_, _02087_);
  and (_02790_, _01715_, _02076_);
  or (_02791_, _02790_, _02789_);
  and (_02792_, _01731_, _02071_);
  and (_02793_, _01719_, _02101_);
  or (_02794_, _02793_, _02792_);
  or (_02795_, _02794_, _02791_);
  or (_02796_, _02795_, _02788_);
  or (_02797_, _02796_, _02787_);
  and (_02798_, _01743_, _02085_);
  and (_02799_, _01747_, _02090_);
  and (_02800_, _01779_, _02103_);
  or (_02801_, _02800_, _02799_);
  or (_02802_, _02801_, _02798_);
  and (_02803_, _01751_, _02112_);
  and (_02804_, _01767_, _02110_);
  and (_02805_, _01763_, _02069_);
  and (_02806_, _01760_, _02062_);
  or (_02807_, _02806_, _02805_);
  or (_02808_, _02807_, _02804_);
  or (_02809_, _02808_, _02803_);
  and (_02810_, _01775_, _02098_);
  and (_02811_, _01756_, _02095_);
  or (_02812_, _02811_, _02810_);
  or (_02813_, _02812_, _02809_);
  or (_02814_, _02813_, _02802_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _02814_, _02797_);
  and (_02815_, _01702_, _02122_);
  and (_02816_, _01719_, _02159_);
  and (_02817_, _01715_, _02124_);
  or (_02818_, _02817_, _02816_);
  and (_02819_, _01731_, _02126_);
  and (_02820_, _01727_, _02151_);
  or (_02821_, _02820_, _02819_);
  or (_02822_, _02821_, _02818_);
  or (_02823_, _02822_, _02815_);
  and (_02824_, _01711_, _02119_);
  and (_02825_, _01706_, _02133_);
  or (_02826_, _02825_, _02824_);
  or (_02827_, _02826_, _02823_);
  and (_02828_, _01751_, _02141_);
  and (_02829_, _01756_, _02165_);
  and (_02830_, _01743_, _02146_);
  or (_02831_, _02830_, _02829_);
  or (_02832_, _02831_, _02828_);
  and (_02833_, _01775_, _02154_);
  and (_02834_, _01747_, _02167_);
  or (_02835_, _02834_, _02833_);
  and (_02836_, _01779_, _02157_);
  and (_02837_, _01767_, _02143_);
  and (_02838_, _01760_, _02117_);
  and (_02839_, _01763_, _02130_);
  or (_02840_, _02839_, _02838_);
  or (_02841_, _02840_, _02837_);
  or (_02842_, _02841_, _02836_);
  or (_02843_, _02842_, _02835_);
  or (_02845_, _02843_, _02832_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _02845_, _02827_);
  and (_02846_, _01702_, _02177_);
  and (_02847_, _01711_, _02174_);
  or (_02848_, _02847_, _02846_);
  and (_02849_, _01779_, _02213_);
  and (_02850_, _01756_, _02220_);
  and (_02851_, _01715_, _02179_);
  and (_02852_, _01719_, _02215_);
  or (_02853_, _02852_, _02851_);
  and (_02854_, _01767_, _02199_);
  or (_02855_, _02854_, _02853_);
  or (_02856_, _02855_, _02850_);
  or (_02857_, _02856_, _02849_);
  or (_02858_, _02857_, _02848_);
  and (_02859_, _01706_, _02189_);
  and (_02860_, _01727_, _02207_);
  and (_02861_, _01743_, _02202_);
  or (_02862_, _02861_, _02860_);
  or (_02863_, _02862_, _02859_);
  and (_02864_, _01747_, _02222_);
  and (_02865_, _01775_, _02210_);
  or (_02866_, _02865_, _02864_);
  and (_02867_, _01731_, _02182_);
  and (_02868_, _01763_, _02186_);
  or (_02869_, _02868_, _02867_);
  or (_02870_, _02869_, _02866_);
  or (_02871_, _02870_, _02863_);
  and (_02872_, _01751_, _02197_);
  and (_02873_, _01760_, _02172_);
  or (_02874_, _02873_, _02872_);
  or (_02875_, _02874_, _02871_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _02875_, _02858_);
  and (_02876_, _01702_, _02232_);
  and (_02877_, _01719_, _02261_);
  and (_02878_, _01715_, _02234_);
  or (_02879_, _02878_, _02877_);
  and (_02880_, _01727_, _02255_);
  and (_02881_, _01731_, _02239_);
  or (_02882_, _02881_, _02880_);
  or (_02883_, _02882_, _02879_);
  or (_02884_, _02883_, _02876_);
  and (_02885_, _01711_, _02229_);
  and (_02886_, _01706_, _02241_);
  or (_02887_, _02886_, _02885_);
  or (_02888_, _02887_, _02884_);
  and (_02889_, _01751_, _02247_);
  and (_02890_, _01756_, _02266_);
  and (_02891_, _01743_, _02251_);
  or (_02892_, _02891_, _02890_);
  or (_02893_, _02892_, _02889_);
  and (_02894_, _01775_, _02257_);
  and (_02895_, _01747_, _02268_);
  or (_02896_, _02895_, _02894_);
  and (_02897_, _01779_, _02259_);
  and (_02898_, _01767_, _02249_);
  and (_02899_, _01760_, _02227_);
  and (_02900_, _01763_, _02236_);
  or (_02901_, _02900_, _02899_);
  or (_02902_, _02901_, _02898_);
  or (_02903_, _02902_, _02897_);
  or (_02904_, _02903_, _02896_);
  or (_02905_, _02904_, _02893_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _02905_, _02888_);
  nand (_02906_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02907_, \oc8051_golden_model_1.PC [3]);
  or (_02908_, \oc8051_golden_model_1.PC [2], _02907_);
  or (_02909_, _02908_, _02906_);
  or (_02910_, _02909_, _42373_);
  not (_02911_, \oc8051_golden_model_1.PC [1]);
  or (_02912_, _02911_, \oc8051_golden_model_1.PC [0]);
  or (_02913_, _02912_, _02908_);
  or (_02914_, _02913_, _42332_);
  and (_02915_, _02914_, _02910_);
  not (_02916_, \oc8051_golden_model_1.PC [2]);
  or (_02917_, _02916_, \oc8051_golden_model_1.PC [3]);
  or (_02918_, _02917_, _02906_);
  or (_02919_, _02918_, _42209_);
  or (_02920_, _02917_, _02912_);
  or (_02921_, _02920_, _42168_);
  and (_02922_, _02921_, _02919_);
  and (_02923_, _02922_, _02915_);
  nand (_02924_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02925_, _02924_, _02906_);
  or (_02926_, _02925_, _42537_);
  or (_02927_, _02924_, _02912_);
  or (_02928_, _02927_, _42496_);
  and (_02929_, _02928_, _02926_);
  or (_02930_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02931_, _02930_, _02906_);
  or (_02932_, _02931_, _42045_);
  or (_02933_, _02930_, _02912_);
  or (_02934_, _02933_, _42004_);
  and (_02935_, _02934_, _02932_);
  and (_02936_, _02935_, _02929_);
  and (_02937_, _02936_, _02923_);
  not (_02938_, \oc8051_golden_model_1.PC [0]);
  or (_02939_, \oc8051_golden_model_1.PC [1], _02938_);
  or (_02940_, _02939_, _02924_);
  or (_02941_, _02940_, _42455_);
  or (_02942_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02943_, _02942_, _02924_);
  or (_02944_, _02943_, _42414_);
  and (_02945_, _02944_, _02941_);
  or (_02946_, _02930_, _02942_);
  or (_02947_, _02946_, _41907_);
  or (_02948_, _02930_, _02939_);
  or (_02949_, _02948_, _41955_);
  and (_02950_, _02949_, _02947_);
  and (_02951_, _02950_, _02945_);
  or (_02952_, _02939_, _02908_);
  or (_02953_, _02952_, _42291_);
  or (_02954_, _02942_, _02908_);
  or (_02955_, _02954_, _42250_);
  and (_02956_, _02955_, _02953_);
  or (_02957_, _02939_, _02917_);
  or (_02958_, _02957_, _42127_);
  or (_02959_, _02942_, _02917_);
  or (_02960_, _02959_, _42086_);
  and (_02961_, _02960_, _02958_);
  and (_02962_, _02961_, _02956_);
  and (_02963_, _02962_, _02951_);
  and (_02964_, _02963_, _02937_);
  or (_02965_, _02909_, _42338_);
  or (_02966_, _02913_, _42297_);
  and (_02967_, _02966_, _02965_);
  or (_02968_, _02918_, _42174_);
  or (_02969_, _02920_, _42133_);
  and (_02970_, _02969_, _02968_);
  and (_02971_, _02970_, _02967_);
  or (_02972_, _02925_, _42502_);
  or (_02973_, _02927_, _42461_);
  and (_02974_, _02973_, _02972_);
  or (_02975_, _02931_, _42010_);
  or (_02976_, _02933_, _41961_);
  and (_02977_, _02976_, _02975_);
  and (_02978_, _02977_, _02974_);
  and (_02979_, _02978_, _02971_);
  or (_02980_, _02940_, _42420_);
  or (_02981_, _02943_, _42379_);
  and (_02982_, _02981_, _02980_);
  or (_02983_, _02946_, _41872_);
  or (_02984_, _02948_, _41913_);
  and (_02985_, _02984_, _02983_);
  and (_02986_, _02985_, _02982_);
  or (_02987_, _02952_, _42256_);
  or (_02988_, _02954_, _42215_);
  and (_02989_, _02988_, _02987_);
  or (_02990_, _02957_, _42092_);
  or (_02991_, _02959_, _42051_);
  and (_02992_, _02991_, _02990_);
  and (_02993_, _02992_, _02989_);
  and (_02994_, _02993_, _02986_);
  and (_02995_, _02994_, _02979_);
  and (_02996_, _02995_, _02964_);
  or (_02997_, _02909_, _42363_);
  or (_02998_, _02913_, _42322_);
  and (_02999_, _02998_, _02997_);
  or (_03000_, _02918_, _42199_);
  or (_03001_, _02920_, _42158_);
  and (_03003_, _03001_, _03000_);
  and (_03004_, _03003_, _02999_);
  or (_03005_, _02925_, _42527_);
  or (_03006_, _02927_, _42486_);
  and (_03007_, _03006_, _03005_);
  or (_03008_, _02931_, _42035_);
  or (_03009_, _02933_, _41994_);
  and (_03010_, _03009_, _03008_);
  and (_03011_, _03010_, _03007_);
  and (_03012_, _03011_, _03004_);
  or (_03014_, _02940_, _42445_);
  or (_03015_, _02943_, _42404_);
  and (_03016_, _03015_, _03014_);
  or (_03017_, _02946_, _41897_);
  or (_03018_, _02948_, _41943_);
  and (_03019_, _03018_, _03017_);
  and (_03020_, _03019_, _03016_);
  or (_03021_, _02952_, _42281_);
  or (_03022_, _02954_, _42240_);
  and (_03023_, _03022_, _03021_);
  or (_03024_, _02957_, _42117_);
  or (_03025_, _02959_, _42076_);
  and (_03026_, _03025_, _03024_);
  and (_03027_, _03026_, _03023_);
  and (_03028_, _03027_, _03020_);
  and (_03029_, _03028_, _03012_);
  or (_03030_, _02909_, _42368_);
  or (_03031_, _02913_, _42327_);
  and (_03032_, _03031_, _03030_);
  or (_03033_, _02918_, _42204_);
  or (_03035_, _02920_, _42163_);
  and (_03036_, _03035_, _03033_);
  and (_03037_, _03036_, _03032_);
  or (_03038_, _02925_, _42532_);
  or (_03039_, _02927_, _42491_);
  and (_03040_, _03039_, _03038_);
  or (_03041_, _02931_, _42040_);
  or (_03042_, _02933_, _41999_);
  and (_03043_, _03042_, _03041_);
  and (_03044_, _03043_, _03040_);
  and (_03046_, _03044_, _03037_);
  or (_03047_, _02940_, _42450_);
  or (_03048_, _02943_, _42409_);
  and (_03049_, _03048_, _03047_);
  or (_03050_, _02946_, _41902_);
  or (_03051_, _02948_, _41950_);
  and (_03052_, _03051_, _03050_);
  and (_03053_, _03052_, _03049_);
  or (_03054_, _02952_, _42286_);
  or (_03055_, _02954_, _42245_);
  and (_03057_, _03055_, _03054_);
  or (_03058_, _02957_, _42122_);
  or (_03059_, _02959_, _42081_);
  and (_03060_, _03059_, _03058_);
  and (_03061_, _03060_, _03057_);
  and (_03062_, _03061_, _03053_);
  nand (_03063_, _03062_, _03046_);
  or (_03064_, _03063_, _03029_);
  not (_03065_, _03064_);
  and (_03066_, _03065_, _02996_);
  or (_03067_, _02909_, _42353_);
  or (_03068_, _02913_, _42312_);
  and (_03069_, _03068_, _03067_);
  or (_03070_, _02918_, _42189_);
  or (_03071_, _02920_, _42148_);
  and (_03072_, _03071_, _03070_);
  and (_03073_, _03072_, _03069_);
  or (_03074_, _02925_, _42517_);
  or (_03075_, _02927_, _42476_);
  and (_03076_, _03075_, _03074_);
  or (_03078_, _02931_, _42025_);
  or (_03079_, _02933_, _41976_);
  and (_03080_, _03079_, _03078_);
  and (_03081_, _03080_, _03076_);
  and (_03082_, _03081_, _03073_);
  or (_03083_, _02940_, _42435_);
  or (_03084_, _02943_, _42394_);
  and (_03085_, _03084_, _03083_);
  or (_03086_, _02946_, _41887_);
  or (_03087_, _02948_, _41928_);
  and (_03089_, _03087_, _03086_);
  and (_03090_, _03089_, _03085_);
  or (_03091_, _02952_, _42271_);
  or (_03092_, _02954_, _42230_);
  and (_03093_, _03092_, _03091_);
  or (_03094_, _02957_, _42107_);
  or (_03095_, _02959_, _42066_);
  and (_03096_, _03095_, _03094_);
  and (_03097_, _03096_, _03093_);
  and (_03098_, _03097_, _03090_);
  nand (_03100_, _03098_, _03082_);
  or (_03101_, _02909_, _42358_);
  or (_03102_, _02913_, _42317_);
  and (_03103_, _03102_, _03101_);
  or (_03104_, _02918_, _42194_);
  or (_03105_, _02920_, _42153_);
  and (_03106_, _03105_, _03104_);
  and (_03107_, _03106_, _03103_);
  or (_03108_, _02925_, _42522_);
  or (_03109_, _02927_, _42481_);
  and (_03111_, _03109_, _03108_);
  or (_03112_, _02931_, _42030_);
  or (_03113_, _02933_, _41986_);
  and (_03114_, _03113_, _03112_);
  and (_03115_, _03114_, _03111_);
  and (_03116_, _03115_, _03107_);
  or (_03117_, _02940_, _42440_);
  or (_03118_, _02943_, _42399_);
  and (_03119_, _03118_, _03117_);
  or (_03120_, _02946_, _41892_);
  or (_03122_, _02948_, _41934_);
  and (_03123_, _03122_, _03120_);
  and (_03124_, _03123_, _03119_);
  or (_03125_, _02952_, _42276_);
  or (_03126_, _02954_, _42235_);
  and (_03127_, _03126_, _03125_);
  or (_03128_, _02957_, _42112_);
  or (_03129_, _02959_, _42071_);
  and (_03130_, _03129_, _03128_);
  and (_03131_, _03130_, _03127_);
  and (_03133_, _03131_, _03124_);
  nand (_03134_, _03133_, _03116_);
  or (_03135_, _03134_, _03100_);
  not (_03136_, _03135_);
  or (_03137_, _02909_, _42343_);
  or (_03138_, _02913_, _42302_);
  and (_03139_, _03138_, _03137_);
  or (_03140_, _02918_, _42179_);
  or (_03141_, _02920_, _42138_);
  and (_03142_, _03141_, _03140_);
  and (_03144_, _03142_, _03139_);
  or (_03145_, _02925_, _42507_);
  or (_03146_, _02927_, _42466_);
  and (_03147_, _03146_, _03145_);
  or (_03148_, _02931_, _42015_);
  or (_03149_, _02933_, _41966_);
  and (_03150_, _03149_, _03148_);
  and (_03151_, _03150_, _03147_);
  and (_03152_, _03151_, _03144_);
  or (_03153_, _02940_, _42425_);
  or (_03155_, _02943_, _42384_);
  and (_03156_, _03155_, _03153_);
  or (_03157_, _02946_, _41877_);
  or (_03158_, _02948_, _41918_);
  and (_03159_, _03158_, _03157_);
  and (_03160_, _03159_, _03156_);
  or (_03161_, _02952_, _42261_);
  or (_03162_, _02954_, _42220_);
  and (_03163_, _03162_, _03161_);
  or (_03164_, _02957_, _42097_);
  or (_03166_, _02959_, _42056_);
  and (_03167_, _03166_, _03164_);
  and (_03168_, _03167_, _03163_);
  and (_03169_, _03168_, _03160_);
  and (_03170_, _03169_, _03152_);
  or (_03171_, _02909_, _42348_);
  or (_03172_, _02913_, _42307_);
  and (_03173_, _03172_, _03171_);
  or (_03174_, _02918_, _42184_);
  or (_03175_, _02920_, _42143_);
  and (_03176_, _03175_, _03174_);
  and (_03177_, _03176_, _03173_);
  or (_03178_, _02925_, _42512_);
  or (_03179_, _02927_, _42471_);
  and (_03180_, _03179_, _03178_);
  or (_03181_, _02931_, _42020_);
  or (_03182_, _02933_, _41971_);
  and (_03183_, _03182_, _03181_);
  and (_03184_, _03183_, _03180_);
  and (_03185_, _03184_, _03177_);
  or (_03186_, _02940_, _42430_);
  or (_03187_, _02943_, _42389_);
  and (_03188_, _03187_, _03186_);
  or (_03189_, _02946_, _41882_);
  or (_03190_, _02948_, _41923_);
  and (_03191_, _03190_, _03189_);
  and (_03192_, _03191_, _03188_);
  or (_03193_, _02952_, _42266_);
  or (_03194_, _02954_, _42225_);
  and (_03195_, _03194_, _03193_);
  or (_03196_, _02957_, _42102_);
  or (_03197_, _02959_, _42061_);
  and (_03198_, _03197_, _03196_);
  and (_03199_, _03198_, _03195_);
  and (_03200_, _03199_, _03192_);
  nand (_03201_, _03200_, _03185_);
  not (_03202_, _03201_);
  and (_03203_, _03202_, _03170_);
  and (_03204_, _03203_, _03136_);
  and (_03205_, _03204_, _03066_);
  not (_03206_, _03205_);
  nor (_03207_, _02924_, _02911_);
  and (_03208_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03209_, _03208_, \oc8051_golden_model_1.PC [3]);
  nor (_03210_, _03209_, _03207_);
  not (_03211_, _03210_);
  or (_03212_, _03201_, _03170_);
  or (_03213_, _03212_, _03135_);
  not (_03214_, _03213_);
  nand (_03215_, _03028_, _03012_);
  or (_03216_, _03063_, _03215_);
  nand (_03217_, _02963_, _02937_);
  or (_03218_, _02995_, _03217_);
  nor (_03219_, _03218_, _03216_);
  and (_03220_, _03219_, _03214_);
  not (_03221_, _03220_);
  and (_03222_, _02995_, _03217_);
  and (_03223_, _03062_, _03046_);
  or (_03224_, _03223_, _03029_);
  not (_03225_, _03224_);
  and (_03226_, _03225_, _03222_);
  and (_03227_, _03226_, _03214_);
  or (_03228_, _03223_, _03215_);
  not (_03229_, _03228_);
  and (_03230_, _03222_, _03229_);
  and (_03231_, _03230_, _03214_);
  nor (_03232_, _03231_, _03227_);
  and (_03233_, _03232_, _03221_);
  not (_03234_, _03216_);
  and (_03235_, _03222_, _03234_);
  and (_03236_, _03235_, _03214_);
  and (_03237_, _03222_, _03065_);
  and (_03238_, _03237_, _03214_);
  nor (_03239_, _03238_, _03236_);
  and (_03240_, _03239_, _03233_);
  and (_03241_, _03234_, _02996_);
  and (_03242_, _03241_, _03214_);
  and (_03243_, _03214_, _03066_);
  nor (_03244_, _03243_, _03242_);
  and (_03245_, _03229_, _02996_);
  and (_03246_, _03245_, _03214_);
  and (_03247_, _03225_, _02996_);
  and (_03248_, _03247_, _03214_);
  nor (_03249_, _03248_, _03246_);
  and (_03250_, _03249_, _03244_);
  and (_03251_, _03250_, _03240_);
  or (_03252_, _03218_, _03224_);
  or (_03253_, _03252_, _03213_);
  or (_03254_, _02995_, _02964_);
  or (_03255_, _03254_, _03064_);
  or (_03257_, _03255_, _03213_);
  and (_03258_, _03257_, _03253_);
  or (_03259_, _03254_, _03216_);
  or (_03260_, _03259_, _03213_);
  or (_03261_, _03254_, _03228_);
  or (_03262_, _03261_, _03213_);
  and (_03263_, _03262_, _03260_);
  or (_03264_, _03218_, _03228_);
  or (_03265_, _03264_, _03213_);
  or (_03266_, _03254_, _03224_);
  or (_03267_, _03266_, _03213_);
  and (_03268_, _03267_, _03265_);
  and (_03269_, _03268_, _03263_);
  and (_03270_, _03269_, _03258_);
  not (_03271_, _03219_);
  not (_03272_, _03100_);
  or (_03273_, _03134_, _03272_);
  or (_03274_, _03273_, _03212_);
  or (_03275_, _03274_, _03271_);
  nor (_03276_, _03218_, _03064_);
  not (_03277_, _03276_);
  or (_03278_, _03277_, _03213_);
  and (_03279_, _03278_, _03275_);
  and (_03280_, _03279_, _03270_);
  nand (_03281_, _03280_, _03251_);
  nand (_03282_, _03281_, _03211_);
  or (_03283_, _03202_, _03170_);
  or (_03284_, _03283_, _03135_);
  or (_03285_, _03284_, _03277_);
  and (_03286_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  and (_03287_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_03288_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03289_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_03290_, _03289_, _03287_);
  and (_03291_, _03290_, _03288_);
  nor (_03292_, _03291_, _03287_);
  nor (_03293_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_03294_, _03293_, _03286_);
  not (_03295_, _03294_);
  nor (_03296_, _03295_, _03292_);
  nor (_03297_, _03296_, _03286_);
  and (_03298_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03299_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_03300_, _03299_, _03298_);
  not (_03301_, _03300_);
  nor (_03302_, _03301_, _03297_);
  and (_03303_, _03301_, _03297_);
  nor (_03304_, _03303_, _03302_);
  or (_03305_, _03304_, _03285_);
  not (_03306_, _02918_);
  nor (_03307_, _02906_, _02916_);
  nor (_03308_, _03307_, _02907_);
  nor (_03309_, _03308_, _03306_);
  and (_03310_, _03285_, _03309_);
  nand (_03311_, _03310_, _03270_);
  nand (_03312_, _03311_, _03305_);
  nor (_03313_, _03284_, _03271_);
  not (_03314_, _03313_);
  and (_03315_, _03314_, _03279_);
  and (_03316_, _03315_, _03312_);
  and (_03317_, _02906_, _02916_);
  nor (_03318_, _03317_, _03307_);
  and (_03319_, _03318_, \oc8051_golden_model_1.ACC [2]);
  not (_03320_, \oc8051_golden_model_1.ACC [1]);
  and (_03321_, _02939_, _02912_);
  nor (_03322_, _03321_, _03320_);
  and (_03323_, \oc8051_golden_model_1.ACC [0], _02938_);
  and (_03324_, _03321_, _03320_);
  nor (_03325_, _03324_, _03322_);
  and (_03326_, _03325_, _03323_);
  nor (_03327_, _03326_, _03322_);
  nor (_03328_, _03318_, \oc8051_golden_model_1.ACC [2]);
  nor (_03329_, _03328_, _03319_);
  not (_03330_, _03329_);
  nor (_03331_, _03330_, _03327_);
  nor (_03332_, _03331_, _03319_);
  nor (_03333_, _03309_, \oc8051_golden_model_1.ACC [3]);
  and (_03334_, _03309_, \oc8051_golden_model_1.ACC [3]);
  nor (_03335_, _03334_, _03333_);
  and (_03336_, _03335_, _03332_);
  nor (_03337_, _03335_, _03332_);
  nor (_03338_, _03337_, _03336_);
  nor (_03339_, _03338_, _03314_);
  or (_03340_, _03339_, _03316_);
  nand (_03341_, _03340_, _03251_);
  nand (_03342_, _03341_, _03282_);
  and (_03343_, _03330_, _03327_);
  nor (_03344_, _03343_, _03331_);
  and (_03345_, _03344_, _03313_);
  and (_03346_, _03295_, _03292_);
  nor (_03347_, _03346_, _03296_);
  not (_03348_, _03347_);
  or (_03349_, _03348_, _03285_);
  and (_03350_, _03349_, _03279_);
  nand (_03351_, _03269_, _03258_);
  or (_03352_, _03318_, _03351_);
  nand (_03353_, _03352_, _03285_);
  nand (_03354_, _03353_, _03350_);
  nor (_03355_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_03356_, _03355_, _03208_);
  or (_03357_, _03356_, _03280_);
  and (_03358_, _03357_, _03314_);
  and (_03359_, _03358_, _03354_);
  or (_03360_, _03359_, _03345_);
  nand (_03361_, _03360_, _03251_);
  not (_03362_, _03356_);
  or (_03363_, _03362_, _03251_);
  and (_03364_, _03363_, _03361_);
  or (_03365_, _03364_, _03342_);
  or (_03366_, _03251_, _02911_);
  or (_03367_, _03270_, \oc8051_golden_model_1.PC [1]);
  or (_03368_, _03321_, _03351_);
  nand (_03369_, _03368_, _03367_);
  nand (_03370_, _03369_, _03285_);
  not (_03371_, _03285_);
  nor (_03372_, _03290_, _03288_);
  nor (_03373_, _03372_, _03291_);
  nand (_03374_, _03373_, _03371_);
  and (_03375_, _03374_, _03279_);
  nand (_03376_, _03375_, _03370_);
  or (_03377_, _03279_, _02911_);
  and (_03378_, _03377_, _03314_);
  nand (_03379_, _03378_, _03376_);
  not (_03380_, _03251_);
  nor (_03381_, _03325_, _03323_);
  nor (_03382_, _03381_, _03326_);
  and (_03383_, _03382_, _03313_);
  nor (_03384_, _03383_, _03380_);
  nand (_03385_, _03384_, _03379_);
  nand (_03386_, _03385_, _03366_);
  nor (_03387_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_03388_, _03387_, _03288_);
  nand (_03389_, _03388_, _03371_);
  and (_03390_, _03285_, _02938_);
  nand (_03391_, _03390_, _03270_);
  nand (_03392_, _03391_, _03389_);
  nand (_03393_, _03392_, _03279_);
  or (_03394_, _03280_, _02938_);
  nand (_03395_, _03394_, _03393_);
  nand (_03396_, _03395_, _03314_);
  not (_03397_, \oc8051_golden_model_1.ACC [0]);
  and (_03398_, _03397_, \oc8051_golden_model_1.PC [0]);
  nor (_03399_, _03398_, _03323_);
  and (_03400_, _03399_, _03313_);
  nor (_03401_, _03400_, _03380_);
  nand (_03402_, _03401_, _03396_);
  or (_03403_, _03251_, \oc8051_golden_model_1.PC [0]);
  nand (_03404_, _03403_, _03402_);
  or (_03405_, _03404_, _03386_);
  or (_03406_, _03405_, _03365_);
  or (_03407_, _03406_, _42502_);
  and (_03408_, _03385_, _03366_);
  or (_03409_, _03404_, _03408_);
  nand (_03410_, _03363_, _03361_);
  or (_03411_, _03410_, _03342_);
  or (_03412_, _03411_, _03409_);
  or (_03413_, _03412_, _42256_);
  and (_03414_, _03413_, _03407_);
  and (_03415_, _03341_, _03282_);
  or (_03416_, _03364_, _03415_);
  or (_03417_, _03416_, _03409_);
  or (_03418_, _03417_, _42092_);
  or (_03419_, _03410_, _03415_);
  or (_03420_, _03419_, _03409_);
  or (_03421_, _03420_, _41913_);
  and (_03422_, _03421_, _03418_);
  and (_03423_, _03422_, _03414_);
  or (_03424_, _03416_, _03405_);
  or (_03425_, _03424_, _42174_);
  and (_03426_, _03403_, _03402_);
  or (_03427_, _03426_, _03408_);
  or (_03428_, _03416_, _03427_);
  or (_03429_, _03428_, _42051_);
  and (_03430_, _03429_, _03425_);
  or (_03431_, _03409_, _03365_);
  or (_03432_, _03431_, _42420_);
  or (_03433_, _03427_, _03365_);
  or (_03434_, _03433_, _42379_);
  and (_03435_, _03434_, _03432_);
  and (_03436_, _03435_, _03430_);
  and (_03437_, _03436_, _03423_);
  or (_03438_, _03426_, _03386_);
  or (_03439_, _03411_, _03438_);
  or (_03440_, _03439_, _42297_);
  or (_03441_, _03411_, _03427_);
  or (_03442_, _03441_, _42215_);
  and (_03443_, _03442_, _03440_);
  or (_03444_, _03419_, _03405_);
  or (_03445_, _03444_, _42010_);
  or (_03446_, _03419_, _03427_);
  or (_03447_, _03446_, _41872_);
  and (_03448_, _03447_, _03445_);
  and (_03449_, _03448_, _03443_);
  or (_03450_, _03438_, _03365_);
  or (_03451_, _03450_, _42461_);
  or (_03452_, _03416_, _03438_);
  or (_03453_, _03452_, _42133_);
  and (_03454_, _03453_, _03451_);
  or (_03455_, _03411_, _03405_);
  or (_03456_, _03455_, _42338_);
  or (_03458_, _03419_, _03438_);
  or (_03459_, _03458_, _41961_);
  and (_03460_, _03459_, _03456_);
  and (_03461_, _03460_, _03454_);
  and (_03462_, _03461_, _03449_);
  nand (_03463_, _03462_, _03437_);
  or (_03464_, _03431_, _42440_);
  or (_03465_, _03424_, _42194_);
  and (_03466_, _03465_, _03464_);
  or (_03467_, _03452_, _42153_);
  or (_03468_, _03446_, _41892_);
  and (_03469_, _03468_, _03467_);
  and (_03470_, _03469_, _03466_);
  or (_03471_, _03412_, _42276_);
  or (_03472_, _03439_, _42317_);
  and (_03473_, _03472_, _03471_);
  or (_03474_, _03455_, _42358_);
  or (_03475_, _03444_, _42030_);
  and (_03476_, _03475_, _03474_);
  and (_03477_, _03476_, _03473_);
  and (_03478_, _03477_, _03470_);
  or (_03479_, _03417_, _42112_);
  or (_03480_, _03428_, _42071_);
  and (_03481_, _03480_, _03479_);
  or (_03482_, _03450_, _42481_);
  or (_03483_, _03420_, _41934_);
  and (_03484_, _03483_, _03482_);
  and (_03485_, _03484_, _03481_);
  or (_03486_, _03406_, _42522_);
  or (_03487_, _03458_, _41986_);
  and (_03488_, _03487_, _03486_);
  or (_03489_, _03433_, _42399_);
  or (_03490_, _03441_, _42235_);
  and (_03491_, _03490_, _03489_);
  and (_03492_, _03491_, _03488_);
  and (_03493_, _03492_, _03485_);
  and (_03494_, _03493_, _03478_);
  or (_03495_, _03494_, _03463_);
  nor (_03496_, _03495_, _03206_);
  not (_03497_, _03278_);
  and (_03498_, _03201_, _03170_);
  and (_03499_, _03498_, _03136_);
  and (_03500_, _03499_, _03276_);
  not (_03501_, _03500_);
  nor (_03502_, _03501_, _03495_);
  not (_03503_, _03252_);
  and (_03504_, _03499_, _03503_);
  not (_03505_, _03504_);
  nor (_03506_, _03505_, _03495_);
  nor (_03507_, _03505_, _03463_);
  not (_03508_, _03507_);
  not (_03509_, _03259_);
  and (_03510_, _03509_, _03204_);
  and (_03511_, _03499_, _03509_);
  not (_03512_, _03511_);
  nor (_03513_, _03512_, _03495_);
  not (_03514_, _03255_);
  and (_03515_, _03499_, _03514_);
  not (_03516_, _03515_);
  or (_03517_, _03516_, _03495_);
  not (_03518_, _03267_);
  and (_03519_, _03245_, _03204_);
  not (_03520_, _03519_);
  and (_03521_, _03499_, _03245_);
  not (_03522_, _03521_);
  not (_03523_, _03274_);
  and (_03524_, _03523_, _03245_);
  not (_03525_, _03524_);
  nor (_03526_, _03424_, _42209_);
  nor (_03527_, _03420_, _41955_);
  nor (_03528_, _03527_, _03526_);
  nor (_03529_, _03441_, _42250_);
  nor (_03530_, _03444_, _42045_);
  nor (_03531_, _03530_, _03529_);
  and (_03532_, _03531_, _03528_);
  nor (_03533_, _03455_, _42373_);
  nor (_03534_, _03446_, _41907_);
  nor (_03535_, _03534_, _03533_);
  nor (_03536_, _03431_, _42455_);
  nor (_03537_, _03433_, _42414_);
  nor (_03538_, _03537_, _03536_);
  and (_03539_, _03538_, _03535_);
  and (_03540_, _03539_, _03532_);
  nor (_03541_, _03450_, _42496_);
  nor (_03542_, _03458_, _42004_);
  nor (_03543_, _03542_, _03541_);
  nor (_03544_, _03412_, _42291_);
  nor (_03545_, _03452_, _42168_);
  nor (_03546_, _03545_, _03544_);
  and (_03547_, _03546_, _03543_);
  nor (_03548_, _03439_, _42332_);
  nor (_03549_, _03428_, _42086_);
  nor (_03550_, _03549_, _03548_);
  nor (_03551_, _03406_, _42537_);
  nor (_03552_, _03417_, _42127_);
  nor (_03553_, _03552_, _03551_);
  and (_03554_, _03553_, _03550_);
  and (_03555_, _03554_, _03547_);
  and (_03556_, _03555_, _03540_);
  nor (_03557_, _03556_, _03463_);
  not (_03558_, _03494_);
  and (_03559_, _03558_, _03463_);
  nor (_03560_, _03559_, _03557_);
  and (_03561_, _03499_, _03226_);
  and (_03562_, _03499_, _03219_);
  nor (_03563_, _03562_, _03561_);
  not (_03564_, _03563_);
  and (_03565_, _03564_, _03560_);
  not (_03566_, _03264_);
  and (_03567_, _03134_, _03272_);
  and (_03568_, _03567_, _03498_);
  and (_03569_, _03568_, _03566_);
  and (_03570_, _03567_, _03203_);
  and (_03571_, _03570_, _03566_);
  nor (_03572_, _03571_, _03569_);
  not (_03573_, _03212_);
  and (_03574_, _03134_, _03100_);
  and (_03575_, _03574_, _03573_);
  and (_03576_, _03575_, _03566_);
  and (_03577_, _03574_, _03498_);
  and (_03578_, _03577_, _03566_);
  nor (_03579_, _03578_, _03576_);
  and (_03580_, _03579_, _03572_);
  not (_03581_, _03283_);
  and (_03582_, _03574_, _03581_);
  and (_03583_, _03582_, _03566_);
  and (_03584_, _03567_, _03581_);
  and (_03585_, _03584_, _03566_);
  nor (_03586_, _03585_, _03583_);
  and (_03587_, _03574_, _03203_);
  and (_03588_, _03587_, _03566_);
  and (_03589_, _03567_, _03573_);
  and (_03590_, _03589_, _03566_);
  nor (_03591_, _03590_, _03588_);
  and (_03592_, _03591_, _03586_);
  and (_03593_, _03592_, _03580_);
  not (_03594_, _03593_);
  and (_03595_, _03515_, _03560_);
  not (_03596_, \oc8051_golden_model_1.SP [3]);
  and (_03597_, _03514_, _03204_);
  and (_03598_, _03597_, _03596_);
  nor (_03599_, _03274_, _03255_);
  nor (_03600_, _03274_, _03261_);
  nor (_03601_, _03600_, _03599_);
  or (_03602_, _03601_, _03494_);
  nor (_03603_, _03274_, _03259_);
  nor (_03604_, _03597_, _03515_);
  nand (_03605_, _03601_, \oc8051_golden_model_1.PSW [3]);
  and (_03606_, _03605_, _03604_);
  or (_03607_, _03606_, _03603_);
  and (_03608_, _03607_, _03602_);
  or (_03609_, _03608_, _03598_);
  or (_03610_, _03609_, _03595_);
  not (_03611_, _03603_);
  or (_03612_, _03611_, _03494_);
  and (_03613_, _03612_, _03610_);
  or (_03614_, _03613_, _03511_);
  nor (_03615_, _03274_, _03252_);
  nor (_03616_, _03615_, _03510_);
  or (_03617_, _03560_, _03512_);
  and (_03618_, _03617_, _03616_);
  and (_03619_, _03618_, _03614_);
  nor (_03620_, _03616_, _03558_);
  and (_03621_, _03503_, _03204_);
  nor (_03622_, _03504_, _03621_);
  not (_03623_, _03622_);
  or (_03624_, _03623_, _03620_);
  or (_03625_, _03624_, _03619_);
  or (_03626_, _03622_, _03560_);
  and (_03627_, _03626_, _03625_);
  or (_03628_, _03627_, _03594_);
  and (_03629_, _03566_, _03204_);
  and (_03630_, _03499_, _03566_);
  nor (_03631_, _03630_, _03629_);
  or (_03632_, _03593_, _03494_);
  and (_03633_, _03632_, _03631_);
  and (_03634_, _03633_, _03628_);
  nor (_03635_, _03277_, _03274_);
  not (_03636_, _03631_);
  and (_03637_, _03636_, _03560_);
  or (_03638_, _03637_, _03635_);
  or (_03639_, _03638_, _03634_);
  not (_03640_, _03635_);
  or (_03641_, _03640_, _03494_);
  and (_03642_, _03641_, _03501_);
  and (_03643_, _03642_, _03639_);
  not (_03644_, _03275_);
  and (_03645_, _03560_, _03500_);
  or (_03646_, _03645_, _03644_);
  or (_03647_, _03646_, _03643_);
  not (_03648_, _03284_);
  and (_03649_, _03648_, _03230_);
  and (_03650_, _03523_, _03226_);
  nor (_03651_, _03650_, _03649_);
  and (_03652_, _03247_, _03204_);
  and (_03653_, _03648_, _03235_);
  nor (_03654_, _03653_, _03652_);
  and (_03655_, _03648_, _03237_);
  and (_03656_, _03276_, _03204_);
  nor (_03657_, _03656_, _03655_);
  and (_03659_, _03657_, _03654_);
  and (_03660_, _03659_, _03651_);
  and (_03661_, _03575_, _03503_);
  and (_03662_, _03577_, _03503_);
  nor (_03663_, _03662_, _03661_);
  and (_03664_, _03587_, _03503_);
  not (_03665_, _03664_);
  and (_03666_, _03567_, _03202_);
  and (_03667_, _03666_, _03503_);
  and (_03668_, _03567_, _03201_);
  and (_03669_, _03668_, _03503_);
  nor (_03670_, _03669_, _03667_);
  and (_03671_, _03670_, _03665_);
  and (_03672_, _03671_, _03663_);
  and (_03673_, _03672_, _03660_);
  not (_03674_, _03273_);
  and (_03675_, _03674_, _03203_);
  and (_03676_, _03675_, _03503_);
  and (_03677_, _03498_, _03674_);
  and (_03678_, _03677_, _03503_);
  nor (_03679_, _03678_, _03676_);
  nor (_03680_, _03283_, _03273_);
  and (_03681_, _03680_, _03503_);
  nor (_03682_, _03681_, _03615_);
  and (_03683_, _03682_, _03679_);
  and (_03684_, _03499_, _03241_);
  nor (_03685_, _03684_, _03205_);
  and (_03686_, _03499_, _03066_);
  nor (_03687_, _03686_, _03519_);
  and (_03688_, _03687_, _03685_);
  not (_03689_, _03170_);
  and (_03690_, _03574_, _03201_);
  and (_03691_, _03690_, _03503_);
  and (_03692_, _03691_, _03689_);
  nor (_03693_, _03692_, _03599_);
  and (_03694_, _03693_, _03688_);
  and (_03695_, _03694_, _03683_);
  and (_03696_, _03695_, _03673_);
  nor (_03697_, _03696_, _03362_);
  and (_03698_, _03696_, _03318_);
  nor (_03699_, _03698_, _03697_);
  nor (_03700_, _03696_, _03211_);
  not (_03701_, _03309_);
  and (_03702_, _03696_, _03701_);
  nor (_03703_, _03702_, _03700_);
  nor (_03704_, _03703_, _03699_);
  nor (_03705_, _03696_, _02938_);
  and (_03706_, _03696_, _02938_);
  nor (_03707_, _03706_, _03705_);
  nor (_03708_, _03706_, \oc8051_golden_model_1.PC [1]);
  and (_03709_, _03706_, \oc8051_golden_model_1.PC [1]);
  nor (_03710_, _03709_, _03708_);
  nor (_03711_, _03710_, _03707_);
  and (_03712_, _03711_, _03704_);
  and (_03713_, _03712_, _02067_);
  and (_03714_, _03710_, _03707_);
  and (_03715_, _03703_, _03699_);
  and (_03716_, _03715_, _03714_);
  and (_03717_, _03716_, _02074_);
  nor (_03718_, _03717_, _03713_);
  not (_03719_, _03699_);
  nor (_03720_, _03703_, _03719_);
  and (_03721_, _03720_, _03711_);
  and (_03722_, _03721_, _02112_);
  not (_03723_, _03707_);
  and (_03724_, _03710_, _03723_);
  and (_03725_, _03715_, _03724_);
  and (_03726_, _03725_, _02087_);
  nor (_03727_, _03726_, _03722_);
  and (_03728_, _03727_, _03718_);
  and (_03729_, _03720_, _03724_);
  and (_03730_, _03729_, _02110_);
  nor (_03731_, _03710_, _03723_);
  and (_03732_, _03715_, _03731_);
  and (_03733_, _03732_, _02085_);
  nor (_03734_, _03733_, _03730_);
  and (_03735_, _03703_, _03719_);
  and (_03736_, _03735_, _03731_);
  and (_03737_, _03736_, _02071_);
  and (_03738_, _03735_, _03714_);
  and (_03739_, _03738_, _02098_);
  nor (_03740_, _03739_, _03737_);
  and (_03741_, _03740_, _03734_);
  and (_03742_, _03741_, _03728_);
  and (_03743_, _03735_, _03724_);
  and (_03744_, _03743_, _02069_);
  and (_03745_, _03715_, _03711_);
  and (_03746_, _03745_, _02090_);
  nor (_03747_, _03746_, _03744_);
  and (_03748_, _03731_, _03704_);
  and (_03749_, _03748_, _02064_);
  and (_03750_, _03720_, _03731_);
  and (_03751_, _03750_, _02095_);
  nor (_03752_, _03751_, _03749_);
  and (_03753_, _03752_, _03747_);
  and (_03754_, _03714_, _03704_);
  and (_03755_, _03754_, _02103_);
  and (_03756_, _03714_, _03720_);
  and (_03757_, _03756_, _02101_);
  nor (_03758_, _03757_, _03755_);
  and (_03759_, _03724_, _03704_);
  and (_03760_, _03759_, _02062_);
  and (_03761_, _03735_, _03711_);
  and (_03762_, _03761_, _02076_);
  nor (_03763_, _03762_, _03760_);
  and (_03764_, _03763_, _03758_);
  and (_03765_, _03764_, _03753_);
  and (_03766_, _03765_, _03742_);
  or (_03767_, _03766_, _03275_);
  and (_03768_, _03767_, _03563_);
  and (_03769_, _03768_, _03647_);
  or (_03770_, _03769_, _03565_);
  and (_03771_, _03523_, _03237_);
  not (_03772_, _03771_);
  and (_03773_, _03499_, _03237_);
  nor (_03774_, _03773_, _03655_);
  and (_03775_, _03774_, _03772_);
  and (_03776_, _03523_, _03230_);
  not (_03777_, _03776_);
  and (_03778_, _03499_, _03230_);
  nor (_03779_, _03778_, _03649_);
  and (_03780_, _03779_, _03777_);
  and (_03781_, _03780_, _03775_);
  and (_03782_, _03523_, _03247_);
  not (_03783_, _03782_);
  and (_03784_, _03523_, _03235_);
  not (_03785_, _03784_);
  and (_03786_, _03499_, _03235_);
  nor (_03787_, _03786_, _03653_);
  and (_03788_, _03787_, _03785_);
  and (_03789_, _03788_, _03783_);
  and (_03790_, _03789_, _03781_);
  and (_03791_, _03790_, _03770_);
  and (_03792_, _03499_, _03247_);
  nor (_03793_, _03790_, _03558_);
  or (_03794_, _03793_, _03792_);
  or (_03795_, _03794_, _03791_);
  not (_03796_, _03652_);
  nand (_03797_, _03792_, \oc8051_golden_model_1.SP [3]);
  and (_03798_, _03797_, _03796_);
  and (_03799_, _03798_, _03795_);
  and (_03800_, _03652_, _03560_);
  or (_03801_, _03800_, _03799_);
  and (_03802_, _03801_, _03525_);
  and (_03803_, _03524_, _03494_);
  nor (_03804_, _03803_, _03802_);
  and (_03805_, _03804_, _03522_);
  and (_03806_, _03521_, \oc8051_golden_model_1.SP [3]);
  or (_03807_, _03806_, _03805_);
  and (_03808_, _03807_, _03520_);
  and (_03809_, _03523_, _03066_);
  nor (_03810_, _03560_, _03520_);
  or (_03811_, _03810_, _03809_);
  or (_03812_, _03811_, _03808_);
  nand (_03813_, _03809_, _03494_);
  and (_03814_, _03813_, _03812_);
  nor (_03815_, _03814_, _03205_);
  and (_03816_, _03523_, _03241_);
  and (_03817_, _03560_, _03205_);
  or (_03818_, _03817_, _03816_);
  nor (_03819_, _03818_, _03815_);
  not (_03820_, _03816_);
  nor (_03821_, _03820_, _03494_);
  nor (_03822_, _03821_, _03819_);
  nor (_03823_, _03424_, _42204_);
  nor (_03824_, _03420_, _41950_);
  nor (_03825_, _03824_, _03823_);
  nor (_03826_, _03441_, _42245_);
  nor (_03827_, _03444_, _42040_);
  nor (_03828_, _03827_, _03826_);
  and (_03829_, _03828_, _03825_);
  nor (_03830_, _03455_, _42368_);
  nor (_03831_, _03446_, _41902_);
  nor (_03832_, _03831_, _03830_);
  nor (_03833_, _03431_, _42450_);
  nor (_03834_, _03433_, _42409_);
  nor (_03835_, _03834_, _03833_);
  and (_03836_, _03835_, _03832_);
  and (_03837_, _03836_, _03829_);
  nor (_03838_, _03450_, _42491_);
  nor (_03839_, _03458_, _41999_);
  nor (_03840_, _03839_, _03838_);
  nor (_03841_, _03412_, _42286_);
  nor (_03842_, _03452_, _42163_);
  nor (_03843_, _03842_, _03841_);
  and (_03844_, _03843_, _03840_);
  nor (_03845_, _03439_, _42327_);
  nor (_03846_, _03428_, _42081_);
  nor (_03847_, _03846_, _03845_);
  nor (_03848_, _03406_, _42532_);
  nor (_03849_, _03417_, _42122_);
  nor (_03850_, _03849_, _03848_);
  and (_03851_, _03850_, _03847_);
  and (_03852_, _03851_, _03844_);
  and (_03853_, _03852_, _03837_);
  nor (_03854_, _03853_, _03463_);
  not (_03855_, _03854_);
  nor (_03856_, _03519_, _03205_);
  nor (_03857_, _03515_, _03652_);
  and (_03858_, _03857_, _03856_);
  and (_03860_, _03858_, _03563_);
  and (_03861_, _03631_, _03622_);
  and (_03862_, _03861_, _03501_);
  and (_03863_, _03862_, _03860_);
  nor (_03864_, _03863_, _03855_);
  not (_03865_, _03864_);
  and (_03866_, _03854_, _03511_);
  not (_03867_, _03866_);
  nor (_03868_, _03406_, _42517_);
  nor (_03869_, _03412_, _42271_);
  nor (_03870_, _03869_, _03868_);
  nor (_03871_, _03439_, _42312_);
  nor (_03872_, _03444_, _42025_);
  nor (_03873_, _03872_, _03871_);
  and (_03874_, _03873_, _03870_);
  nor (_03875_, _03450_, _42476_);
  nor (_03876_, _03431_, _42435_);
  nor (_03877_, _03876_, _03875_);
  nor (_03878_, _03424_, _42189_);
  nor (_03879_, _03428_, _42066_);
  nor (_03880_, _03879_, _03878_);
  and (_03881_, _03880_, _03877_);
  and (_03882_, _03881_, _03874_);
  nor (_03883_, _03417_, _42107_);
  nor (_03884_, _03458_, _41976_);
  nor (_03885_, _03884_, _03883_);
  nor (_03886_, _03446_, _41887_);
  nor (_03887_, _03420_, _41928_);
  nor (_03888_, _03887_, _03886_);
  and (_03889_, _03888_, _03885_);
  nor (_03890_, _03433_, _42394_);
  nor (_03891_, _03452_, _42148_);
  nor (_03892_, _03891_, _03890_);
  nor (_03893_, _03455_, _42353_);
  nor (_03894_, _03441_, _42230_);
  nor (_03895_, _03894_, _03893_);
  and (_03896_, _03895_, _03892_);
  and (_03897_, _03896_, _03889_);
  and (_03898_, _03897_, _03882_);
  not (_03899_, _03898_);
  or (_03900_, _03524_, _03782_);
  or (_03901_, _03635_, _03603_);
  nor (_03902_, _03901_, _03900_);
  and (_03903_, _03601_, _03616_);
  and (_03904_, _03903_, _03902_);
  nand (_03905_, _03904_, _03593_);
  nand (_03906_, _03788_, _03780_);
  nor (_03907_, _03816_, _03809_);
  nand (_03908_, _03907_, _03775_);
  or (_03909_, _03908_, _03906_);
  or (_03910_, _03909_, _03905_);
  and (_03911_, _03910_, _03899_);
  not (_03912_, _03911_);
  and (_03913_, _03759_, _02012_);
  and (_03914_, _03721_, _02057_);
  nor (_03915_, _03914_, _03913_);
  and (_03916_, _03738_, _02045_);
  and (_03917_, _03725_, _02031_);
  nor (_03918_, _03917_, _03916_);
  and (_03919_, _03918_, _03915_);
  and (_03920_, _03750_, _02034_);
  and (_03921_, _03729_, _02039_);
  nor (_03922_, _03921_, _03920_);
  and (_03923_, _03748_, _02009_);
  and (_03924_, _03754_, _02042_);
  nor (_03925_, _03924_, _03923_);
  and (_03926_, _03925_, _03922_);
  and (_03927_, _03926_, _03919_);
  and (_03928_, _03761_, _02021_);
  and (_03929_, _03736_, _02019_);
  nor (_03930_, _03929_, _03928_);
  and (_03931_, _03743_, _02014_);
  and (_03932_, _03745_, _02029_);
  nor (_03933_, _03932_, _03931_);
  and (_03934_, _03933_, _03930_);
  and (_03935_, _03712_, _02007_);
  and (_03936_, _03756_, _02047_);
  nor (_03937_, _03936_, _03935_);
  and (_03938_, _03716_, _02016_);
  and (_03939_, _03732_, _02054_);
  nor (_03940_, _03939_, _03938_);
  and (_03941_, _03940_, _03937_);
  and (_03942_, _03941_, _03934_);
  and (_03943_, _03942_, _03927_);
  nor (_03944_, _03943_, _03275_);
  not (_03945_, _03261_);
  and (_03946_, _03690_, _03945_);
  and (_03947_, _03575_, _03945_);
  nor (_03948_, _03947_, _03946_);
  and (_03949_, _03574_, _03202_);
  and (_03950_, _03949_, _03245_);
  and (_03951_, _03574_, _03241_);
  nor (_03952_, _03951_, _03950_);
  and (_03953_, _03690_, _03066_);
  and (_03954_, _03574_, _03235_);
  nor (_03955_, _03954_, _03953_);
  and (_03956_, _03955_, _03952_);
  and (_03957_, _03956_, _03948_);
  and (_03958_, _03574_, _03514_);
  not (_03959_, _03958_);
  and (_03960_, _03587_, _03230_);
  and (_03961_, _03575_, _03230_);
  nor (_03962_, _03961_, _03960_);
  and (_03963_, _03962_, _03959_);
  and (_03964_, _03963_, _03957_);
  and (_03965_, _03575_, _03247_);
  and (_03966_, _03587_, _03945_);
  nor (_03967_, _03966_, _03965_);
  and (_03968_, _03597_, \oc8051_golden_model_1.SP [2]);
  and (_03969_, _03587_, _03247_);
  and (_03970_, _03587_, _03219_);
  or (_03971_, _03970_, _03969_);
  nor (_03972_, _03971_, _03968_);
  and (_03973_, _03972_, _03967_);
  and (_03974_, _03949_, _03503_);
  and (_03975_, _03949_, _03066_);
  nor (_03976_, _03975_, _03974_);
  and (_03977_, _03690_, _03219_);
  and (_03978_, _03949_, _03237_);
  nor (_03979_, _03978_, _03977_);
  and (_03980_, _03979_, _03976_);
  and (_03981_, _03587_, _03276_);
  not (_03982_, _03981_);
  and (_03983_, _03690_, _03230_);
  nor (_03984_, _03983_, _03691_);
  and (_03985_, _03984_, _03982_);
  and (_03986_, _03985_, _03980_);
  and (_03987_, _03986_, _03973_);
  and (_03988_, _03690_, _03245_);
  and (_03989_, _03690_, _03237_);
  nor (_03990_, _03989_, _03988_);
  and (_03991_, _03521_, \oc8051_golden_model_1.SP [2]);
  nor (_03992_, _03218_, _03063_);
  and (_03993_, _03992_, _03575_);
  nor (_03994_, _03993_, _03991_);
  and (_03995_, _03994_, _03990_);
  and (_03996_, _03574_, _03509_);
  not (_03997_, _03996_);
  and (_03998_, _03792_, \oc8051_golden_model_1.SP [2]);
  not (_03999_, _03690_);
  nor (_04000_, _03276_, _03247_);
  nor (_04001_, _04000_, _03999_);
  nor (_04002_, _04001_, _03998_);
  and (_04003_, _04002_, _03997_);
  and (_04004_, _04003_, _03995_);
  and (_04005_, _04004_, _03987_);
  and (_04006_, _04005_, _03964_);
  not (_04007_, _04006_);
  nor (_04008_, _04007_, _03944_);
  and (_04009_, _04008_, _03912_);
  and (_04010_, _04009_, _03867_);
  and (_04011_, _04010_, _03865_);
  or (_04012_, _03444_, _42015_);
  or (_04013_, _03458_, _41966_);
  and (_04014_, _04013_, _04012_);
  or (_04015_, _03455_, _42343_);
  or (_04016_, _03439_, _42302_);
  and (_04017_, _04016_, _04015_);
  and (_04018_, _04017_, _04014_);
  or (_04019_, _03424_, _42179_);
  or (_04020_, _03417_, _42097_);
  and (_04021_, _04020_, _04019_);
  or (_04022_, _03406_, _42507_);
  or (_04023_, _03433_, _42384_);
  and (_04024_, _04023_, _04022_);
  and (_04025_, _04024_, _04021_);
  and (_04026_, _04025_, _04018_);
  or (_04027_, _03412_, _42261_);
  or (_04028_, _03441_, _42220_);
  and (_04029_, _04028_, _04027_);
  or (_04030_, _03450_, _42466_);
  or (_04031_, _03420_, _41918_);
  and (_04032_, _04031_, _04030_);
  and (_04033_, _04032_, _04029_);
  or (_04034_, _03452_, _42138_);
  or (_04035_, _03428_, _42056_);
  and (_04036_, _04035_, _04034_);
  or (_04037_, _03431_, _42425_);
  or (_04038_, _03446_, _41877_);
  and (_04039_, _04038_, _04037_);
  and (_04040_, _04039_, _04036_);
  and (_04041_, _04040_, _04033_);
  and (_04042_, _04041_, _04026_);
  nor (_04043_, _04042_, _03820_);
  not (_04044_, _04043_);
  nor (_04045_, _04042_, _03640_);
  not (_04046_, _03615_);
  nor (_04047_, _04042_, _04046_);
  or (_04048_, _04042_, _03611_);
  nor (_04049_, _04042_, _03601_);
  and (_04050_, _03574_, _03170_);
  nor (_04051_, _03568_, _04050_);
  nor (_04052_, _04051_, _03255_);
  not (_04053_, _04052_);
  and (_04054_, _03677_, _03514_);
  and (_04055_, _03570_, _03514_);
  nor (_04056_, _04055_, _04054_);
  and (_04057_, _04056_, _04053_);
  and (_04058_, _03568_, _03945_);
  not (_04059_, _04058_);
  not (_04061_, _03266_);
  and (_04062_, _03677_, _04061_);
  and (_04063_, _03577_, _03945_);
  nor (_04064_, _04063_, _04062_);
  and (_04065_, _04064_, _04059_);
  nor (_04066_, _03677_, _03523_);
  nor (_04067_, _04066_, _03261_);
  not (_04068_, _04067_);
  not (_04069_, _03966_);
  and (_04070_, _03570_, _03945_);
  nor (_04071_, _04070_, _03599_);
  and (_04072_, _04071_, _04069_);
  and (_04073_, _04072_, _04068_);
  and (_04074_, _04073_, _04065_);
  and (_04075_, _04074_, _04057_);
  or (_04076_, _04075_, _04049_);
  nand (_04077_, _04076_, _03516_);
  nand (_04078_, _03517_, _04077_);
  not (_04079_, \oc8051_golden_model_1.SP [0]);
  and (_04080_, _03597_, _04079_);
  nor (_04081_, _04080_, _03603_);
  and (_04082_, _03677_, _03509_);
  and (_04083_, _03170_, _03134_);
  and (_04084_, _04083_, _03509_);
  nor (_04085_, _04084_, _04082_);
  and (_04086_, _04085_, _04081_);
  nand (_04087_, _04086_, _04078_);
  nand (_04088_, _04087_, _04048_);
  and (_04089_, _04088_, _03512_);
  or (_04090_, _03513_, _04089_);
  and (_04091_, _04042_, _03510_);
  and (_04092_, _03568_, _03503_);
  nor (_04093_, _04092_, _03664_);
  or (_04094_, _03678_, _03615_);
  and (_04095_, _03570_, _03503_);
  nor (_04096_, _04095_, _03662_);
  not (_04097_, _04096_);
  nor (_04098_, _04097_, _04094_);
  and (_04099_, _04098_, _04093_);
  not (_04100_, _04099_);
  nor (_04101_, _04100_, _04091_);
  and (_04102_, _04101_, _04090_);
  or (_04103_, _04102_, _04047_);
  and (_04104_, _04103_, _03622_);
  nor (_04105_, _03622_, _03495_);
  or (_04106_, _04105_, _04104_);
  and (_04107_, _04042_, _03594_);
  and (_04108_, _03677_, _03566_);
  nor (_04109_, _04108_, _03636_);
  not (_04110_, _04109_);
  nor (_04111_, _04110_, _04107_);
  and (_04112_, _04111_, _04106_);
  nor (_04113_, _03631_, _03495_);
  or (_04114_, _04113_, _04112_);
  not (_04115_, _03677_);
  nor (_04116_, _04050_, _03523_);
  and (_04117_, _04116_, _04115_);
  nor (_04118_, _04117_, _03277_);
  and (_04119_, _03568_, _03276_);
  and (_04120_, _03666_, _03276_);
  and (_04121_, _04120_, _03170_);
  nor (_04122_, _04121_, _04119_);
  not (_04123_, _04122_);
  nor (_04124_, _04123_, _04118_);
  and (_04125_, _04124_, _04114_);
  or (_04126_, _04125_, _04045_);
  and (_04127_, _04126_, _03501_);
  or (_04128_, _04127_, _03502_);
  and (_04129_, _03568_, _03219_);
  not (_04130_, _04129_);
  and (_04131_, _03570_, _03219_);
  nor (_04132_, _04131_, _03644_);
  and (_04133_, _04132_, _04130_);
  and (_04134_, _03577_, _03219_);
  not (_04135_, _04134_);
  and (_04136_, _03677_, _03219_);
  nor (_04137_, _04136_, _03970_);
  and (_04138_, _04137_, _04135_);
  and (_04139_, _04138_, _04133_);
  and (_04140_, _04139_, _04128_);
  and (_04141_, _03761_, _01904_);
  and (_04142_, _03716_, _01911_);
  nor (_04143_, _04142_, _04141_);
  and (_04144_, _03748_, _01898_);
  and (_04145_, _03745_, _01945_);
  nor (_04146_, _04145_, _04144_);
  and (_04147_, _04146_, _04143_);
  and (_04148_, _03736_, _01906_);
  and (_04149_, _03743_, _01909_);
  nor (_04150_, _04149_, _04148_);
  and (_04151_, _03759_, _01896_);
  and (_04152_, _03754_, _01933_);
  nor (_04153_, _04152_, _04151_);
  and (_04154_, _04153_, _04150_);
  and (_04155_, _04154_, _04147_);
  and (_04156_, _03732_, _01922_);
  and (_04157_, _03725_, _01927_);
  nor (_04158_, _04157_, _04156_);
  and (_04159_, _03750_, _01942_);
  and (_04160_, _03756_, _01935_);
  nor (_04162_, _04160_, _04159_);
  and (_04163_, _04162_, _04158_);
  and (_04164_, _03712_, _01902_);
  and (_04165_, _03738_, _01930_);
  nor (_04166_, _04165_, _04164_);
  and (_04167_, _03721_, _01917_);
  and (_04168_, _03729_, _01919_);
  nor (_04169_, _04168_, _04167_);
  and (_04170_, _04169_, _04166_);
  and (_04171_, _04170_, _04163_);
  and (_04172_, _04171_, _04155_);
  nor (_04173_, _04172_, _03275_);
  or (_04174_, _04173_, _04140_);
  and (_04175_, _03562_, _03495_);
  and (_04176_, _03677_, _03226_);
  nor (_04177_, _04176_, _03561_);
  not (_04178_, _04177_);
  nor (_04179_, _04178_, _04175_);
  and (_04180_, _04179_, _04174_);
  not (_04181_, _03561_);
  nor (_04182_, _04181_, _03495_);
  or (_04183_, _04182_, _04180_);
  and (_04184_, _03677_, _03230_);
  not (_04185_, _04184_);
  and (_04186_, _04050_, _03230_);
  and (_04187_, _03567_, _03170_);
  and (_04188_, _04187_, _03230_);
  nor (_04189_, _04188_, _04186_);
  and (_04190_, _04189_, _04185_);
  and (_04191_, _04190_, _04183_);
  not (_04192_, _04042_);
  nor (_04193_, _04192_, _03781_);
  not (_04194_, _03237_);
  nor (_04195_, _04051_, _04194_);
  not (_04196_, _04195_);
  nor (_04197_, _03273_, _03202_);
  and (_04198_, _04197_, _03237_);
  and (_04199_, _04198_, _03170_);
  and (_04200_, _03666_, _03237_);
  and (_04201_, _04200_, _03170_);
  nor (_04202_, _04201_, _04199_);
  and (_04203_, _04202_, _04196_);
  not (_04204_, _03235_);
  nor (_04205_, _04051_, _04204_);
  and (_04206_, _03666_, _03235_);
  and (_04207_, _04197_, _03235_);
  or (_04208_, _04207_, _04206_);
  and (_04209_, _04208_, _03170_);
  nor (_04210_, _04209_, _04205_);
  and (_04211_, _04210_, _04203_);
  not (_04212_, _04211_);
  nor (_04213_, _04212_, _04193_);
  and (_04214_, _04213_, _04191_);
  nor (_04215_, _04192_, _03788_);
  and (_04216_, _03568_, _03247_);
  and (_04217_, _03677_, _03247_);
  nor (_04218_, _04217_, _04216_);
  and (_04219_, _03570_, _03247_);
  not (_04220_, _03247_);
  nor (_04221_, _04116_, _04220_);
  nor (_04222_, _04221_, _04219_);
  and (_04223_, _04222_, _04218_);
  not (_04224_, _04223_);
  nor (_04225_, _04224_, _04215_);
  and (_04226_, _04225_, _04214_);
  nor (_04227_, _04042_, _03783_);
  nor (_04228_, _04227_, _04226_);
  and (_04229_, _03792_, _04079_);
  nor (_04230_, _04229_, _04228_);
  and (_04231_, _03652_, _03495_);
  and (_04232_, _03677_, _03245_);
  and (_04233_, _03570_, _03245_);
  nor (_04234_, _04233_, _04232_);
  and (_04235_, _03577_, _03245_);
  and (_04236_, _03568_, _03245_);
  nor (_04237_, _04236_, _04235_);
  and (_04238_, _03587_, _03245_);
  nor (_04239_, _04238_, _03524_);
  and (_04240_, _04239_, _04237_);
  and (_04241_, _04240_, _04234_);
  not (_04242_, _04241_);
  nor (_04243_, _04242_, _04231_);
  and (_04244_, _04243_, _04230_);
  nor (_04245_, _04042_, _03525_);
  nor (_04246_, _04245_, _04244_);
  and (_04247_, _03521_, _04079_);
  nor (_04248_, _04247_, _04246_);
  and (_04249_, _03519_, _03495_);
  and (_04250_, _03570_, _03066_);
  nor (_04251_, _04250_, _03809_);
  not (_04252_, _04251_);
  not (_04253_, _03066_);
  and (_04254_, _04051_, _04115_);
  nor (_04255_, _04254_, _04253_);
  nor (_04256_, _04255_, _04252_);
  not (_04257_, _04256_);
  nor (_04258_, _04257_, _04249_);
  and (_04259_, _04258_, _04248_);
  not (_04260_, _03809_);
  nor (_04261_, _04042_, _04260_);
  or (_04263_, _04261_, _04259_);
  and (_04264_, _04263_, _03206_);
  or (_04265_, _04264_, _03496_);
  and (_04266_, _03568_, _03241_);
  and (_04267_, _04050_, _03241_);
  or (_04268_, _04267_, _03816_);
  or (_04269_, _04268_, _04266_);
  and (_04270_, _03570_, _03241_);
  and (_04271_, _04197_, _03241_);
  and (_04272_, _04271_, _03170_);
  or (_04273_, _04272_, _04270_);
  nor (_04274_, _04273_, _04269_);
  nand (_04275_, _04274_, _04265_);
  and (_04276_, _04275_, _04044_);
  nand (_04277_, _04276_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_04278_, _03420_, _41943_);
  nor (_04279_, _03458_, _41994_);
  nor (_04280_, _04279_, _04278_);
  nor (_04281_, _03433_, _42404_);
  nor (_04282_, _03452_, _42158_);
  nor (_04283_, _04282_, _04281_);
  and (_04284_, _04283_, _04280_);
  nor (_04285_, _03444_, _42035_);
  nor (_04286_, _03428_, _42076_);
  nor (_04287_, _04286_, _04285_);
  nor (_04288_, _03455_, _42363_);
  nor (_04289_, _03412_, _42281_);
  nor (_04290_, _04289_, _04288_);
  and (_04291_, _04290_, _04287_);
  and (_04292_, _04291_, _04284_);
  nor (_04293_, _03406_, _42527_);
  nor (_04294_, _03450_, _42486_);
  nor (_04295_, _04294_, _04293_);
  nor (_04296_, _03431_, _42445_);
  nor (_04297_, _03441_, _42240_);
  nor (_04298_, _04297_, _04296_);
  and (_04299_, _04298_, _04295_);
  nor (_04300_, _03439_, _42322_);
  nor (_04301_, _03446_, _41897_);
  nor (_04302_, _04301_, _04300_);
  nor (_04303_, _03424_, _42199_);
  nor (_04304_, _03417_, _42117_);
  nor (_04305_, _04304_, _04303_);
  and (_04306_, _04305_, _04302_);
  and (_04307_, _04306_, _04299_);
  and (_04308_, _04307_, _04292_);
  nor (_04309_, _04308_, _03463_);
  and (_04310_, _03861_, _03512_);
  and (_04311_, _04310_, _03860_);
  not (_04312_, _04311_);
  and (_04313_, _04312_, _04309_);
  not (_04314_, _04313_);
  and (_04315_, _04309_, _03500_);
  not (_04316_, _04315_);
  and (_04317_, _03725_, _01975_);
  and (_04318_, _03732_, _01998_);
  nor (_04319_, _04318_, _04317_);
  and (_04320_, _03748_, _01954_);
  and (_04321_, _03754_, _01986_);
  nor (_04322_, _04321_, _04320_);
  and (_04323_, _04322_, _04319_);
  and (_04324_, _03721_, _01978_);
  and (_04325_, _03756_, _01991_);
  nor (_04326_, _04325_, _04324_);
  and (_04327_, _03738_, _01989_);
  and (_04328_, _03716_, _01964_);
  nor (_04329_, _04328_, _04327_);
  and (_04330_, _04329_, _04326_);
  and (_04331_, _04330_, _04323_);
  and (_04332_, _03736_, _01961_);
  and (_04333_, _03743_, _01959_);
  nor (_04334_, _04333_, _04332_);
  and (_04335_, _03712_, _01957_);
  and (_04336_, _03759_, _01952_);
  nor (_04337_, _04336_, _04335_);
  and (_04338_, _04337_, _04334_);
  and (_04339_, _03750_, _01983_);
  and (_04340_, _03745_, _02001_);
  nor (_04341_, _04340_, _04339_);
  and (_04342_, _03729_, _01972_);
  and (_04343_, _03761_, _01966_);
  nor (_04344_, _04343_, _04342_);
  and (_04345_, _04344_, _04341_);
  and (_04346_, _04345_, _04338_);
  and (_04347_, _04346_, _04331_);
  nor (_04348_, _04347_, _03275_);
  not (_04349_, _03584_);
  nor (_04350_, _03219_, _03241_);
  and (_04351_, _04350_, _04000_);
  nor (_04352_, _04351_, _04349_);
  not (_04353_, _04352_);
  and (_04354_, _03668_, _03245_);
  not (_04355_, _04354_);
  and (_04356_, _03668_, _03945_);
  and (_04357_, _03668_, _03237_);
  nor (_04358_, _04357_, _04356_);
  and (_04359_, _04358_, _04355_);
  and (_04360_, _04359_, _04353_);
  and (_04361_, _03690_, _03509_);
  nor (_04362_, _04361_, _03953_);
  not (_04364_, _04362_);
  not (_04365_, \oc8051_golden_model_1.SP [1]);
  nor (_04366_, _03597_, _03792_);
  nor (_04367_, _04366_, _04365_);
  nor (_04368_, _04367_, _04364_);
  and (_04369_, _04368_, _04360_);
  not (_04370_, _04001_);
  and (_04371_, _04370_, _03990_);
  and (_04372_, _03521_, \oc8051_golden_model_1.SP [1]);
  nor (_04373_, _04372_, _04266_);
  and (_04374_, _04373_, _04371_);
  and (_04375_, _03668_, _03230_);
  nor (_04376_, _04375_, _03977_);
  and (_04377_, _03668_, _03235_);
  and (_04378_, _03668_, _03509_);
  nor (_04379_, _04378_, _04377_);
  and (_04380_, _04379_, _04376_);
  nor (_04381_, _03669_, _03946_);
  and (_04382_, _04381_, _03984_);
  and (_04383_, _04382_, _04380_);
  and (_04384_, _04383_, _04374_);
  and (_04385_, _03567_, _03066_);
  and (_04386_, _04385_, _03201_);
  not (_04387_, _04386_);
  and (_04388_, _03690_, _03235_);
  and (_04389_, _03690_, _03241_);
  nor (_04390_, _04389_, _04388_);
  and (_04391_, _04390_, _04387_);
  nor (_04392_, _04216_, _04129_);
  not (_04393_, _04119_);
  and (_04394_, _03690_, _03514_);
  and (_04395_, _03668_, _03514_);
  nor (_04396_, _04395_, _04394_);
  and (_04397_, _04396_, _04393_);
  and (_04398_, _04397_, _04392_);
  and (_04399_, _04398_, _04391_);
  and (_04400_, _04399_, _04384_);
  and (_04401_, _04400_, _04369_);
  not (_04402_, _04401_);
  nor (_04403_, _04402_, _04348_);
  nor (_04404_, _03406_, _42512_);
  nor (_04405_, _03420_, _41923_);
  nor (_04406_, _04405_, _04404_);
  nor (_04407_, _03439_, _42307_);
  nor (_04408_, _03446_, _41882_);
  nor (_04409_, _04408_, _04407_);
  and (_04410_, _04409_, _04406_);
  nor (_04411_, _03441_, _42225_);
  nor (_04412_, _03458_, _41971_);
  nor (_04413_, _04412_, _04411_);
  nor (_04414_, _03424_, _42184_);
  nor (_04415_, _03428_, _42061_);
  nor (_04416_, _04415_, _04414_);
  and (_04417_, _04416_, _04413_);
  and (_04418_, _04417_, _04410_);
  nor (_04419_, _03417_, _42102_);
  nor (_04420_, _03444_, _42020_);
  nor (_04421_, _04420_, _04419_);
  nor (_04422_, _03450_, _42471_);
  nor (_04423_, _03455_, _42348_);
  nor (_04424_, _04423_, _04422_);
  and (_04425_, _04424_, _04421_);
  nor (_04426_, _03433_, _42389_);
  nor (_04427_, _03412_, _42266_);
  nor (_04428_, _04427_, _04426_);
  nor (_04429_, _03431_, _42430_);
  nor (_04430_, _03452_, _42143_);
  nor (_04431_, _04430_, _04429_);
  and (_04432_, _04431_, _04428_);
  and (_04433_, _04432_, _04425_);
  and (_04434_, _04433_, _04418_);
  not (_04435_, _04434_);
  and (_04436_, _04435_, _03910_);
  not (_04437_, _04436_);
  and (_04438_, _04437_, _04403_);
  and (_04439_, _04438_, _04316_);
  and (_04440_, _04439_, _04314_);
  nand (_04441_, _04275_, _04044_);
  nand (_04442_, _04441_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_04443_, _04442_, _04440_);
  nand (_04444_, _04443_, _04277_);
  nand (_04445_, _04441_, \oc8051_golden_model_1.IRAM[3] [0]);
  not (_04446_, _04440_);
  nand (_04447_, _04276_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_04448_, _04447_, _04446_);
  nand (_04449_, _04448_, _04445_);
  nand (_04450_, _04449_, _04444_);
  nand (_04451_, _04450_, _04011_);
  not (_04452_, _04011_);
  nand (_04453_, _04441_, \oc8051_golden_model_1.IRAM[7] [0]);
  nand (_04454_, _04276_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_04455_, _04454_, _04446_);
  nand (_04456_, _04455_, _04453_);
  nand (_04457_, _04276_, \oc8051_golden_model_1.IRAM[4] [0]);
  nand (_04458_, _04441_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_04459_, _04458_, _04440_);
  nand (_04460_, _04459_, _04457_);
  nand (_04461_, _04460_, _04456_);
  nand (_04462_, _04461_, _04452_);
  nand (_04463_, _04462_, _04451_);
  nand (_04465_, _04463_, _03822_);
  not (_04466_, _03822_);
  nand (_04467_, _04441_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_04468_, _04276_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_04469_, _04468_, _04446_);
  nand (_04470_, _04469_, _04467_);
  nand (_04471_, _04276_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_04472_, _04441_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_04473_, _04472_, _04440_);
  nand (_04474_, _04473_, _04471_);
  nand (_04475_, _04474_, _04470_);
  nand (_04476_, _04475_, _04011_);
  not (_04477_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_04478_, _04276_, _04477_);
  nand (_04479_, _04276_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_04480_, _04479_, _04446_);
  nand (_04481_, _04480_, _04478_);
  not (_04482_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_04483_, _04441_, _04482_);
  nand (_04484_, _04441_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_04485_, _04484_, _04440_);
  nand (_04486_, _04485_, _04483_);
  nand (_04487_, _04486_, _04481_);
  nand (_04488_, _04487_, _04452_);
  nand (_04489_, _04488_, _04476_);
  nand (_04490_, _04489_, _04466_);
  and (_04491_, _04490_, _04465_);
  and (_04492_, _04491_, _03518_);
  nor (_04493_, _03675_, _03214_);
  nor (_04494_, _03677_, _03570_);
  nand (_04495_, _04494_, _04493_);
  and (_04496_, _04495_, _04061_);
  not (_04497_, _04496_);
  nor (_04498_, _04497_, _04492_);
  and (_04499_, _03582_, _03945_);
  not (_04500_, _04499_);
  nor (_04501_, _04500_, _03463_);
  and (_04502_, _04042_, _04501_);
  or (_04503_, _04502_, _04498_);
  and (_04504_, _03947_, \oc8051_golden_model_1.SP [0]);
  and (_04505_, _04083_, _03514_);
  nor (_04506_, _04505_, _04504_);
  not (_04507_, _04506_);
  nor (_04508_, _04507_, _04503_);
  and (_04509_, _04197_, _03514_);
  nand (_04510_, _04490_, _04465_);
  and (_04511_, _04510_, _04509_);
  not (_04512_, _04511_);
  and (_04513_, _04512_, _04508_);
  nor (_04514_, _03516_, _03463_);
  not (_04515_, _03599_);
  nor (_04516_, _04515_, _03463_);
  and (_04517_, _04516_, _04042_);
  nor (_04518_, _04517_, _04514_);
  and (_04519_, _04518_, _04513_);
  not (_04520_, _04519_);
  and (_04521_, _04520_, _03517_);
  nor (_04522_, _03257_, _04079_);
  nor (_04523_, _04522_, _04521_);
  not (_04524_, _03597_);
  nor (_04525_, _04524_, _03463_);
  and (_04526_, _04525_, _04042_);
  nor (_04527_, _04526_, _04084_);
  and (_04528_, _04527_, _04523_);
  and (_04529_, _04197_, _03509_);
  and (_04530_, _04529_, _04510_);
  not (_04531_, _04530_);
  and (_04532_, _04531_, _04528_);
  nor (_04533_, _03512_, _03463_);
  nor (_04534_, _03611_, _03463_);
  and (_04535_, _04534_, _04042_);
  nor (_04536_, _04535_, _04533_);
  and (_04537_, _04536_, _04532_);
  nor (_04538_, _04537_, _03513_);
  nor (_04539_, _04538_, _03510_);
  and (_04540_, _03510_, _04079_);
  or (_04541_, _04540_, _04539_);
  and (_04542_, _04541_, _03508_);
  nor (_04543_, _04542_, _03506_);
  nor (_04544_, _03253_, _04079_);
  and (_04545_, _04050_, _03566_);
  nor (_04546_, _04545_, _04544_);
  and (_04547_, _04546_, _03572_);
  not (_04548_, _04547_);
  nor (_04549_, _04548_, _04543_);
  nor (_04550_, _03501_, _03463_);
  and (_04551_, _04197_, _03566_);
  and (_04552_, _04551_, _04510_);
  nor (_04553_, _04552_, _04550_);
  and (_04554_, _04553_, _04549_);
  nor (_04555_, _04554_, _03502_);
  nor (_04556_, _04555_, _03497_);
  nor (_04557_, _03278_, \oc8051_golden_model_1.SP [0]);
  nor (_04558_, _04557_, _04556_);
  not (_04559_, _03463_);
  and (_04560_, _03970_, _04559_);
  nor (_04561_, _03463_, _03271_);
  not (_04562_, _03203_);
  and (_04563_, _03574_, _04562_);
  nor (_04564_, _04563_, _03567_);
  not (_04566_, _04564_);
  and (_04567_, _04566_, _04561_);
  nor (_04568_, _04567_, _04560_);
  nor (_04569_, _03463_, _03275_);
  and (_04570_, _04561_, _04197_);
  nor (_04571_, _04570_, _04569_);
  and (_04572_, _04571_, _04568_);
  nor (_04573_, _04572_, _04192_);
  and (_04574_, _04083_, _03226_);
  nor (_04575_, _04574_, _04573_);
  not (_04576_, _04575_);
  nor (_04577_, _04576_, _04558_);
  and (_04578_, _04197_, _03226_);
  and (_04579_, _04578_, _04510_);
  not (_04580_, _04579_);
  and (_04581_, _04580_, _04577_);
  not (_04582_, _03650_);
  nor (_04583_, _04582_, _03463_);
  and (_04584_, _04583_, _04042_);
  nor (_04585_, _04584_, _03227_);
  and (_04586_, _04585_, _04581_);
  and (_04587_, _03227_, _04079_);
  nor (_04588_, _04587_, _04586_);
  not (_04589_, _03778_);
  nor (_04590_, _04589_, _03463_);
  not (_04591_, _03649_);
  nor (_04592_, _04591_, _03463_);
  nor (_04593_, _04592_, _04590_);
  not (_04594_, _03773_);
  nor (_04595_, _04594_, _03463_);
  not (_04596_, _03655_);
  nor (_04597_, _04596_, _03463_);
  nor (_04598_, _04597_, _04595_);
  and (_04599_, _04598_, _04593_);
  nor (_04600_, _04599_, _04192_);
  nor (_04601_, _04600_, _03238_);
  not (_04602_, _04601_);
  nor (_04603_, _04602_, _04588_);
  and (_04604_, _03238_, _04079_);
  nor (_04605_, _04604_, _04603_);
  not (_04606_, _03786_);
  nor (_04607_, _04606_, _03463_);
  not (_04608_, _03653_);
  nor (_04609_, _04608_, _03463_);
  nor (_04610_, _04609_, _04607_);
  nor (_04611_, _04610_, _04192_);
  nor (_04612_, _04611_, _04605_);
  and (_04613_, _03248_, \oc8051_golden_model_1.SP [0]);
  and (_04614_, _04083_, _03066_);
  nor (_04615_, _04614_, _04613_);
  and (_04616_, _04615_, _04612_);
  nor (_04617_, _04260_, _03463_);
  and (_04618_, _04197_, _03066_);
  and (_04619_, _04618_, _04510_);
  nor (_04620_, _04619_, _04617_);
  and (_04621_, _04620_, _04616_);
  and (_04622_, _04617_, _04192_);
  nor (_04623_, _04622_, _04621_);
  nor (_04624_, _03463_, _03206_);
  nor (_04625_, _03686_, _03243_);
  nor (_04626_, _04625_, _04079_);
  nor (_04627_, _04626_, _04624_);
  not (_04628_, _04627_);
  nor (_04629_, _04628_, _04623_);
  nor (_04630_, _04629_, _03496_);
  and (_04631_, _04083_, _03241_);
  nor (_04632_, _04631_, _04630_);
  nor (_04633_, _03820_, _03463_);
  and (_04634_, _04510_, _04271_);
  nor (_04635_, _04634_, _04633_);
  and (_04636_, _04635_, _04632_);
  and (_04637_, _04633_, _04192_);
  nor (_04638_, _04637_, _04636_);
  not (_04639_, _04638_);
  and (_04640_, _04633_, _04435_);
  and (_04641_, _03949_, _03241_);
  and (_04642_, _03666_, _03241_);
  and (_04643_, _04309_, _03205_);
  and (_04644_, _04365_, \oc8051_golden_model_1.SP [0]);
  and (_04645_, \oc8051_golden_model_1.SP [1], _04079_);
  nor (_04646_, _04645_, _04644_);
  not (_04647_, _04646_);
  and (_04648_, _04647_, _03248_);
  and (_04649_, _04647_, _03510_);
  not (_04650_, _03510_);
  and (_04651_, _04525_, _04435_);
  or (_04652_, _04197_, _03214_);
  and (_04653_, _04652_, _04061_);
  nand (_04654_, _04276_, \oc8051_golden_model_1.IRAM[0] [1]);
  nand (_04655_, _04441_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_04656_, _04655_, _04440_);
  nand (_04657_, _04656_, _04654_);
  nand (_04658_, _04441_, \oc8051_golden_model_1.IRAM[3] [1]);
  nand (_04659_, _04276_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_04660_, _04659_, _04446_);
  nand (_04661_, _04660_, _04658_);
  nand (_04662_, _04661_, _04657_);
  nand (_04663_, _04662_, _04011_);
  nand (_04664_, _04441_, \oc8051_golden_model_1.IRAM[7] [1]);
  nand (_04665_, _04276_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_04667_, _04665_, _04446_);
  nand (_04668_, _04667_, _04664_);
  nand (_04669_, _04276_, \oc8051_golden_model_1.IRAM[4] [1]);
  nand (_04670_, _04441_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_04671_, _04670_, _04440_);
  nand (_04672_, _04671_, _04669_);
  nand (_04673_, _04672_, _04668_);
  nand (_04674_, _04673_, _04452_);
  nand (_04675_, _04674_, _04663_);
  nand (_04676_, _04675_, _03822_);
  nand (_04677_, _04441_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_04678_, _04276_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_04679_, _04678_, _04446_);
  nand (_04680_, _04679_, _04677_);
  nand (_04681_, _04276_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_04682_, _04441_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_04683_, _04682_, _04440_);
  nand (_04684_, _04683_, _04681_);
  nand (_04685_, _04684_, _04680_);
  nand (_04686_, _04685_, _04011_);
  nand (_04687_, _04441_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_04688_, _04276_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_04689_, _04688_, _04446_);
  nand (_04690_, _04689_, _04687_);
  nand (_04691_, _04276_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_04692_, _04441_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_04693_, _04692_, _04440_);
  nand (_04694_, _04693_, _04691_);
  nand (_04695_, _04694_, _04690_);
  nand (_04696_, _04695_, _04452_);
  nand (_04697_, _04696_, _04686_);
  nand (_04698_, _04697_, _04466_);
  nand (_04699_, _04698_, _04676_);
  or (_04700_, _04699_, _03213_);
  and (_04701_, _04700_, _04653_);
  and (_04702_, _04434_, _04501_);
  nor (_04703_, _04702_, _04701_);
  and (_04704_, _03949_, _03514_);
  and (_04705_, _03666_, _03514_);
  nor (_04706_, _04705_, _04704_);
  not (_04707_, _04706_);
  and (_04708_, _04646_, _03947_);
  nor (_04709_, _04708_, _04707_);
  and (_04710_, _04709_, _04703_);
  and (_04711_, _04699_, _04509_);
  nor (_04712_, _04711_, _04516_);
  and (_04713_, _04712_, _04710_);
  and (_04714_, _04516_, _04435_);
  nor (_04715_, _04714_, _04713_);
  and (_04716_, _04308_, _04514_);
  nor (_04717_, _04716_, _04715_);
  nor (_04718_, _04647_, _03257_);
  nor (_04719_, _04718_, _04525_);
  and (_04720_, _04719_, _04717_);
  nor (_04721_, _04720_, _04651_);
  and (_04722_, _03949_, _03509_);
  and (_04723_, _03666_, _03509_);
  nor (_04724_, _04723_, _04722_);
  not (_04725_, _04724_);
  nor (_04726_, _04725_, _04721_);
  and (_04727_, _04699_, _04529_);
  nor (_04728_, _04727_, _04534_);
  and (_04729_, _04728_, _04726_);
  and (_04730_, _04534_, _04435_);
  nor (_04731_, _04730_, _04729_);
  and (_04732_, _04308_, _04533_);
  nor (_04733_, _04732_, _04731_);
  and (_04734_, _04733_, _04650_);
  nor (_04735_, _04734_, _04649_);
  and (_04736_, _03507_, _04308_);
  or (_04737_, _04736_, _04735_);
  and (_04738_, _03666_, _03566_);
  and (_04739_, _04738_, _03689_);
  or (_04740_, _04739_, _03588_);
  and (_04741_, _04738_, _03170_);
  nor (_04742_, _04647_, _03253_);
  or (_04743_, _04742_, _04741_);
  or (_04744_, _04743_, _03576_);
  nor (_04745_, _04744_, _04740_);
  not (_04746_, _04745_);
  nor (_04747_, _04746_, _04737_);
  and (_04748_, _04699_, _04551_);
  nor (_04749_, _04748_, _04550_);
  and (_04750_, _04749_, _04747_);
  nor (_04751_, _04750_, _04315_);
  nor (_04752_, _04751_, _03497_);
  nor (_04753_, _04646_, _03278_);
  nor (_04754_, _04753_, _04752_);
  nor (_04755_, _04572_, _04435_);
  and (_04756_, _03226_, _03202_);
  and (_04757_, _04756_, _03134_);
  nor (_04758_, _04757_, _04755_);
  not (_04759_, _04758_);
  nor (_04760_, _04759_, _04754_);
  and (_04761_, _04699_, _04578_);
  nor (_04762_, _04761_, _04583_);
  and (_04763_, _04762_, _04760_);
  and (_04764_, _04583_, _04435_);
  nor (_04765_, _04764_, _04763_);
  nor (_04766_, _04765_, _03227_);
  and (_04768_, _04647_, _03227_);
  nor (_04769_, _04768_, _04766_);
  nor (_04770_, _04599_, _04435_);
  nor (_04771_, _04770_, _03238_);
  not (_04772_, _04771_);
  nor (_04773_, _04772_, _04769_);
  and (_04774_, _04647_, _03238_);
  nor (_04775_, _04774_, _04773_);
  nor (_04776_, _03787_, _03463_);
  and (_04777_, _04776_, _04434_);
  or (_04778_, _04777_, _03248_);
  nor (_04779_, _04778_, _04775_);
  nor (_04780_, _04779_, _04648_);
  and (_04781_, _03666_, _03066_);
  nor (_04782_, _04781_, _03975_);
  not (_04783_, _04782_);
  nor (_04784_, _04783_, _04780_);
  and (_04785_, _04699_, _04618_);
  nor (_04786_, _04785_, _04617_);
  and (_04787_, _04786_, _04784_);
  and (_04788_, _04617_, _04435_);
  nor (_04789_, _04788_, _04787_);
  nor (_04790_, _04647_, _04625_);
  nor (_04791_, _04790_, _04624_);
  not (_04792_, _04791_);
  nor (_04793_, _04792_, _04789_);
  nor (_04794_, _04793_, _04643_);
  or (_04795_, _04794_, _04642_);
  nor (_04796_, _04795_, _04641_);
  and (_04797_, _04699_, _04271_);
  nor (_04798_, _04797_, _04633_);
  and (_04799_, _04798_, _04796_);
  nor (_04800_, _04799_, _04640_);
  not (_04801_, _00000_);
  nor (_04802_, _04590_, _04595_);
  nor (_04803_, _04592_, _04597_);
  and (_04804_, _04803_, _04802_);
  not (_04805_, _04633_);
  nor (_04806_, _04560_, _04624_);
  and (_04807_, _04806_, _04805_);
  and (_04808_, _04807_, _04804_);
  and (_04809_, _04808_, _04571_);
  not (_04810_, _04567_);
  not (_04811_, _04617_);
  and (_04812_, _03575_, _03241_);
  not (_04813_, _03226_);
  nor (_04814_, _04197_, _03666_);
  or (_04815_, _04814_, _04813_);
  not (_04816_, _04815_);
  nor (_04817_, _04816_, _04812_);
  and (_04818_, _03589_, _03509_);
  nor (_04819_, _04818_, _04378_);
  and (_04820_, _04819_, _04706_);
  nor (_04821_, _04814_, _03266_);
  and (_04822_, _03567_, _03226_);
  and (_04823_, _04822_, _03498_);
  nor (_04824_, _04823_, _04821_);
  and (_04825_, _04824_, _04820_);
  nor (_04826_, _04389_, _04386_);
  nor (_04827_, _04814_, _04253_);
  and (_04828_, _04822_, _03581_);
  nor (_04829_, _04828_, _04827_);
  and (_04830_, _04829_, _04826_);
  and (_04831_, _04830_, _04825_);
  and (_04832_, _04831_, _04817_);
  and (_04833_, _04493_, _03274_);
  nor (_04834_, _04833_, _03266_);
  not (_04835_, _04834_);
  and (_04836_, _03668_, _03566_);
  nor (_04837_, _04836_, _03590_);
  not (_04838_, _03241_);
  nor (_04839_, _03587_, _03668_);
  nor (_04840_, _04839_, _04838_);
  not (_04841_, _04840_);
  and (_04842_, _04841_, _04837_);
  and (_04843_, _04842_, _04835_);
  and (_04844_, _03582_, _03226_);
  and (_04845_, _03574_, _03283_);
  and (_04846_, _04845_, _03566_);
  nor (_04847_, _04846_, _04844_);
  and (_04848_, _03570_, _03509_);
  and (_04849_, _04845_, _03226_);
  nor (_04850_, _04849_, _04848_);
  and (_04851_, _04850_, _04847_);
  nor (_04852_, _04642_, _04509_);
  nor (_04853_, _04551_, _04529_);
  and (_04854_, _04853_, _04852_);
  and (_04855_, _04854_, _04851_);
  and (_04856_, _03278_, _03253_);
  not (_04857_, _03257_);
  nor (_04858_, _04857_, _03227_);
  and (_04859_, _04858_, _04856_);
  and (_04860_, _04859_, _04362_);
  and (_04861_, _04860_, _04855_);
  nor (_04862_, _03238_, _03248_);
  not (_04863_, _04862_);
  nor (_04864_, _04741_, _04863_);
  not (_04865_, _04722_);
  and (_04866_, _04396_, _04865_);
  and (_04867_, _04866_, _04864_);
  not (_04868_, _03947_);
  and (_04869_, _04625_, _04868_);
  nor (_04870_, _04271_, _03510_);
  nor (_04871_, _03975_, _03583_);
  and (_04872_, _04871_, _04870_);
  and (_04873_, _04872_, _04869_);
  and (_04874_, _04873_, _04867_);
  and (_04875_, _04874_, _04861_);
  and (_04876_, _04875_, _04843_);
  and (_04877_, _04876_, _04832_);
  and (_04878_, _04877_, _04811_);
  nor (_04879_, _04776_, _04583_);
  and (_04880_, _04879_, _04878_);
  and (_04881_, _04880_, _04810_);
  nor (_04882_, _03507_, _04550_);
  nor (_04883_, _04514_, _04501_);
  and (_04884_, _04883_, _04882_);
  nor (_04885_, _04534_, _04533_);
  nor (_04886_, _04525_, _04516_);
  and (_04887_, _04886_, _04885_);
  and (_04888_, _04887_, _04884_);
  and (_04889_, _04888_, _04881_);
  and (_04890_, _04889_, _04809_);
  nor (_04891_, _04890_, _04801_);
  not (_04892_, _04891_);
  nor (_04893_, _04892_, _04800_);
  and (_04894_, _04893_, _04639_);
  and (_04895_, _03821_, _04559_);
  nand (_04896_, _04276_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand (_04897_, _04441_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_04898_, _04897_, _04440_);
  nand (_04899_, _04898_, _04896_);
  nand (_04900_, _04441_, \oc8051_golden_model_1.IRAM[3] [3]);
  not (_04901_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_04902_, _04441_, _04901_);
  and (_04903_, _04902_, _04446_);
  nand (_04904_, _04903_, _04900_);
  nand (_04905_, _04904_, _04899_);
  nand (_04906_, _04905_, _04011_);
  nand (_04907_, _04441_, \oc8051_golden_model_1.IRAM[7] [3]);
  nand (_04908_, _04276_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_04909_, _04908_, _04446_);
  nand (_04910_, _04909_, _04907_);
  nand (_04911_, _04276_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand (_04912_, _04441_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_04913_, _04912_, _04440_);
  nand (_04914_, _04913_, _04911_);
  nand (_04915_, _04914_, _04910_);
  nand (_04916_, _04915_, _04452_);
  nand (_04917_, _04916_, _04906_);
  nand (_04918_, _04917_, _03822_);
  nand (_04919_, _04441_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_04920_, _04276_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_04921_, _04920_, _04446_);
  nand (_04922_, _04921_, _04919_);
  nand (_04923_, _04276_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_04924_, _04441_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_04925_, _04924_, _04440_);
  nand (_04926_, _04925_, _04923_);
  nand (_04927_, _04926_, _04922_);
  nand (_04928_, _04927_, _04011_);
  not (_04929_, \oc8051_golden_model_1.IRAM[15] [3]);
  or (_04930_, _04276_, _04929_);
  not (_04931_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_04932_, _04441_, _04931_);
  and (_04933_, _04932_, _04446_);
  nand (_04934_, _04933_, _04930_);
  nand (_04935_, _04276_, \oc8051_golden_model_1.IRAM[12] [3]);
  not (_04936_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_04937_, _04276_, _04936_);
  and (_04938_, _04937_, _04440_);
  nand (_04939_, _04938_, _04935_);
  nand (_04940_, _04939_, _04934_);
  nand (_04941_, _04940_, _04452_);
  nand (_04942_, _04941_, _04928_);
  nand (_04943_, _04942_, _04466_);
  nand (_04944_, _04943_, _04918_);
  and (_04945_, _04944_, _04578_);
  and (_04946_, _04514_, _03556_);
  and (_04947_, _04944_, _04509_);
  and (_04948_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04949_, _04948_, \oc8051_golden_model_1.SP [2]);
  nor (_04950_, _04949_, \oc8051_golden_model_1.SP [3]);
  and (_04951_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04952_, _04951_, \oc8051_golden_model_1.SP [3]);
  and (_04953_, _04952_, \oc8051_golden_model_1.SP [0]);
  nor (_04954_, _04953_, _04950_);
  and (_04955_, _04954_, _03947_);
  and (_04956_, _04944_, _03518_);
  not (_04957_, \oc8051_golden_model_1.PSW [3]);
  and (_04958_, _03267_, _04957_);
  nor (_04959_, _04958_, _04956_);
  nor (_04960_, _04959_, _04501_);
  and (_04961_, _04501_, _03494_);
  nor (_04962_, _04961_, _03947_);
  not (_04963_, _04962_);
  nor (_04964_, _04963_, _04960_);
  or (_04965_, _04964_, _04509_);
  nor (_04966_, _04965_, _04955_);
  or (_04967_, _04966_, _04516_);
  nor (_04968_, _04967_, _04947_);
  and (_04969_, _04516_, _03558_);
  or (_04970_, _04969_, _04514_);
  nor (_04971_, _04970_, _04968_);
  nor (_04972_, _04971_, _04946_);
  nor (_04973_, _04972_, _04857_);
  nor (_04974_, _04954_, _03257_);
  nor (_04975_, _04974_, _04525_);
  not (_04976_, _04975_);
  nor (_04977_, _04976_, _04973_);
  and (_04978_, _04525_, _03558_);
  nor (_04979_, _04978_, _04529_);
  not (_04980_, _04979_);
  nor (_04981_, _04980_, _04977_);
  and (_04982_, _04944_, _04529_);
  nor (_04983_, _04982_, _04534_);
  not (_04984_, _04983_);
  nor (_04985_, _04984_, _04981_);
  and (_04986_, _04534_, _03558_);
  or (_04987_, _04986_, _04533_);
  nor (_04988_, _04987_, _04985_);
  and (_04989_, _03556_, _04533_);
  nor (_04990_, _04989_, _04988_);
  and (_04991_, _04990_, _04650_);
  and (_04992_, _04954_, _03510_);
  nor (_04993_, _04992_, _04991_);
  nor (_04994_, _04993_, _03507_);
  nor (_04995_, _03508_, _03560_);
  or (_04996_, _04995_, _04994_);
  and (_04997_, _04996_, _03253_);
  not (_04998_, _03253_);
  nor (_04999_, _04551_, _04998_);
  nor (_05000_, _04954_, _04551_);
  nor (_05001_, _05000_, _04999_);
  nor (_05002_, _05001_, _04997_);
  and (_05003_, _04944_, _04551_);
  nor (_05004_, _05003_, _04550_);
  not (_05005_, _05004_);
  nor (_05006_, _05005_, _05002_);
  not (_05007_, _04550_);
  nor (_05008_, _05007_, _03560_);
  nor (_05009_, _05008_, _05006_);
  nor (_05010_, _05009_, _03497_);
  and (_05011_, _04954_, _03497_);
  not (_05012_, _05011_);
  and (_05013_, _05012_, _04572_);
  not (_05014_, _05013_);
  nor (_05015_, _05014_, _05010_);
  nor (_05016_, _04572_, _03558_);
  nor (_05017_, _05016_, _05015_);
  nor (_05018_, _05017_, _04578_);
  or (_05019_, _05018_, _04583_);
  nor (_05020_, _05019_, _04945_);
  and (_05021_, _04583_, _03558_);
  nor (_05022_, _05021_, _05020_);
  nor (_05023_, _05022_, _03227_);
  and (_05024_, _04954_, _03227_);
  not (_05025_, _05024_);
  and (_05026_, _05025_, _04804_);
  not (_05027_, _05026_);
  nor (_05028_, _05027_, _05023_);
  nor (_05029_, _04599_, _03558_);
  nor (_05030_, _05029_, _03238_);
  not (_05031_, _05030_);
  nor (_05032_, _05031_, _05028_);
  and (_05033_, _04954_, _03238_);
  or (_05034_, _05033_, _04776_);
  nor (_05035_, _05034_, _05032_);
  and (_05036_, _04776_, _03494_);
  or (_05037_, _05036_, _03248_);
  nor (_05038_, _05037_, _05035_);
  and (_05039_, _04954_, _03248_);
  nor (_05040_, _05039_, _04618_);
  not (_05041_, _05040_);
  nor (_05042_, _05041_, _05038_);
  and (_05043_, _04944_, _04618_);
  nor (_05044_, _05043_, _04617_);
  not (_05045_, _05044_);
  nor (_05046_, _05045_, _05042_);
  not (_05047_, _04625_);
  and (_05048_, _04617_, _03558_);
  nor (_05049_, _05048_, _05047_);
  not (_05050_, _05049_);
  nor (_05051_, _05050_, _05046_);
  nor (_05052_, _04954_, _04625_);
  nor (_05053_, _05052_, _04624_);
  not (_05054_, _05053_);
  nor (_05055_, _05054_, _05051_);
  not (_05056_, _03556_);
  and (_05057_, _04624_, _05056_);
  nor (_05058_, _05057_, _04271_);
  not (_05059_, _05058_);
  nor (_05060_, _05059_, _05055_);
  and (_05061_, _04944_, _04271_);
  nor (_05062_, _05061_, _04633_);
  not (_05063_, _05062_);
  nor (_05064_, _05063_, _05060_);
  nor (_05065_, _05064_, _04895_);
  and (_05066_, _03854_, _03205_);
  nor (_05067_, _04948_, \oc8051_golden_model_1.SP [2]);
  nor (_05068_, _05067_, _04949_);
  and (_05069_, _05068_, _03248_);
  nor (_05070_, _04572_, _03899_);
  and (_05071_, _03854_, _03500_);
  nor (_05072_, _05068_, _03253_);
  and (_05073_, _03567_, _03566_);
  nor (_05074_, _05073_, _05072_);
  and (_05075_, _04534_, _03899_);
  not (_05076_, _05068_);
  and (_05077_, _05076_, _03947_);
  not (_05078_, _05077_);
  and (_05079_, _03584_, _03514_);
  nor (_05080_, _03589_, _03568_);
  nor (_05081_, _05080_, _03255_);
  or (_05082_, _05081_, _05079_);
  nor (_05083_, _05082_, _04055_);
  and (_05084_, _05083_, _05078_);
  and (_05085_, _03898_, _04501_);
  nand (_05086_, _04276_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand (_05087_, _04441_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_05088_, _05087_, _04440_);
  nand (_05089_, _05088_, _05086_);
  nand (_05090_, _04441_, \oc8051_golden_model_1.IRAM[3] [2]);
  nand (_05091_, _04276_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_05092_, _05091_, _04446_);
  nand (_05093_, _05092_, _05090_);
  nand (_05094_, _05093_, _05089_);
  nand (_05095_, _05094_, _04011_);
  nand (_05096_, _04441_, \oc8051_golden_model_1.IRAM[7] [2]);
  nand (_05097_, _04276_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_05098_, _05097_, _04446_);
  nand (_05099_, _05098_, _05096_);
  nand (_05100_, _04276_, \oc8051_golden_model_1.IRAM[4] [2]);
  nand (_05101_, _04441_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_05102_, _05101_, _04440_);
  nand (_05103_, _05102_, _05100_);
  nand (_05104_, _05103_, _05099_);
  nand (_05105_, _05104_, _04452_);
  nand (_05106_, _05105_, _05095_);
  nand (_05107_, _05106_, _03822_);
  nand (_05108_, _04441_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_05109_, _04276_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_05110_, _05109_, _04446_);
  nand (_05111_, _05110_, _05108_);
  nand (_05112_, _04276_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_05113_, _04441_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_05114_, _05113_, _04440_);
  nand (_05115_, _05114_, _05112_);
  nand (_05116_, _05115_, _05111_);
  nand (_05117_, _05116_, _04011_);
  nand (_05118_, _04441_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_05119_, _04276_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_05120_, _05119_, _04446_);
  nand (_05121_, _05120_, _05118_);
  nand (_05122_, _04276_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_05123_, _04441_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_05124_, _05123_, _04440_);
  nand (_05125_, _05124_, _05122_);
  nand (_05126_, _05125_, _05121_);
  nand (_05127_, _05126_, _04452_);
  nand (_05128_, _05127_, _05117_);
  nand (_05129_, _05128_, _04466_);
  nand (_05130_, _05129_, _05107_);
  nor (_05131_, _05130_, _03213_);
  nor (_05132_, _05131_, _04835_);
  nor (_05133_, _05132_, _05085_);
  and (_05134_, _05133_, _05084_);
  and (_05135_, _05130_, _04509_);
  nor (_05136_, _05135_, _04516_);
  and (_05137_, _05136_, _05134_);
  and (_05138_, _04516_, _03899_);
  nor (_05139_, _05138_, _05137_);
  and (_05140_, _04514_, _03853_);
  nor (_05141_, _05140_, _05139_);
  nor (_05142_, _05068_, _03257_);
  nor (_05143_, _05142_, _04525_);
  and (_05144_, _05143_, _05141_);
  and (_05145_, _04525_, _03899_);
  nor (_05146_, _05145_, _05144_);
  and (_05147_, _03567_, _03509_);
  nor (_05148_, _05147_, _05146_);
  and (_05149_, _05130_, _04529_);
  nor (_05150_, _05149_, _04534_);
  and (_05151_, _05150_, _05148_);
  nor (_05152_, _05151_, _05075_);
  nor (_05153_, _05152_, _04533_);
  nor (_05154_, _05153_, _03866_);
  nor (_05155_, _05154_, _03510_);
  and (_05156_, _05068_, _03510_);
  nor (_05157_, _05156_, _05155_);
  and (_05158_, _03507_, _03853_);
  nor (_05159_, _05158_, _05157_);
  and (_05160_, _05159_, _05074_);
  and (_05161_, _05130_, _04551_);
  nor (_05162_, _05161_, _04550_);
  and (_05163_, _05162_, _05160_);
  nor (_05164_, _05163_, _05071_);
  nor (_05165_, _05164_, _03497_);
  nor (_05166_, _05076_, _03278_);
  nor (_05167_, _05166_, _05165_);
  or (_05168_, _05167_, _04822_);
  nor (_05169_, _05168_, _05070_);
  and (_05170_, _05130_, _04578_);
  nor (_05171_, _05170_, _04583_);
  and (_05172_, _05171_, _05169_);
  and (_05173_, _04583_, _03899_);
  nor (_05174_, _05173_, _05172_);
  nor (_05175_, _05174_, _03227_);
  and (_05176_, _05068_, _03227_);
  nor (_05177_, _05176_, _05175_);
  nor (_05178_, _04599_, _03899_);
  nor (_05179_, _05178_, _03238_);
  not (_05180_, _05179_);
  nor (_05181_, _05180_, _05177_);
  and (_05182_, _05068_, _03238_);
  nor (_05183_, _05182_, _05181_);
  and (_05184_, _04776_, _03898_);
  or (_05185_, _05184_, _03248_);
  nor (_05186_, _05185_, _05183_);
  nor (_05187_, _05186_, _05069_);
  nor (_05188_, _05187_, _04385_);
  and (_05189_, _05130_, _04618_);
  nor (_05190_, _05189_, _04617_);
  and (_05191_, _05190_, _05188_);
  and (_05192_, _04617_, _03899_);
  nor (_05193_, _05192_, _05191_);
  nor (_05194_, _05068_, _04625_);
  nor (_05195_, _05194_, _04624_);
  not (_05196_, _05195_);
  nor (_05197_, _05196_, _05193_);
  nor (_05198_, _05197_, _05066_);
  and (_05199_, _03567_, _03241_);
  nor (_05200_, _05199_, _05198_);
  and (_05201_, _05130_, _04271_);
  nor (_05202_, _05201_, _04633_);
  and (_05203_, _05202_, _05200_);
  and (_05204_, _04633_, _03899_);
  nor (_05205_, _05204_, _05203_);
  nor (_05206_, _05205_, _04892_);
  not (_05207_, _05206_);
  nor (_05208_, _05207_, _05065_);
  and (_05209_, _05208_, _04894_);
  or (_05210_, _05209_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_05211_, _04951_, _04079_);
  nor (_05212_, _05068_, _04645_);
  nor (_05213_, _05212_, _05211_);
  and (_05214_, _04952_, _04079_);
  nor (_05215_, _05211_, _04954_);
  nor (_05216_, _05215_, _05214_);
  and (_05217_, _44104_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_05218_, _05217_);
  and (_05219_, _04869_, _04862_);
  and (_05220_, _05219_, _04859_);
  nor (_05221_, _05220_, _05218_);
  and (_05222_, _05221_, _05216_);
  and (_05223_, _05222_, _05213_);
  and (_05224_, _05223_, _04644_);
  not (_05225_, _05224_);
  and (_05226_, _05225_, _05210_);
  nor (_05227_, _05218_, _04890_);
  not (_05228_, _05227_);
  nor (_05229_, _05228_, _04638_);
  not (_05230_, _05229_);
  nor (_05231_, _05230_, _04800_);
  not (_05232_, _05205_);
  nor (_05233_, _05228_, _05065_);
  and (_05234_, _05233_, _05232_);
  and (_05235_, _05234_, _05231_);
  not (_05236_, _05235_);
  not (_05237_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_05238_, _04441_, _05237_);
  not (_05239_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_05240_, _04276_, _05239_);
  and (_05241_, _05240_, _04440_);
  nand (_05242_, _05241_, _05238_);
  not (_05243_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_05244_, _04276_, _05243_);
  not (_05245_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_05246_, _04441_, _05245_);
  and (_05247_, _05246_, _04446_);
  nand (_05248_, _05247_, _05244_);
  nand (_05249_, _05248_, _05242_);
  nand (_05250_, _05249_, _04011_);
  not (_05251_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_05252_, _04276_, _05251_);
  not (_05253_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_05254_, _04441_, _05253_);
  and (_05255_, _05254_, _04446_);
  nand (_05256_, _05255_, _05252_);
  not (_05257_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_05258_, _04441_, _05257_);
  not (_05259_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_05260_, _04276_, _05259_);
  and (_05261_, _05260_, _04440_);
  nand (_05262_, _05261_, _05258_);
  nand (_05263_, _05262_, _05256_);
  nand (_05264_, _05263_, _04452_);
  nand (_05265_, _05264_, _05250_);
  nand (_05266_, _05265_, _03822_);
  nand (_05267_, _04441_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_05268_, _04276_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_05269_, _05268_, _04446_);
  nand (_05270_, _05269_, _05267_);
  nand (_05271_, _04276_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_05272_, _04441_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_05273_, _05272_, _04440_);
  nand (_05274_, _05273_, _05271_);
  nand (_05275_, _05274_, _05270_);
  nand (_05276_, _05275_, _04011_);
  nand (_05277_, _04441_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_05278_, _04276_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_05279_, _05278_, _04446_);
  nand (_05280_, _05279_, _05277_);
  nand (_05281_, _04276_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_05282_, _04441_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_05283_, _05282_, _04440_);
  nand (_05284_, _05283_, _05281_);
  nand (_05285_, _05284_, _05280_);
  nand (_05286_, _05285_, _04452_);
  nand (_05287_, _05286_, _05276_);
  nand (_05288_, _05287_, _04466_);
  nand (_05289_, _05288_, _05266_);
  or (_05290_, _05289_, _03463_);
  and (_05291_, _03556_, _03463_);
  and (_05292_, _05291_, _03853_);
  and (_05293_, _05292_, _04308_);
  and (_05294_, _05293_, _03494_);
  nor (_05295_, _04434_, _04042_);
  and (_05296_, _05295_, _03898_);
  and (_05297_, _05296_, _05294_);
  and (_05298_, _05297_, \oc8051_golden_model_1.DPH [7]);
  not (_05299_, _05298_);
  not (_05300_, _05293_);
  and (_05301_, _04434_, _04042_);
  nor (_05302_, _03898_, _03494_);
  nand (_05303_, _05302_, _05301_);
  nor (_05304_, _05303_, _05300_);
  and (_05305_, _05304_, \oc8051_golden_model_1.TH0 [7]);
  not (_05306_, _05295_);
  nand (_05307_, _03898_, _03558_);
  or (_05308_, _05307_, _05306_);
  nor (_05309_, _05308_, _05300_);
  and (_05310_, _05309_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05311_, _05310_, _05305_);
  and (_05312_, _05311_, _05299_);
  and (_05313_, _04434_, _04192_);
  and (_05314_, _05313_, _03898_);
  and (_05315_, _05314_, _05294_);
  and (_05316_, _05315_, \oc8051_golden_model_1.SP [7]);
  nor (_05317_, _04434_, _04192_);
  and (_05318_, _05317_, _03898_);
  and (_05319_, _05318_, _05294_);
  and (_05320_, _05319_, \oc8051_golden_model_1.DPL [7]);
  nor (_05321_, _05320_, _05316_);
  and (_05322_, _05295_, _03899_);
  and (_05323_, _05322_, _05294_);
  and (_05324_, _05323_, \oc8051_golden_model_1.PCON [7]);
  not (_05325_, _05324_);
  and (_05326_, _05314_, _03558_);
  not (_05327_, _04308_);
  and (_05328_, _05327_, _03853_);
  and (_05329_, _05328_, _05291_);
  and (_05330_, _05329_, _05326_);
  and (_05331_, _05330_, \oc8051_golden_model_1.SBUF [7]);
  and (_05332_, _05301_, _03898_);
  and (_05333_, _05332_, _03558_);
  not (_05334_, _03853_);
  and (_05335_, _04308_, _05334_);
  and (_05336_, _05335_, _05291_);
  and (_05337_, _05336_, _05333_);
  and (_05338_, _05337_, \oc8051_golden_model_1.IE [7]);
  nor (_05339_, _05338_, _05331_);
  and (_05340_, _05339_, _05325_);
  and (_05341_, _05340_, _05321_);
  and (_05342_, _05341_, _05312_);
  and (_05343_, _05326_, _05293_);
  and (_05344_, _05343_, \oc8051_golden_model_1.TMOD [7]);
  and (_05345_, _05333_, _05329_);
  and (_05346_, _05345_, \oc8051_golden_model_1.SCON [7]);
  nor (_05347_, _05346_, _05344_);
  not (_05348_, _05317_);
  or (_05349_, _05348_, _05307_);
  nor (_05350_, _05349_, _05300_);
  and (_05351_, _05350_, \oc8051_golden_model_1.TL0 [7]);
  not (_05352_, _05351_);
  and (_05353_, _05333_, _05293_);
  and (_05354_, _05353_, \oc8051_golden_model_1.TCON [7]);
  nand (_05355_, _05313_, _05302_);
  nor (_05356_, _05355_, _05300_);
  and (_05357_, _05356_, \oc8051_golden_model_1.TH1 [7]);
  nor (_05358_, _05357_, _05354_);
  and (_05359_, _05358_, _05352_);
  and (_05360_, _05359_, _05347_);
  and (_05361_, _03898_, _03494_);
  and (_05362_, _05301_, _05361_);
  and (_05363_, _05362_, _05293_);
  and (_05364_, _05363_, \oc8051_golden_model_1.P0 [7]);
  not (_05365_, _05364_);
  nor (_05366_, _03556_, _04559_);
  and (_05367_, _05366_, _05328_);
  and (_05368_, _05367_, _05362_);
  and (_05369_, _05368_, \oc8051_golden_model_1.PSW [7]);
  and (_05370_, _05366_, _05335_);
  and (_05371_, _05370_, _05362_);
  and (_05372_, _05371_, \oc8051_golden_model_1.ACC [7]);
  nor (_05373_, _05372_, _05369_);
  nor (_05374_, _04308_, _03853_);
  and (_05375_, _05374_, _05291_);
  and (_05376_, _05375_, _05333_);
  and (_05377_, _05376_, \oc8051_golden_model_1.IP [7]);
  and (_05378_, _05374_, _05366_);
  and (_05379_, _05378_, _05362_);
  and (_05380_, _05379_, \oc8051_golden_model_1.B [7]);
  nor (_05381_, _05380_, _05377_);
  and (_05382_, _05381_, _05373_);
  and (_05383_, _05362_, _05329_);
  and (_05384_, _05383_, \oc8051_golden_model_1.P1 [7]);
  not (_05385_, _05384_);
  and (_05386_, _05362_, _05336_);
  and (_05387_, _05386_, \oc8051_golden_model_1.P2 [7]);
  and (_05388_, _05375_, _05362_);
  and (_05389_, _05388_, \oc8051_golden_model_1.P3 [7]);
  nor (_05390_, _05389_, _05387_);
  and (_05391_, _05390_, _05385_);
  and (_05392_, _05391_, _05382_);
  and (_05393_, _05392_, _05365_);
  and (_05394_, _05393_, _05360_);
  and (_05395_, _05394_, _05342_);
  and (_05396_, _05395_, _05290_);
  not (_05397_, _05396_);
  nand (_05398_, _04276_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand (_05399_, _04441_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_05400_, _05399_, _04440_);
  nand (_05401_, _05400_, _05398_);
  nand (_05402_, _04441_, \oc8051_golden_model_1.IRAM[3] [6]);
  nand (_05403_, _04276_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_05404_, _05403_, _04446_);
  nand (_05405_, _05404_, _05402_);
  nand (_05406_, _05405_, _05401_);
  nand (_05407_, _05406_, _04011_);
  nand (_05408_, _04441_, \oc8051_golden_model_1.IRAM[7] [6]);
  nand (_05409_, _04276_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_05410_, _05409_, _04446_);
  nand (_05411_, _05410_, _05408_);
  nand (_05412_, _04276_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand (_05413_, _04441_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_05414_, _05413_, _04440_);
  nand (_05415_, _05414_, _05412_);
  nand (_05416_, _05415_, _05411_);
  nand (_05417_, _05416_, _04452_);
  nand (_05418_, _05417_, _05407_);
  nand (_05419_, _05418_, _03822_);
  nand (_05420_, _04441_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_05421_, _04276_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_05422_, _05421_, _04446_);
  nand (_05423_, _05422_, _05420_);
  nand (_05424_, _04276_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_05425_, _04441_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_05426_, _05425_, _04440_);
  nand (_05427_, _05426_, _05424_);
  nand (_05428_, _05427_, _05423_);
  nand (_05429_, _05428_, _04011_);
  nand (_05430_, _04441_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_05431_, _04276_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_05432_, _05431_, _04446_);
  nand (_05433_, _05432_, _05430_);
  nand (_05434_, _04276_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_05435_, _04441_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_05436_, _05435_, _04440_);
  nand (_05437_, _05436_, _05434_);
  nand (_05438_, _05437_, _05433_);
  nand (_05439_, _05438_, _04452_);
  nand (_05440_, _05439_, _05429_);
  nand (_05441_, _05440_, _04466_);
  nand (_05442_, _05441_, _05419_);
  or (_05443_, _05442_, _03463_);
  and (_05444_, _05297_, \oc8051_golden_model_1.DPH [6]);
  not (_05445_, _05444_);
  and (_05446_, _05304_, \oc8051_golden_model_1.TH0 [6]);
  and (_05447_, _05309_, \oc8051_golden_model_1.TL1 [6]);
  nor (_05448_, _05447_, _05446_);
  and (_05449_, _05448_, _05445_);
  and (_05450_, _05315_, \oc8051_golden_model_1.SP [6]);
  and (_05451_, _05319_, \oc8051_golden_model_1.DPL [6]);
  nor (_05452_, _05451_, _05450_);
  and (_05453_, _05323_, \oc8051_golden_model_1.PCON [6]);
  not (_05454_, _05453_);
  and (_05455_, _05330_, \oc8051_golden_model_1.SBUF [6]);
  and (_05456_, _05337_, \oc8051_golden_model_1.IE [6]);
  nor (_05457_, _05456_, _05455_);
  and (_05458_, _05457_, _05454_);
  and (_05459_, _05458_, _05452_);
  and (_05460_, _05459_, _05449_);
  and (_05461_, _05343_, \oc8051_golden_model_1.TMOD [6]);
  and (_05462_, _05345_, \oc8051_golden_model_1.SCON [6]);
  nor (_05463_, _05462_, _05461_);
  and (_05464_, _05350_, \oc8051_golden_model_1.TL0 [6]);
  not (_05465_, _05464_);
  and (_05466_, _05353_, \oc8051_golden_model_1.TCON [6]);
  and (_05467_, _05356_, \oc8051_golden_model_1.TH1 [6]);
  nor (_05468_, _05467_, _05466_);
  and (_05469_, _05468_, _05465_);
  and (_05470_, _05469_, _05463_);
  and (_05471_, _05376_, \oc8051_golden_model_1.IP [6]);
  and (_05472_, _05379_, \oc8051_golden_model_1.B [6]);
  nor (_05473_, _05472_, _05471_);
  and (_05474_, _05368_, \oc8051_golden_model_1.PSW [6]);
  and (_05475_, _05371_, \oc8051_golden_model_1.ACC [6]);
  nor (_05476_, _05475_, _05474_);
  and (_05477_, _05476_, _05473_);
  and (_05478_, _05363_, \oc8051_golden_model_1.P0 [6]);
  not (_05479_, _05478_);
  and (_05480_, _05383_, \oc8051_golden_model_1.P1 [6]);
  not (_05481_, _05480_);
  and (_05482_, _05386_, \oc8051_golden_model_1.P2 [6]);
  and (_05483_, _05388_, \oc8051_golden_model_1.P3 [6]);
  nor (_05484_, _05483_, _05482_);
  and (_05485_, _05484_, _05481_);
  and (_05486_, _05485_, _05479_);
  and (_05487_, _05486_, _05477_);
  and (_05488_, _05487_, _05470_);
  and (_05489_, _05488_, _05460_);
  and (_05490_, _05489_, _05443_);
  not (_05491_, _05490_);
  not (_05492_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_05493_, _04441_, _05492_);
  not (_05494_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_05495_, _04276_, _05494_);
  and (_05496_, _05495_, _04440_);
  nand (_05497_, _05496_, _05493_);
  not (_05498_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_05499_, _04276_, _05498_);
  not (_05500_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05501_, _04441_, _05500_);
  and (_05502_, _05501_, _04446_);
  nand (_05503_, _05502_, _05499_);
  nand (_05504_, _05503_, _05497_);
  nand (_05505_, _05504_, _04011_);
  not (_05506_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_05507_, _04276_, _05506_);
  not (_05508_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_05509_, _04441_, _05508_);
  and (_05510_, _05509_, _04446_);
  nand (_05511_, _05510_, _05507_);
  not (_05512_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_05513_, _04441_, _05512_);
  not (_05514_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_05515_, _04276_, _05514_);
  and (_05516_, _05515_, _04440_);
  nand (_05517_, _05516_, _05513_);
  nand (_05518_, _05517_, _05511_);
  nand (_05519_, _05518_, _04452_);
  nand (_05520_, _05519_, _05505_);
  nand (_05521_, _05520_, _03822_);
  not (_05522_, \oc8051_golden_model_1.IRAM[11] [5]);
  or (_05523_, _04276_, _05522_);
  not (_05524_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_05525_, _04441_, _05524_);
  and (_05526_, _05525_, _04446_);
  nand (_05527_, _05526_, _05523_);
  not (_05528_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_05529_, _04441_, _05528_);
  not (_05530_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_05531_, _04276_, _05530_);
  and (_05532_, _05531_, _04440_);
  nand (_05533_, _05532_, _05529_);
  nand (_05534_, _05533_, _05527_);
  nand (_05535_, _05534_, _04011_);
  not (_05536_, \oc8051_golden_model_1.IRAM[15] [5]);
  or (_05537_, _04276_, _05536_);
  not (_05538_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_05539_, _04441_, _05538_);
  and (_05540_, _05539_, _04446_);
  nand (_05541_, _05540_, _05537_);
  not (_05542_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_05543_, _04441_, _05542_);
  not (_05544_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_05545_, _04276_, _05544_);
  and (_05546_, _05545_, _04440_);
  nand (_05547_, _05546_, _05543_);
  nand (_05548_, _05547_, _05541_);
  nand (_05549_, _05548_, _04452_);
  nand (_05550_, _05549_, _05535_);
  nand (_05551_, _05550_, _04466_);
  nand (_05552_, _05551_, _05521_);
  or (_05553_, _05552_, _03463_);
  and (_05554_, _05297_, \oc8051_golden_model_1.DPH [5]);
  not (_05555_, _05554_);
  and (_05556_, _05304_, \oc8051_golden_model_1.TH0 [5]);
  and (_05557_, _05309_, \oc8051_golden_model_1.TL1 [5]);
  nor (_05558_, _05557_, _05556_);
  and (_05559_, _05558_, _05555_);
  and (_05560_, _05315_, \oc8051_golden_model_1.SP [5]);
  and (_05561_, _05319_, \oc8051_golden_model_1.DPL [5]);
  nor (_05562_, _05561_, _05560_);
  and (_05563_, _05323_, \oc8051_golden_model_1.PCON [5]);
  not (_05564_, _05563_);
  and (_05565_, _05330_, \oc8051_golden_model_1.SBUF [5]);
  and (_05566_, _05337_, \oc8051_golden_model_1.IE [5]);
  nor (_05567_, _05566_, _05565_);
  and (_05568_, _05567_, _05564_);
  and (_05569_, _05568_, _05562_);
  and (_05570_, _05569_, _05559_);
  and (_05571_, _05343_, \oc8051_golden_model_1.TMOD [5]);
  and (_05572_, _05345_, \oc8051_golden_model_1.SCON [5]);
  nor (_05573_, _05572_, _05571_);
  and (_05574_, _05350_, \oc8051_golden_model_1.TL0 [5]);
  not (_05575_, _05574_);
  and (_05576_, _05353_, \oc8051_golden_model_1.TCON [5]);
  and (_05577_, _05356_, \oc8051_golden_model_1.TH1 [5]);
  nor (_05578_, _05577_, _05576_);
  and (_05579_, _05578_, _05575_);
  and (_05580_, _05579_, _05573_);
  and (_05581_, _05376_, \oc8051_golden_model_1.IP [5]);
  and (_05582_, _05371_, \oc8051_golden_model_1.ACC [5]);
  nor (_05583_, _05582_, _05581_);
  and (_05584_, _05368_, \oc8051_golden_model_1.PSW [5]);
  and (_05585_, _05379_, \oc8051_golden_model_1.B [5]);
  nor (_05586_, _05585_, _05584_);
  and (_05587_, _05586_, _05583_);
  and (_05588_, _05363_, \oc8051_golden_model_1.P0 [5]);
  not (_05589_, _05588_);
  and (_05590_, _05383_, \oc8051_golden_model_1.P1 [5]);
  not (_05591_, _05590_);
  and (_05592_, _05386_, \oc8051_golden_model_1.P2 [5]);
  and (_05593_, _05388_, \oc8051_golden_model_1.P3 [5]);
  nor (_05594_, _05593_, _05592_);
  and (_05595_, _05594_, _05591_);
  and (_05596_, _05595_, _05589_);
  and (_05597_, _05596_, _05587_);
  and (_05598_, _05597_, _05580_);
  and (_05599_, _05598_, _05570_);
  and (_05600_, _05599_, _05553_);
  not (_05601_, _05600_);
  or (_05602_, _04944_, _03463_);
  and (_05603_, _05368_, \oc8051_golden_model_1.PSW [3]);
  not (_05604_, _05603_);
  and (_05605_, _05376_, \oc8051_golden_model_1.IP [3]);
  not (_05606_, _05605_);
  and (_05607_, _05379_, \oc8051_golden_model_1.B [3]);
  and (_05608_, _05371_, \oc8051_golden_model_1.ACC [3]);
  nor (_05609_, _05608_, _05607_);
  and (_05610_, _05609_, _05606_);
  and (_05611_, _05610_, _05604_);
  and (_05612_, _05353_, \oc8051_golden_model_1.TCON [3]);
  and (_05613_, _05304_, \oc8051_golden_model_1.TH0 [3]);
  nor (_05614_, _05613_, _05612_);
  and (_05615_, _05309_, \oc8051_golden_model_1.TL1 [3]);
  and (_05616_, _05383_, \oc8051_golden_model_1.P1 [3]);
  nor (_05617_, _05616_, _05615_);
  and (_05618_, _05617_, _05614_);
  and (_05619_, _05345_, \oc8051_golden_model_1.SCON [3]);
  and (_05620_, _05356_, \oc8051_golden_model_1.TH1 [3]);
  nor (_05621_, _05620_, _05619_);
  and (_05622_, _05350_, \oc8051_golden_model_1.TL0 [3]);
  and (_05623_, _05343_, \oc8051_golden_model_1.TMOD [3]);
  nor (_05624_, _05623_, _05622_);
  and (_05625_, _05624_, _05621_);
  and (_05626_, _05625_, _05618_);
  and (_05627_, _05323_, \oc8051_golden_model_1.PCON [3]);
  not (_05628_, _05627_);
  and (_05629_, _05330_, \oc8051_golden_model_1.SBUF [3]);
  and (_05630_, _05337_, \oc8051_golden_model_1.IE [3]);
  nor (_05631_, _05630_, _05629_);
  and (_05632_, _05631_, _05628_);
  and (_05633_, _05386_, \oc8051_golden_model_1.P2 [3]);
  and (_05634_, _05388_, \oc8051_golden_model_1.P3 [3]);
  nor (_05635_, _05634_, _05633_);
  and (_05636_, _05635_, _05632_);
  and (_05637_, _05297_, \oc8051_golden_model_1.DPH [3]);
  not (_05638_, _05637_);
  and (_05639_, _05315_, \oc8051_golden_model_1.SP [3]);
  and (_05640_, _05319_, \oc8051_golden_model_1.DPL [3]);
  nor (_05641_, _05640_, _05639_);
  and (_05642_, _05641_, _05638_);
  and (_05643_, _05363_, \oc8051_golden_model_1.P0 [3]);
  not (_05644_, _05643_);
  and (_05645_, _05644_, _05642_);
  and (_05646_, _05645_, _05636_);
  and (_05647_, _05646_, _05626_);
  and (_05648_, _05647_, _05611_);
  and (_05649_, _05648_, _05602_);
  not (_05650_, _05649_);
  or (_05651_, _04699_, _03463_);
  and (_05652_, _05323_, \oc8051_golden_model_1.PCON [1]);
  not (_05653_, _05652_);
  and (_05654_, _05330_, \oc8051_golden_model_1.SBUF [1]);
  and (_05655_, _05337_, \oc8051_golden_model_1.IE [1]);
  nor (_05656_, _05655_, _05654_);
  and (_05657_, _05656_, _05653_);
  and (_05658_, _05353_, \oc8051_golden_model_1.TCON [1]);
  not (_05659_, _05658_);
  and (_05660_, _05383_, \oc8051_golden_model_1.P1 [1]);
  not (_05661_, _05660_);
  and (_05662_, _05386_, \oc8051_golden_model_1.P2 [1]);
  and (_05663_, _05388_, \oc8051_golden_model_1.P3 [1]);
  nor (_05664_, _05663_, _05662_);
  and (_05665_, _05664_, _05661_);
  and (_05666_, _05665_, _05659_);
  and (_05667_, _05363_, \oc8051_golden_model_1.P0 [1]);
  not (_05668_, _05667_);
  and (_05669_, _05376_, \oc8051_golden_model_1.IP [1]);
  and (_05670_, _05379_, \oc8051_golden_model_1.B [1]);
  nor (_05671_, _05670_, _05669_);
  and (_05672_, _05368_, \oc8051_golden_model_1.PSW [1]);
  and (_05673_, _05371_, \oc8051_golden_model_1.ACC [1]);
  nor (_05674_, _05673_, _05672_);
  and (_05675_, _05674_, _05671_);
  and (_05676_, _05675_, _05668_);
  and (_05677_, _05676_, _05666_);
  and (_05678_, _05677_, _05657_);
  and (_05679_, _05297_, \oc8051_golden_model_1.DPH [1]);
  not (_05680_, _05679_);
  and (_05681_, _05315_, \oc8051_golden_model_1.SP [1]);
  and (_05682_, _05319_, \oc8051_golden_model_1.DPL [1]);
  nor (_05683_, _05682_, _05681_);
  and (_05684_, _05683_, _05680_);
  and (_05685_, _05350_, \oc8051_golden_model_1.TL0 [1]);
  and (_05686_, _05345_, \oc8051_golden_model_1.SCON [1]);
  nor (_05687_, _05686_, _05685_);
  and (_05688_, _05343_, \oc8051_golden_model_1.TMOD [1]);
  and (_05689_, _05304_, \oc8051_golden_model_1.TH0 [1]);
  nor (_05690_, _05689_, _05688_);
  and (_05691_, _05309_, \oc8051_golden_model_1.TL1 [1]);
  and (_05692_, _05356_, \oc8051_golden_model_1.TH1 [1]);
  nor (_05693_, _05692_, _05691_);
  and (_05694_, _05693_, _05690_);
  and (_05695_, _05694_, _05687_);
  and (_05696_, _05695_, _05684_);
  and (_05697_, _05696_, _05678_);
  and (_05698_, _05697_, _05651_);
  not (_05699_, _05698_);
  or (_05700_, _04510_, _03463_);
  and (_05701_, _05356_, \oc8051_golden_model_1.TH1 [0]);
  and (_05702_, _05330_, \oc8051_golden_model_1.SBUF [0]);
  nor (_05703_, _05702_, _05701_);
  and (_05704_, _05343_, \oc8051_golden_model_1.TMOD [0]);
  and (_05705_, _05345_, \oc8051_golden_model_1.SCON [0]);
  nor (_05706_, _05705_, _05704_);
  and (_05707_, _05706_, _05703_);
  and (_05708_, _05319_, \oc8051_golden_model_1.DPL [0]);
  not (_05709_, _05708_);
  and (_05710_, _05350_, \oc8051_golden_model_1.TL0 [0]);
  and (_05711_, _05337_, \oc8051_golden_model_1.IE [0]);
  nor (_05712_, _05711_, _05710_);
  and (_05713_, _05712_, _05709_);
  and (_05714_, _05315_, \oc8051_golden_model_1.SP [0]);
  and (_05715_, _05297_, \oc8051_golden_model_1.DPH [0]);
  nor (_05716_, _05715_, _05714_);
  and (_05717_, _05716_, _05713_);
  and (_05718_, _05717_, _05707_);
  not (_05719_, _05718_);
  and (_05720_, _05383_, \oc8051_golden_model_1.P1 [0]);
  and (_05721_, _05353_, \oc8051_golden_model_1.TCON [0]);
  and (_05722_, _05386_, \oc8051_golden_model_1.P2 [0]);
  and (_05723_, _05388_, \oc8051_golden_model_1.P3 [0]);
  or (_05724_, _05723_, _05722_);
  or (_05725_, _05724_, _05721_);
  or (_05726_, _05725_, _05720_);
  and (_05727_, _05376_, \oc8051_golden_model_1.IP [0]);
  and (_05728_, _05379_, \oc8051_golden_model_1.B [0]);
  nor (_05729_, _05728_, _05727_);
  and (_05730_, _05368_, \oc8051_golden_model_1.PSW [0]);
  and (_05731_, _05371_, \oc8051_golden_model_1.ACC [0]);
  nor (_05732_, _05731_, _05730_);
  and (_05733_, _05732_, _05729_);
  and (_05734_, _05304_, \oc8051_golden_model_1.TH0 [0]);
  and (_05735_, _05309_, \oc8051_golden_model_1.TL1 [0]);
  nor (_05736_, _05735_, _05734_);
  and (_05737_, _05736_, _05733_);
  and (_05738_, _05363_, \oc8051_golden_model_1.P0 [0]);
  and (_05739_, _05323_, \oc8051_golden_model_1.PCON [0]);
  nor (_05740_, _05739_, _05738_);
  nand (_05741_, _05740_, _05737_);
  or (_05742_, _05741_, _05726_);
  nor (_05743_, _05742_, _05719_);
  nand (_05744_, _05743_, _05700_);
  and (_05745_, _05744_, _05699_);
  or (_05746_, _05130_, _03463_);
  and (_05747_, _05356_, \oc8051_golden_model_1.TH1 [2]);
  and (_05748_, _05330_, \oc8051_golden_model_1.SBUF [2]);
  nor (_05749_, _05748_, _05747_);
  and (_05750_, _05343_, \oc8051_golden_model_1.TMOD [2]);
  and (_05751_, _05345_, \oc8051_golden_model_1.SCON [2]);
  nor (_05752_, _05751_, _05750_);
  and (_05753_, _05752_, _05749_);
  and (_05754_, _05319_, \oc8051_golden_model_1.DPL [2]);
  not (_05755_, _05754_);
  and (_05756_, _05350_, \oc8051_golden_model_1.TL0 [2]);
  and (_05757_, _05337_, \oc8051_golden_model_1.IE [2]);
  nor (_05758_, _05757_, _05756_);
  and (_05759_, _05758_, _05755_);
  and (_05760_, _05315_, \oc8051_golden_model_1.SP [2]);
  and (_05761_, _05297_, \oc8051_golden_model_1.DPH [2]);
  nor (_05762_, _05761_, _05760_);
  and (_05763_, _05762_, _05759_);
  and (_05764_, _05763_, _05753_);
  not (_05765_, _05764_);
  and (_05766_, _05353_, \oc8051_golden_model_1.TCON [2]);
  and (_05767_, _05383_, \oc8051_golden_model_1.P1 [2]);
  and (_05768_, _05386_, \oc8051_golden_model_1.P2 [2]);
  and (_05769_, _05388_, \oc8051_golden_model_1.P3 [2]);
  or (_05770_, _05769_, _05768_);
  or (_05771_, _05770_, _05767_);
  or (_05772_, _05771_, _05766_);
  and (_05773_, _05363_, \oc8051_golden_model_1.P0 [2]);
  not (_05774_, _05773_);
  and (_05775_, _05376_, \oc8051_golden_model_1.IP [2]);
  and (_05776_, _05379_, \oc8051_golden_model_1.B [2]);
  nor (_05777_, _05776_, _05775_);
  and (_05778_, _05368_, \oc8051_golden_model_1.PSW [2]);
  and (_05779_, _05371_, \oc8051_golden_model_1.ACC [2]);
  nor (_05780_, _05779_, _05778_);
  and (_05781_, _05780_, _05777_);
  nand (_05782_, _05781_, _05774_);
  and (_05783_, _05323_, \oc8051_golden_model_1.PCON [2]);
  not (_05784_, _05783_);
  and (_05785_, _05304_, \oc8051_golden_model_1.TH0 [2]);
  and (_05786_, _05309_, \oc8051_golden_model_1.TL1 [2]);
  nor (_05787_, _05786_, _05785_);
  nand (_05788_, _05787_, _05784_);
  or (_05789_, _05788_, _05782_);
  or (_05790_, _05789_, _05772_);
  nor (_05791_, _05790_, _05765_);
  and (_05792_, _05791_, _05746_);
  not (_05793_, _05792_);
  and (_05794_, _05793_, _05745_);
  and (_05795_, _05794_, _05650_);
  nand (_05796_, _04276_, \oc8051_golden_model_1.IRAM[0] [4]);
  nand (_05797_, _04441_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_05798_, _05797_, _04440_);
  nand (_05799_, _05798_, _05796_);
  nand (_05800_, _04441_, \oc8051_golden_model_1.IRAM[3] [4]);
  nand (_05801_, _04276_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_05802_, _05801_, _04446_);
  nand (_05803_, _05802_, _05800_);
  nand (_05804_, _05803_, _05799_);
  nand (_05805_, _05804_, _04011_);
  nand (_05806_, _04441_, \oc8051_golden_model_1.IRAM[7] [4]);
  nand (_05807_, _04276_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_05808_, _05807_, _04446_);
  nand (_05809_, _05808_, _05806_);
  nand (_05810_, _04276_, \oc8051_golden_model_1.IRAM[4] [4]);
  nand (_05811_, _04441_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_05812_, _05811_, _04440_);
  nand (_05813_, _05812_, _05810_);
  nand (_05814_, _05813_, _05809_);
  nand (_05815_, _05814_, _04452_);
  nand (_05816_, _05815_, _05805_);
  nand (_05817_, _05816_, _03822_);
  nand (_05818_, _04441_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_05819_, _04276_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_05820_, _05819_, _04446_);
  nand (_05821_, _05820_, _05818_);
  nand (_05822_, _04276_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_05823_, _04441_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_05824_, _05823_, _04440_);
  nand (_05825_, _05824_, _05822_);
  nand (_05826_, _05825_, _05821_);
  nand (_05827_, _05826_, _04011_);
  nand (_05828_, _04441_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_05829_, _04276_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_05830_, _05829_, _04446_);
  nand (_05831_, _05830_, _05828_);
  nand (_05832_, _04276_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_05833_, _04441_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_05834_, _05833_, _04440_);
  nand (_05835_, _05834_, _05832_);
  nand (_05836_, _05835_, _05831_);
  nand (_05837_, _05836_, _04452_);
  nand (_05838_, _05837_, _05827_);
  nand (_05839_, _05838_, _04466_);
  nand (_05840_, _05839_, _05817_);
  or (_05841_, _05840_, _03463_);
  and (_05842_, _05323_, \oc8051_golden_model_1.PCON [4]);
  not (_05843_, _05842_);
  and (_05844_, _05330_, \oc8051_golden_model_1.SBUF [4]);
  and (_05845_, _05337_, \oc8051_golden_model_1.IE [4]);
  nor (_05846_, _05845_, _05844_);
  and (_05847_, _05846_, _05843_);
  and (_05848_, _05353_, \oc8051_golden_model_1.TCON [4]);
  not (_05849_, _05848_);
  and (_05850_, _05383_, \oc8051_golden_model_1.P1 [4]);
  not (_05851_, _05850_);
  and (_05852_, _05386_, \oc8051_golden_model_1.P2 [4]);
  and (_05853_, _05388_, \oc8051_golden_model_1.P3 [4]);
  nor (_05854_, _05853_, _05852_);
  and (_05855_, _05854_, _05851_);
  and (_05856_, _05855_, _05849_);
  and (_05857_, _05363_, \oc8051_golden_model_1.P0 [4]);
  not (_05858_, _05857_);
  and (_05859_, _05368_, \oc8051_golden_model_1.PSW [4]);
  and (_05860_, _05379_, \oc8051_golden_model_1.B [4]);
  nor (_05861_, _05860_, _05859_);
  and (_05862_, _05376_, \oc8051_golden_model_1.IP [4]);
  and (_05863_, _05371_, \oc8051_golden_model_1.ACC [4]);
  nor (_05864_, _05863_, _05862_);
  and (_05865_, _05864_, _05861_);
  and (_05866_, _05865_, _05858_);
  and (_05867_, _05866_, _05856_);
  and (_05868_, _05867_, _05847_);
  and (_05869_, _05297_, \oc8051_golden_model_1.DPH [4]);
  not (_05870_, _05869_);
  and (_05871_, _05315_, \oc8051_golden_model_1.SP [4]);
  and (_05872_, _05319_, \oc8051_golden_model_1.DPL [4]);
  nor (_05873_, _05872_, _05871_);
  and (_05874_, _05873_, _05870_);
  and (_05875_, _05343_, \oc8051_golden_model_1.TMOD [4]);
  and (_05876_, _05345_, \oc8051_golden_model_1.SCON [4]);
  nor (_05877_, _05876_, _05875_);
  and (_05878_, _05304_, \oc8051_golden_model_1.TH0 [4]);
  and (_05879_, _05356_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05880_, _05879_, _05878_);
  and (_05881_, _05350_, \oc8051_golden_model_1.TL0 [4]);
  and (_05882_, _05309_, \oc8051_golden_model_1.TL1 [4]);
  nor (_05883_, _05882_, _05881_);
  and (_05884_, _05883_, _05880_);
  and (_05885_, _05884_, _05877_);
  and (_05886_, _05885_, _05874_);
  and (_05887_, _05886_, _05868_);
  and (_05888_, _05887_, _05841_);
  not (_05889_, _05888_);
  and (_05890_, _05889_, _05795_);
  and (_05891_, _05890_, _05601_);
  and (_05892_, _05891_, _05491_);
  nor (_05893_, _05892_, _05397_);
  and (_05894_, _05892_, _05397_);
  nor (_05895_, _05894_, _05893_);
  and (_05896_, _05895_, _04633_);
  not (_05897_, _05289_);
  and (_05898_, _04698_, _04676_);
  and (_05899_, _05898_, _04491_);
  nor (_05900_, _05130_, _04944_);
  and (_05901_, _05900_, _05899_);
  nor (_05902_, _05840_, _05552_);
  and (_05903_, _05902_, _05901_);
  or (_05904_, _05903_, _05897_);
  and (_05905_, _05442_, _05289_);
  nor (_05906_, _05442_, _05289_);
  nor (_05907_, _05906_, _05905_);
  not (_05908_, _05907_);
  nand (_05909_, _05908_, _05903_);
  and (_05910_, _05909_, _05904_);
  and (_05911_, _04563_, _03241_);
  or (_05912_, _05911_, _04840_);
  nor (_05913_, _05912_, _04642_);
  or (_05914_, _05913_, _05910_);
  and (_05915_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_05916_, _05915_, \oc8051_golden_model_1.PC [6]);
  and (_05917_, _02942_, \oc8051_golden_model_1.PC [2]);
  and (_05918_, _05917_, \oc8051_golden_model_1.PC [3]);
  and (_05919_, _05918_, _05916_);
  and (_05920_, _05919_, \oc8051_golden_model_1.PC [7]);
  nor (_05921_, _05919_, \oc8051_golden_model_1.PC [7]);
  nor (_05922_, _05921_, _05920_);
  not (_05923_, _05922_);
  nand (_05924_, _05923_, _03686_);
  not (_05925_, _04595_);
  not (_05926_, _04597_);
  not (_05927_, _04590_);
  and (_05928_, _03712_, _01758_);
  and (_05929_, _03745_, _01723_);
  nor (_05930_, _05929_, _05928_);
  and (_05931_, _03748_, _01778_);
  and (_05932_, _03729_, _01714_);
  nor (_05933_, _05932_, _05931_);
  and (_05934_, _05933_, _05930_);
  and (_05935_, _03743_, _01746_);
  and (_05936_, _03736_, _01774_);
  nor (_05937_, _05936_, _05935_);
  and (_05938_, _03721_, _01765_);
  and (_05939_, _03761_, _01762_);
  nor (_05940_, _05939_, _05938_);
  and (_05941_, _05940_, _05937_);
  and (_05942_, _05941_, _05934_);
  and (_05943_, _03759_, _01749_);
  and (_05944_, _03754_, _01755_);
  nor (_05945_, _05944_, _05943_);
  and (_05946_, _03756_, _01730_);
  and (_05947_, _03732_, _01704_);
  nor (_05948_, _05947_, _05946_);
  and (_05949_, _05948_, _05945_);
  and (_05950_, _03750_, _01718_);
  and (_05951_, _03738_, _01739_);
  nor (_05952_, _05951_, _05950_);
  and (_05953_, _03716_, _01709_);
  and (_05954_, _03725_, _01673_);
  nor (_05955_, _05954_, _05953_);
  and (_05956_, _05955_, _05952_);
  and (_05957_, _05956_, _05949_);
  and (_05958_, _05957_, _05942_);
  and (_05959_, _05958_, _05396_);
  nor (_05960_, _05958_, _05396_);
  nor (_05961_, _05960_, _05959_);
  and (_05962_, _05961_, _04592_);
  not (_05963_, _04563_);
  and (_05964_, _04839_, _05963_);
  nor (_05965_, _05964_, _04813_);
  nor (_05966_, _05965_, _04816_);
  and (_05967_, _05966_, _04582_);
  or (_05968_, _05967_, _03463_);
  and (_05969_, _04197_, _03219_);
  not (_05970_, _05969_);
  nor (_05971_, _05970_, _03463_);
  not (_05972_, _03495_);
  nor (_05973_, _04309_, _05972_);
  nor (_05974_, _03854_, _03560_);
  and (_05975_, _05974_, _05973_);
  and (_05976_, _05975_, _05329_);
  and (_05977_, _05976_, \oc8051_golden_model_1.SCON [7]);
  not (_05978_, _05977_);
  and (_05979_, _05975_, _05336_);
  and (_05980_, _05979_, \oc8051_golden_model_1.IE [7]);
  and (_05981_, _03855_, _03560_);
  and (_05982_, _05981_, _05973_);
  and (_05983_, _05370_, _05982_);
  and (_05985_, _05983_, \oc8051_golden_model_1.ACC [7]);
  nor (_05986_, _05985_, _05980_);
  and (_05988_, _05986_, _05978_);
  and (_05989_, _05975_, _05375_);
  and (_05991_, _05989_, \oc8051_golden_model_1.IP [7]);
  and (_05992_, _05378_, _05982_);
  and (_05994_, _05992_, \oc8051_golden_model_1.B [7]);
  nor (_05995_, _05994_, _05991_);
  and (_05997_, _05975_, _05293_);
  and (_05998_, _05997_, \oc8051_golden_model_1.TCON [7]);
  and (_06000_, _05367_, _05982_);
  and (_06001_, _06000_, \oc8051_golden_model_1.PSW [7]);
  nor (_06003_, _06001_, _05998_);
  and (_06004_, _06003_, _05995_);
  and (_06006_, _06004_, _05988_);
  and (_06007_, _05294_, \oc8051_golden_model_1.P0INREG [7]);
  and (_06009_, _05336_, _05982_);
  and (_06010_, _06009_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_06012_, _06010_, _06007_);
  and (_06013_, _05329_, _05982_);
  and (_06015_, _06013_, \oc8051_golden_model_1.P1INREG [7]);
  and (_06016_, _05375_, _05982_);
  and (_06018_, _06016_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06019_, _06018_, _06015_);
  and (_06021_, _06019_, _06012_);
  and (_06022_, _06021_, _06006_);
  and (_06023_, _06022_, _05290_);
  nor (_06024_, _06023_, _05322_);
  and (_06025_, _05322_, \oc8051_golden_model_1.PSW [7]);
  nor (_06026_, _06025_, _06024_);
  nor (_06027_, _06026_, _05007_);
  not (_06028_, _04533_);
  and (_06029_, _05294_, \oc8051_golden_model_1.P0 [7]);
  and (_06030_, _06016_, \oc8051_golden_model_1.P3 [7]);
  nor (_06031_, _06030_, _06029_);
  and (_06032_, _06013_, \oc8051_golden_model_1.P1 [7]);
  and (_06033_, _06009_, \oc8051_golden_model_1.P2 [7]);
  nor (_06034_, _06033_, _06032_);
  and (_06035_, _06034_, _06031_);
  and (_06036_, _06035_, _06006_);
  and (_06037_, _06036_, _05290_);
  nor (_06038_, _06037_, _05322_);
  or (_06039_, _06038_, _06028_);
  not (_06040_, _04514_);
  not (_06041_, _05322_);
  nand (_06042_, _06037_, _06041_);
  or (_06043_, _06042_, _06040_);
  and (_06044_, _05840_, _05552_);
  and (_06045_, _04699_, _04510_);
  and (_06046_, _05130_, _04944_);
  and (_06047_, _06046_, _06045_);
  and (_06048_, _06047_, _06044_);
  and (_06049_, _06048_, _05442_);
  or (_06050_, _06049_, _05897_);
  nand (_06051_, _06049_, _05897_);
  and (_06052_, _06051_, _06050_);
  or (_06053_, _04395_, _03958_);
  nor (_06054_, _06053_, _04705_);
  or (_06055_, _06054_, _06052_);
  and (_06056_, _05916_, _03207_);
  and (_06057_, _06056_, \oc8051_golden_model_1.PC [7]);
  nor (_06058_, _06056_, \oc8051_golden_model_1.PC [7]);
  nor (_06059_, _06058_, _06057_);
  and (_06060_, _06059_, _03947_);
  not (_06061_, \oc8051_golden_model_1.ACC [7]);
  nor (_06062_, _03947_, _06061_);
  or (_06063_, _06062_, _03958_);
  nor (_06064_, _06063_, _06060_);
  nand (_06065_, _06064_, _05083_);
  and (_06066_, _06065_, _06055_);
  or (_06067_, _06066_, _04509_);
  not (_06068_, _04509_);
  not (_06069_, \oc8051_golden_model_1.SP [2]);
  nor (_06070_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_06071_, _06070_, _06069_);
  nor (_06072_, _06071_, _03596_);
  nor (_06073_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_06074_, _06073_, _03596_);
  and (_06075_, _06074_, _04079_);
  nor (_06076_, _06075_, _06072_);
  nor (_06077_, _03792_, _03521_);
  nor (_06078_, _06077_, _06076_);
  not (_06080_, _06078_);
  not (_06082_, _04551_);
  nand (_06083_, _04944_, _06082_);
  not (_06085_, _06077_);
  and (_06086_, _04551_, _03494_);
  nor (_06088_, _06086_, _06085_);
  nand (_06089_, _06088_, _06083_);
  and (_06091_, _06089_, _06080_);
  not (_06092_, _06091_);
  or (_06094_, _05130_, _04551_);
  nor (_06095_, _06082_, _03898_);
  nor (_06097_, _06095_, _06085_);
  nand (_06098_, _06097_, _06094_);
  nor (_06100_, _06070_, _06069_);
  nor (_06101_, _06100_, _06071_);
  not (_06103_, _06101_);
  nor (_06104_, _06103_, _06077_);
  not (_06106_, _06104_);
  and (_06107_, _06106_, _06098_);
  or (_06109_, _04551_, _04491_);
  and (_06110_, _04551_, _04042_);
  nor (_06112_, _06110_, _06085_);
  nand (_06113_, _06112_, _06109_);
  nor (_06114_, _06077_, \oc8051_golden_model_1.SP [0]);
  not (_06115_, _06114_);
  and (_06116_, _06115_, _06113_);
  or (_06117_, _06116_, \oc8051_golden_model_1.IRAM[13] [7]);
  nor (_06118_, _06077_, _04646_);
  not (_06119_, _06118_);
  and (_06120_, _05898_, _06082_);
  nor (_06121_, _06082_, _04434_);
  or (_06122_, _06121_, _06085_);
  or (_06123_, _06122_, _06120_);
  nand (_06124_, _06123_, _06119_);
  nand (_06125_, _06115_, _06113_);
  or (_06126_, _06125_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_06127_, _06126_, _06124_);
  and (_06128_, _06127_, _06117_);
  or (_06129_, _06125_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_06130_, _06123_, _06119_);
  or (_06131_, _06116_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_06132_, _06131_, _06130_);
  and (_06133_, _06132_, _06129_);
  nor (_06134_, _06133_, _06128_);
  nand (_06135_, _06134_, _06107_);
  not (_06136_, _06107_);
  or (_06137_, _06116_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_06138_, _06125_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_06139_, _06138_, _06124_);
  and (_06140_, _06139_, _06137_);
  or (_06141_, _06125_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_06142_, _06116_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_06143_, _06142_, _06130_);
  and (_06144_, _06143_, _06141_);
  nor (_06145_, _06144_, _06140_);
  nand (_06146_, _06145_, _06136_);
  nand (_06147_, _06146_, _06135_);
  nand (_06148_, _06147_, _06092_);
  or (_06149_, _06125_, _05257_);
  or (_06150_, _06116_, _05259_);
  and (_06151_, _06150_, _06124_);
  nand (_06152_, _06151_, _06149_);
  or (_06153_, _06125_, _05253_);
  or (_06154_, _06116_, _05251_);
  and (_06155_, _06154_, _06130_);
  nand (_06156_, _06155_, _06153_);
  nand (_06157_, _06156_, _06152_);
  nand (_06158_, _06157_, _06107_);
  or (_06159_, _06116_, _05239_);
  or (_06160_, _06125_, _05237_);
  and (_06161_, _06160_, _06124_);
  nand (_06162_, _06161_, _06159_);
  or (_06163_, _06125_, _05245_);
  or (_06164_, _06116_, _05243_);
  and (_06165_, _06164_, _06130_);
  nand (_06166_, _06165_, _06163_);
  nand (_06167_, _06166_, _06162_);
  nand (_06168_, _06167_, _06136_);
  nand (_06169_, _06168_, _06158_);
  nand (_06170_, _06169_, _06091_);
  and (_06171_, _06170_, _06148_);
  or (_06172_, _06171_, _06068_);
  and (_06173_, _06172_, _06067_);
  or (_06174_, _06173_, _04516_);
  not (_06175_, _04516_);
  and (_06176_, _05888_, _05600_);
  not (_06177_, _05744_);
  and (_06178_, _06177_, _05698_);
  and (_06179_, _05792_, _05649_);
  and (_06180_, _06179_, _06178_);
  and (_06181_, _06180_, _06176_);
  and (_06182_, _06181_, _05490_);
  nor (_06183_, _06182_, _05397_);
  and (_06184_, _06182_, _05397_);
  nor (_06185_, _06184_, _06183_);
  or (_06186_, _06185_, _06175_);
  and (_06187_, _06186_, _06174_);
  or (_06188_, _06187_, _04514_);
  and (_06189_, _06188_, _06043_);
  or (_06190_, _06189_, _04857_);
  nor (_06191_, _06059_, _03257_);
  nor (_06192_, _06191_, _04525_);
  and (_06193_, _06192_, _06190_);
  and (_06194_, _05897_, _04525_);
  or (_06195_, _06194_, _04533_);
  or (_06196_, _06195_, _06193_);
  and (_06197_, _06196_, _06039_);
  or (_06198_, _06197_, _03510_);
  and (_06199_, _05363_, \oc8051_golden_model_1.P0INREG [7]);
  not (_06200_, _06199_);
  and (_06201_, _05383_, \oc8051_golden_model_1.P1INREG [7]);
  not (_06202_, _06201_);
  and (_06203_, _05386_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06204_, _05388_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06205_, _06204_, _06203_);
  and (_06206_, _06205_, _06202_);
  and (_06207_, _06206_, _05382_);
  and (_06208_, _06207_, _06200_);
  and (_06209_, _06208_, _05360_);
  and (_06210_, _06209_, _05342_);
  and (_06211_, _06210_, _05290_);
  nand (_06212_, _06211_, _03510_);
  and (_06213_, _06212_, _03508_);
  and (_06214_, _06213_, _06198_);
  nor (_06215_, _06037_, _06041_);
  not (_06216_, _06215_);
  and (_06217_, _06216_, _06042_);
  and (_06218_, _06217_, _03507_);
  or (_06219_, _06218_, _06214_);
  and (_06220_, _06219_, _03253_);
  not (_06221_, _06059_);
  or (_06222_, _06221_, _03253_);
  nand (_06223_, _06222_, _03593_);
  or (_06224_, _06223_, _06220_);
  nand (_06225_, _06211_, _03594_);
  and (_06226_, _06225_, _06224_);
  or (_06227_, _06226_, _04551_);
  and (_06228_, _06171_, _04559_);
  nand (_06229_, _06210_, _04551_);
  or (_06230_, _06229_, _06228_);
  and (_06231_, _06230_, _05007_);
  and (_06232_, _06231_, _06227_);
  or (_06233_, _06232_, _06027_);
  and (_06234_, _06233_, _03278_);
  or (_06235_, _06221_, _03278_);
  nand (_06236_, _06235_, _04568_);
  or (_06237_, _06236_, _06234_);
  not (_06238_, _04568_);
  nand (_06239_, _05289_, _06238_);
  and (_06240_, _06239_, _06237_);
  or (_06241_, _06240_, _05971_);
  not (_06242_, _04569_);
  and (_06243_, _06171_, _06242_);
  or (_06244_, _06243_, _04571_);
  and (_06245_, _06244_, _06241_);
  not (_06246_, _05966_);
  not (_06247_, _05958_);
  nor (_06248_, _06247_, _05289_);
  not (_06249_, _04347_);
  and (_06250_, _06249_, _04172_);
  and (_06251_, _03712_, _02232_);
  and (_06252_, _03745_, _02268_);
  nor (_06253_, _06252_, _06251_);
  and (_06254_, _03748_, _02229_);
  and (_06255_, _03729_, _02249_);
  nor (_06256_, _06255_, _06254_);
  and (_06257_, _06256_, _06253_);
  and (_06258_, _03721_, _02247_);
  and (_06259_, _03761_, _02234_);
  nor (_06260_, _06259_, _06258_);
  and (_06261_, _03736_, _02239_);
  and (_06262_, _03738_, _02257_);
  nor (_06263_, _06262_, _06261_);
  and (_06264_, _06263_, _06260_);
  and (_06265_, _06264_, _06257_);
  and (_06266_, _03759_, _02227_);
  and (_06267_, _03754_, _02259_);
  nor (_06268_, _06267_, _06266_);
  and (_06269_, _03756_, _02261_);
  and (_06270_, _03732_, _02251_);
  nor (_06271_, _06270_, _06269_);
  and (_06272_, _06271_, _06268_);
  and (_06273_, _03750_, _02266_);
  and (_06274_, _03743_, _02236_);
  nor (_06275_, _06274_, _06273_);
  and (_06276_, _03716_, _02241_);
  and (_06277_, _03725_, _02255_);
  nor (_06278_, _06277_, _06276_);
  and (_06279_, _06278_, _06275_);
  and (_06280_, _06279_, _06272_);
  and (_06281_, _06280_, _06265_);
  and (_06282_, _06281_, _06247_);
  and (_06283_, _03761_, _02179_);
  and (_06284_, _03716_, _02189_);
  nor (_06285_, _06284_, _06283_);
  and (_06286_, _03748_, _02174_);
  and (_06287_, _03745_, _02222_);
  nor (_06288_, _06287_, _06286_);
  and (_06289_, _06288_, _06285_);
  and (_06290_, _03759_, _02172_);
  and (_06291_, _03754_, _02213_);
  nor (_06292_, _06291_, _06290_);
  and (_06293_, _03736_, _02182_);
  and (_06294_, _03738_, _02210_);
  nor (_06295_, _06294_, _06293_);
  and (_06296_, _06295_, _06292_);
  and (_06297_, _06296_, _06289_);
  and (_06298_, _03732_, _02202_);
  and (_06299_, _03725_, _02207_);
  nor (_06300_, _06299_, _06298_);
  and (_06301_, _03750_, _02220_);
  and (_06302_, _03756_, _02215_);
  nor (_06303_, _06302_, _06301_);
  and (_06304_, _06303_, _06300_);
  and (_06305_, _03712_, _02177_);
  and (_06306_, _03743_, _02186_);
  nor (_06307_, _06306_, _06305_);
  and (_06308_, _03721_, _02197_);
  and (_06309_, _03729_, _02199_);
  nor (_06310_, _06309_, _06308_);
  and (_06311_, _06310_, _06307_);
  and (_06312_, _06311_, _06304_);
  and (_06313_, _06312_, _06297_);
  and (_06314_, _03761_, _02124_);
  and (_06315_, _03716_, _02133_);
  nor (_06316_, _06315_, _06314_);
  and (_06317_, _03748_, _02119_);
  and (_06318_, _03745_, _02167_);
  nor (_06319_, _06318_, _06317_);
  and (_06320_, _06319_, _06316_);
  and (_06321_, _03736_, _02126_);
  and (_06322_, _03743_, _02130_);
  nor (_06323_, _06322_, _06321_);
  and (_06324_, _03759_, _02117_);
  and (_06325_, _03754_, _02157_);
  nor (_06326_, _06325_, _06324_);
  and (_06327_, _06326_, _06323_);
  and (_06328_, _06327_, _06320_);
  and (_06329_, _03732_, _02146_);
  and (_06330_, _03725_, _02151_);
  nor (_06331_, _06330_, _06329_);
  and (_06332_, _03750_, _02165_);
  and (_06333_, _03756_, _02159_);
  nor (_06334_, _06333_, _06332_);
  and (_06335_, _06334_, _06331_);
  and (_06336_, _03712_, _02122_);
  and (_06337_, _03738_, _02154_);
  nor (_06338_, _06337_, _06336_);
  and (_06339_, _03721_, _02141_);
  and (_06340_, _03729_, _02143_);
  nor (_06341_, _06340_, _06339_);
  and (_06342_, _06341_, _06338_);
  and (_06343_, _06342_, _06335_);
  and (_06344_, _06343_, _06328_);
  and (_06345_, _06344_, _06313_);
  and (_06346_, _06345_, _06282_);
  not (_06347_, _03766_);
  and (_06348_, _03943_, _06347_);
  and (_06349_, _06348_, _06346_);
  and (_06350_, _06349_, _06250_);
  and (_06351_, _06350_, \oc8051_golden_model_1.TL0 [7]);
  not (_06352_, _06351_);
  and (_06353_, _04347_, _04172_);
  and (_06354_, _03943_, _03766_);
  and (_06355_, _06354_, _06353_);
  and (_06356_, _06355_, _06346_);
  and (_06357_, _06356_, \oc8051_golden_model_1.P0INREG [7]);
  not (_06358_, _06313_);
  and (_06359_, _06344_, _06358_);
  and (_06360_, _06359_, _06282_);
  and (_06361_, _06360_, _06355_);
  and (_06362_, _06361_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_06363_, _06362_, _06357_);
  and (_06364_, _06363_, _06352_);
  and (_06365_, _06354_, _06346_);
  not (_06366_, _04172_);
  and (_06367_, _04347_, _06366_);
  and (_06368_, _06367_, _06365_);
  and (_06369_, _06368_, \oc8051_golden_model_1.SP [7]);
  not (_06370_, _06369_);
  and (_06371_, _06367_, _06348_);
  and (_06372_, _06371_, _06346_);
  and (_06373_, _06372_, \oc8051_golden_model_1.TMOD [7]);
  not (_06374_, _06373_);
  not (_06375_, _06344_);
  and (_06376_, _06375_, _06313_);
  and (_06377_, _06376_, _06282_);
  and (_06378_, _06377_, _06355_);
  and (_06379_, _06378_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_06380_, _06344_, _06313_);
  and (_06381_, _06380_, _06282_);
  and (_06382_, _06381_, _06355_);
  and (_06383_, _06382_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_06384_, _06383_, _06379_);
  and (_06385_, _06384_, _06374_);
  and (_06386_, _06385_, _06370_);
  and (_06387_, _06386_, _06364_);
  and (_06388_, _06353_, _06348_);
  and (_06389_, _06388_, _06360_);
  and (_06390_, _06389_, \oc8051_golden_model_1.IE [7]);
  not (_06391_, _06390_);
  and (_06392_, _06388_, _06377_);
  and (_06393_, _06392_, \oc8051_golden_model_1.SCON [7]);
  and (_06394_, _06377_, _06371_);
  and (_06395_, _06394_, \oc8051_golden_model_1.SBUF [7]);
  nor (_06396_, _06395_, _06393_);
  and (_06397_, _06396_, _06391_);
  nor (_06398_, _04347_, _04172_);
  and (_06399_, _06398_, _06346_);
  and (_06400_, _06399_, _06354_);
  and (_06401_, _06400_, \oc8051_golden_model_1.DPH [7]);
  nor (_06402_, _03943_, _03766_);
  and (_06403_, _06402_, _06346_);
  and (_06404_, _06403_, _06367_);
  and (_06405_, _06404_, \oc8051_golden_model_1.TH1 [7]);
  nor (_06406_, _06405_, _06401_);
  and (_06407_, _06406_, _06397_);
  and (_06408_, _06407_, _06387_);
  and (_06409_, _06403_, _06353_);
  and (_06410_, _06409_, \oc8051_golden_model_1.TH0 [7]);
  and (_06411_, _06399_, _06348_);
  and (_06412_, _06411_, \oc8051_golden_model_1.TL1 [7]);
  nor (_06413_, _06412_, _06410_);
  not (_06414_, _03943_);
  and (_06415_, _06414_, _03766_);
  and (_06416_, _06415_, _06399_);
  and (_06417_, _06416_, \oc8051_golden_model_1.PCON [7]);
  and (_06418_, _06353_, _06349_);
  and (_06419_, _06418_, \oc8051_golden_model_1.TCON [7]);
  nor (_06420_, _06419_, _06417_);
  and (_06421_, _06420_, _06413_);
  and (_06422_, _06365_, _06250_);
  and (_06423_, _06422_, \oc8051_golden_model_1.DPL [7]);
  not (_06424_, _06423_);
  nor (_06425_, _06281_, _05958_);
  and (_06426_, _06425_, _06355_);
  and (_06427_, _06426_, _06376_);
  and (_06428_, _06427_, \oc8051_golden_model_1.PSW [7]);
  and (_06429_, _06426_, _06380_);
  and (_06430_, _06429_, \oc8051_golden_model_1.B [7]);
  nor (_06431_, _06430_, _06428_);
  and (_06432_, _06426_, _06359_);
  and (_06433_, _06432_, \oc8051_golden_model_1.ACC [7]);
  and (_06434_, _06388_, _06282_);
  and (_06435_, _06434_, _06380_);
  and (_06436_, _06435_, \oc8051_golden_model_1.IP [7]);
  nor (_06437_, _06436_, _06433_);
  and (_06438_, _06437_, _06431_);
  and (_06439_, _06438_, _06424_);
  and (_06440_, _06439_, _06421_);
  and (_06441_, _06440_, _06408_);
  not (_06442_, _06441_);
  nor (_06443_, _06442_, _06248_);
  nor (_06444_, _06443_, _06242_);
  or (_06445_, _06444_, _06246_);
  or (_06446_, _06445_, _06245_);
  and (_06447_, _06446_, _05968_);
  and (_06448_, _06247_, _04583_);
  or (_06449_, _06448_, _03227_);
  or (_06450_, _06449_, _06447_);
  and (_06451_, _06221_, _03227_);
  nor (_06452_, _06451_, _04592_);
  and (_06453_, _06452_, _06450_);
  or (_06454_, _06453_, _05962_);
  and (_06455_, _06454_, _05927_);
  nor (_06456_, _05396_, _06061_);
  and (_06457_, _05396_, _06061_);
  nor (_06458_, _06457_, _06456_);
  and (_06459_, _06458_, _04590_);
  or (_06460_, _06459_, _06455_);
  and (_06461_, _06460_, _05926_);
  and (_06462_, _05960_, _04597_);
  or (_06463_, _06462_, _06461_);
  and (_06464_, _06463_, _05925_);
  and (_06465_, _06456_, _04595_);
  or (_06466_, _06465_, _03238_);
  or (_06467_, _06466_, _06464_);
  and (_06468_, _06221_, _03238_);
  nor (_06469_, _06468_, _04609_);
  and (_06470_, _06469_, _06467_);
  not (_06471_, _04609_);
  nor (_06472_, _05959_, _06471_);
  or (_06473_, _06472_, _04607_);
  or (_06474_, _06473_, _06470_);
  not (_06475_, _03248_);
  nand (_06476_, _06457_, _04607_);
  and (_06477_, _06476_, _06475_);
  and (_06478_, _06477_, _06474_);
  and (_06479_, _04563_, _03066_);
  nor (_06480_, _04839_, _04253_);
  or (_06481_, _06480_, _06479_);
  and (_06482_, _06059_, _03248_);
  or (_06483_, _06482_, _04827_);
  or (_06484_, _06483_, _06481_);
  or (_06485_, _06484_, _06478_);
  not (_06486_, _04618_);
  or (_06487_, _06116_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_06488_, _06125_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_06489_, _06488_, _06124_);
  and (_06490_, _06489_, _06487_);
  or (_06491_, _06125_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_06492_, _06116_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_06493_, _06492_, _06130_);
  and (_06494_, _06493_, _06491_);
  nor (_06495_, _06494_, _06490_);
  nand (_06496_, _06495_, _06107_);
  or (_06497_, _06116_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_06498_, _06125_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_06499_, _06498_, _06124_);
  and (_06500_, _06499_, _06497_);
  or (_06501_, _06125_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_06502_, _06116_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_06503_, _06502_, _06130_);
  and (_06504_, _06503_, _06501_);
  nor (_06505_, _06504_, _06500_);
  nand (_06506_, _06505_, _06136_);
  nand (_06507_, _06506_, _06496_);
  nand (_06508_, _06507_, _06092_);
  or (_06509_, _06116_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_06510_, _06125_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_06511_, _06510_, _06124_);
  nand (_06512_, _06511_, _06509_);
  or (_06513_, _06125_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_06514_, _06116_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_06515_, _06514_, _06130_);
  nand (_06516_, _06515_, _06513_);
  nand (_06517_, _06516_, _06512_);
  and (_06518_, _06517_, _06136_);
  or (_06519_, _06116_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_06520_, _06125_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_06521_, _06520_, _06124_);
  nand (_06522_, _06521_, _06519_);
  or (_06523_, _06125_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_06524_, _06116_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_06525_, _06524_, _06130_);
  nand (_06526_, _06525_, _06523_);
  nand (_06527_, _06526_, _06522_);
  and (_06528_, _06527_, _06107_);
  nor (_06529_, _06528_, _06518_);
  nand (_06530_, _06529_, _06091_);
  and (_06531_, _06530_, _06508_);
  not (_06532_, _06531_);
  or (_06533_, _06116_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_06534_, _06125_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_06535_, _06534_, _06124_);
  and (_06536_, _06535_, _06533_);
  or (_06537_, _06125_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_06538_, _06116_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_06539_, _06538_, _06130_);
  and (_06540_, _06539_, _06537_);
  nor (_06541_, _06540_, _06536_);
  nand (_06542_, _06541_, _06107_);
  or (_06543_, _06116_, \oc8051_golden_model_1.IRAM[9] [1]);
  or (_06544_, _06125_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_06545_, _06544_, _06124_);
  and (_06546_, _06545_, _06543_);
  or (_06547_, _06125_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_06548_, _06116_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_06549_, _06548_, _06130_);
  and (_06550_, _06549_, _06547_);
  nor (_06551_, _06550_, _06546_);
  nand (_06552_, _06551_, _06136_);
  nand (_06553_, _06552_, _06542_);
  nand (_06554_, _06553_, _06092_);
  or (_06555_, _06116_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_06556_, _06125_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_06557_, _06556_, _06124_);
  nand (_06558_, _06557_, _06555_);
  or (_06559_, _06125_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_06560_, _06116_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_06561_, _06560_, _06130_);
  nand (_06562_, _06561_, _06559_);
  nand (_06563_, _06562_, _06558_);
  and (_06564_, _06563_, _06136_);
  or (_06565_, _06116_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_06566_, _06125_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_06567_, _06566_, _06124_);
  nand (_06568_, _06567_, _06565_);
  or (_06569_, _06125_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_06570_, _06116_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_06571_, _06570_, _06130_);
  nand (_06572_, _06571_, _06569_);
  nand (_06573_, _06572_, _06568_);
  and (_06574_, _06573_, _06107_);
  nor (_06575_, _06574_, _06564_);
  nand (_06576_, _06575_, _06091_);
  nand (_06577_, _06576_, _06554_);
  or (_06578_, _06116_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_06579_, _06125_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_06580_, _06579_, _06124_);
  and (_06581_, _06580_, _06578_);
  or (_06582_, _06125_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_06583_, _06116_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_06584_, _06583_, _06130_);
  and (_06585_, _06584_, _06582_);
  nor (_06586_, _06585_, _06581_);
  nand (_06587_, _06586_, _06107_);
  or (_06588_, _06116_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_06589_, _06125_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_06590_, _06589_, _06124_);
  and (_06591_, _06590_, _06588_);
  or (_06592_, _06125_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_06593_, _06116_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_06594_, _06593_, _06130_);
  and (_06595_, _06594_, _06592_);
  nor (_06596_, _06595_, _06591_);
  nand (_06597_, _06596_, _06136_);
  nand (_06598_, _06597_, _06587_);
  nand (_06599_, _06598_, _06092_);
  or (_06600_, _06116_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_06601_, _06125_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_06602_, _06601_, _06124_);
  nand (_06603_, _06602_, _06600_);
  or (_06604_, _06125_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_06605_, _06116_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_06606_, _06605_, _06130_);
  nand (_06607_, _06606_, _06604_);
  nand (_06608_, _06607_, _06603_);
  and (_06609_, _06608_, _06136_);
  or (_06610_, _06116_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_06611_, _06125_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_06612_, _06611_, _06124_);
  nand (_06613_, _06612_, _06610_);
  or (_06614_, _06125_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_06615_, _06116_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_06616_, _06615_, _06130_);
  nand (_06617_, _06616_, _06614_);
  nand (_06618_, _06617_, _06613_);
  and (_06619_, _06618_, _06107_);
  nor (_06620_, _06619_, _06609_);
  nand (_06621_, _06620_, _06091_);
  nand (_06622_, _06621_, _06599_);
  and (_06623_, _06622_, _06577_);
  or (_06624_, _06116_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_06625_, _06125_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_06626_, _06625_, _06124_);
  and (_06627_, _06626_, _06624_);
  or (_06628_, _06125_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_06629_, _06116_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_06630_, _06629_, _06130_);
  and (_06631_, _06630_, _06628_);
  nor (_06632_, _06631_, _06627_);
  nand (_06633_, _06632_, _06107_);
  or (_06634_, _06116_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_06635_, _06125_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_06636_, _06635_, _06124_);
  and (_06637_, _06636_, _06634_);
  or (_06638_, _06125_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_06639_, _06116_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_06640_, _06639_, _06130_);
  and (_06641_, _06640_, _06638_);
  nor (_06642_, _06641_, _06637_);
  nand (_06643_, _06642_, _06136_);
  nand (_06644_, _06643_, _06633_);
  nand (_06645_, _06644_, _06092_);
  or (_06646_, _06116_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_06647_, _06125_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_06648_, _06647_, _06124_);
  nand (_06649_, _06648_, _06646_);
  or (_06650_, _06125_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_06651_, _06116_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_06652_, _06651_, _06130_);
  nand (_06653_, _06652_, _06650_);
  nand (_06654_, _06653_, _06649_);
  and (_06655_, _06654_, _06136_);
  or (_06656_, _06116_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_06657_, _06125_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_06658_, _06657_, _06124_);
  nand (_06659_, _06658_, _06656_);
  or (_06660_, _06125_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_06661_, _06116_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_06662_, _06661_, _06130_);
  nand (_06663_, _06662_, _06660_);
  nand (_06664_, _06663_, _06659_);
  and (_06665_, _06664_, _06107_);
  nor (_06666_, _06665_, _06655_);
  nand (_06667_, _06666_, _06091_);
  nand (_06668_, _06667_, _06645_);
  or (_06669_, _06116_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_06670_, _06125_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_06671_, _06670_, _06124_);
  and (_06672_, _06671_, _06669_);
  or (_06673_, _06125_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_06674_, _06116_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_06675_, _06674_, _06130_);
  and (_06676_, _06675_, _06673_);
  nor (_06677_, _06676_, _06672_);
  nand (_06678_, _06677_, _06107_);
  or (_06679_, _06116_, \oc8051_golden_model_1.IRAM[9] [2]);
  or (_06680_, _06125_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_06681_, _06680_, _06124_);
  and (_06682_, _06681_, _06679_);
  or (_06684_, _06125_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_06685_, _06116_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_06686_, _06685_, _06130_);
  and (_06687_, _06686_, _06684_);
  nor (_06688_, _06687_, _06682_);
  nand (_06689_, _06688_, _06136_);
  nand (_06690_, _06689_, _06678_);
  nand (_06691_, _06690_, _06092_);
  or (_06692_, _06116_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_06693_, _06125_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_06694_, _06693_, _06124_);
  nand (_06695_, _06694_, _06692_);
  or (_06696_, _06125_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_06697_, _06116_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_06698_, _06697_, _06130_);
  nand (_06699_, _06698_, _06696_);
  nand (_06700_, _06699_, _06695_);
  and (_06701_, _06700_, _06136_);
  or (_06702_, _06116_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_06703_, _06125_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_06704_, _06703_, _06124_);
  nand (_06705_, _06704_, _06702_);
  or (_06706_, _06125_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_06707_, _06116_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_06708_, _06707_, _06130_);
  nand (_06709_, _06708_, _06706_);
  nand (_06710_, _06709_, _06705_);
  and (_06711_, _06710_, _06107_);
  nor (_06712_, _06711_, _06701_);
  nand (_06713_, _06712_, _06091_);
  nand (_06714_, _06713_, _06691_);
  and (_06715_, _06714_, _06668_);
  and (_06716_, _06715_, _06623_);
  or (_06717_, _06116_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_06718_, _06125_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_06719_, _06718_, _06124_);
  and (_06720_, _06719_, _06717_);
  or (_06721_, _06125_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06722_, _06116_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_06723_, _06722_, _06130_);
  and (_06724_, _06723_, _06721_);
  nor (_06725_, _06724_, _06720_);
  nand (_06726_, _06725_, _06107_);
  or (_06727_, _06116_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_06728_, _06125_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_06729_, _06728_, _06124_);
  and (_06730_, _06729_, _06727_);
  or (_06731_, _06125_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06732_, _06116_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_06733_, _06732_, _06130_);
  and (_06734_, _06733_, _06731_);
  nor (_06735_, _06734_, _06730_);
  nand (_06736_, _06735_, _06136_);
  nand (_06737_, _06736_, _06726_);
  nand (_06738_, _06737_, _06092_);
  or (_06739_, _06116_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_06740_, _06125_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_06741_, _06740_, _06124_);
  nand (_06742_, _06741_, _06739_);
  or (_06743_, _06125_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_06744_, _06116_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_06745_, _06744_, _06130_);
  nand (_06746_, _06745_, _06743_);
  nand (_06747_, _06746_, _06742_);
  and (_06748_, _06747_, _06136_);
  or (_06749_, _06116_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_06750_, _06125_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_06751_, _06750_, _06124_);
  nand (_06752_, _06751_, _06749_);
  or (_06753_, _06125_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_06754_, _06116_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_06755_, _06754_, _06130_);
  nand (_06756_, _06755_, _06753_);
  nand (_06757_, _06756_, _06752_);
  and (_06758_, _06757_, _06107_);
  nor (_06759_, _06758_, _06748_);
  nand (_06760_, _06759_, _06091_);
  nand (_06761_, _06760_, _06738_);
  or (_06762_, _06116_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_06763_, _06125_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_06764_, _06763_, _06124_);
  and (_06765_, _06764_, _06762_);
  or (_06766_, _06125_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06767_, _06116_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_06768_, _06767_, _06130_);
  and (_06769_, _06768_, _06766_);
  nor (_06770_, _06769_, _06765_);
  nand (_06771_, _06770_, _06107_);
  or (_06772_, _06116_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_06773_, _06125_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_06774_, _06773_, _06124_);
  and (_06775_, _06774_, _06772_);
  or (_06776_, _06125_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06777_, _06116_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_06778_, _06777_, _06130_);
  and (_06779_, _06778_, _06776_);
  nor (_06780_, _06779_, _06775_);
  nand (_06781_, _06780_, _06136_);
  nand (_06782_, _06781_, _06771_);
  nand (_06783_, _06782_, _06092_);
  or (_06784_, _06116_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_06785_, _06125_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_06786_, _06785_, _06124_);
  nand (_06787_, _06786_, _06784_);
  or (_06788_, _06125_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_06789_, _06116_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_06790_, _06789_, _06130_);
  nand (_06791_, _06790_, _06788_);
  nand (_06792_, _06791_, _06787_);
  and (_06793_, _06792_, _06136_);
  or (_06794_, _06116_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_06795_, _06125_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_06796_, _06795_, _06124_);
  nand (_06797_, _06796_, _06794_);
  or (_06798_, _06125_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_06799_, _06116_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_06800_, _06799_, _06130_);
  nand (_06801_, _06800_, _06798_);
  nand (_06802_, _06801_, _06797_);
  and (_06803_, _06802_, _06107_);
  nor (_06804_, _06803_, _06793_);
  nand (_06805_, _06804_, _06091_);
  nand (_06806_, _06805_, _06783_);
  and (_06807_, _06806_, _06761_);
  and (_06808_, _06807_, _06716_);
  and (_06809_, _06808_, _06532_);
  or (_06810_, _06809_, _06171_);
  nand (_06811_, _06809_, _06171_);
  and (_06812_, _06811_, _06810_);
  or (_06813_, _06812_, _06486_);
  nor (_06814_, _06481_, _04781_);
  or (_06815_, _06814_, _06052_);
  and (_06816_, _06815_, _04811_);
  and (_06817_, _06816_, _06813_);
  and (_06818_, _06817_, _06485_);
  and (_06819_, _06185_, _04617_);
  or (_06820_, _06819_, _03686_);
  or (_06821_, _06820_, _06818_);
  and (_06822_, _06821_, _05924_);
  or (_06823_, _06822_, _03243_);
  and (_06824_, _06221_, _03243_);
  nor (_06825_, _06824_, _04624_);
  and (_06826_, _06825_, _06823_);
  not (_06827_, _05913_);
  and (_06828_, _06024_, _04624_);
  or (_06829_, _06828_, _06827_);
  or (_06830_, _06829_, _06826_);
  and (_06831_, _06830_, _05914_);
  or (_06832_, _06831_, _04271_);
  not (_06833_, _04271_);
  not (_06834_, _06171_);
  and (_06835_, _06576_, _06554_);
  and (_06836_, _06621_, _06599_);
  and (_06837_, _06836_, _06835_);
  and (_06838_, _06667_, _06645_);
  and (_06839_, _06713_, _06691_);
  and (_06840_, _06839_, _06838_);
  and (_06841_, _06840_, _06837_);
  and (_06842_, _06760_, _06738_);
  and (_06843_, _06805_, _06783_);
  and (_06844_, _06843_, _06842_);
  and (_06845_, _06844_, _06841_);
  and (_06846_, _06845_, _06531_);
  nor (_06847_, _06846_, _06834_);
  and (_06848_, _06846_, _06834_);
  or (_06849_, _06848_, _06847_);
  or (_06850_, _06849_, _06833_);
  and (_06851_, _06850_, _04805_);
  and (_06852_, _06851_, _06832_);
  or (_06853_, _06852_, _05896_);
  and (_06854_, _06853_, _05227_);
  or (_06855_, _06854_, _05236_);
  and (_06856_, _06855_, _05226_);
  not (_06857_, \oc8051_golden_model_1.PC [15]);
  and (_06858_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_06859_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_06860_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_06861_, _06860_, _06859_);
  and (_06862_, _06861_, _05920_);
  and (_06863_, _06862_, _06858_);
  and (_06864_, _06863_, \oc8051_golden_model_1.PC [14]);
  and (_06865_, _06864_, _06857_);
  nor (_06866_, _06864_, _06857_);
  or (_06867_, _06866_, _06865_);
  and (_06868_, _06867_, _03686_);
  and (_06869_, _06861_, _06057_);
  and (_06870_, _06869_, _06858_);
  and (_06871_, _06870_, \oc8051_golden_model_1.PC [14]);
  and (_06872_, _06871_, _06857_);
  nor (_06873_, _06871_, _06857_);
  or (_06874_, _06873_, _06872_);
  not (_06875_, _06874_);
  nor (_06876_, _06875_, _03686_);
  or (_06877_, _06876_, _06868_);
  and (_06878_, _06877_, _05221_);
  and (_06879_, _06878_, _05224_);
  or (_40744_, _06879_, _06856_);
  not (_06880_, \oc8051_golden_model_1.B [7]);
  nor (_06881_, _43227_, _06880_);
  nor (_06882_, _05379_, _06880_);
  not (_06883_, _05379_);
  nor (_06884_, _06883_, _05289_);
  or (_06885_, _06884_, _06882_);
  nor (_06886_, _03584_, _03574_);
  and (_06887_, _06886_, _05080_);
  nor (_06888_, _06887_, _03271_);
  nor (_06889_, _06888_, _04131_);
  or (_06890_, _06889_, _06885_);
  nor (_06891_, _05992_, _06880_);
  and (_06892_, _06038_, _05992_);
  or (_06893_, _06892_, _06891_);
  and (_06894_, _06893_, _03511_);
  and (_06895_, _06185_, _05379_);
  or (_06896_, _06895_, _06882_);
  or (_06897_, _06896_, _04515_);
  and (_06898_, _05379_, \oc8051_golden_model_1.ACC [7]);
  or (_06899_, _06898_, _06882_);
  and (_06900_, _06899_, _04499_);
  nor (_06901_, _04499_, _06880_);
  or (_06902_, _06901_, _03599_);
  or (_06903_, _06902_, _06900_);
  and (_06904_, _06903_, _03516_);
  and (_06905_, _06904_, _06897_);
  and (_06906_, _06042_, _05992_);
  or (_06907_, _06906_, _06891_);
  and (_06908_, _06907_, _03515_);
  or (_06909_, _06908_, _03597_);
  or (_06910_, _06909_, _06905_);
  or (_06911_, _06885_, _04524_);
  and (_06912_, _06911_, _06910_);
  or (_06913_, _06912_, _03603_);
  or (_06914_, _06899_, _03611_);
  and (_06915_, _06914_, _03512_);
  and (_06916_, _06915_, _06913_);
  or (_06917_, _06916_, _06894_);
  and (_06918_, _06917_, _03505_);
  and (_06919_, _03675_, _03566_);
  or (_06920_, _06891_, _06216_);
  and (_06921_, _06920_, _03504_);
  and (_06922_, _06921_, _06907_);
  or (_06923_, _06922_, _06919_);
  or (_06924_, _06923_, _06918_);
  not (_06925_, _06919_);
  and (_06926_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_06927_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_06928_, _06927_, _06926_);
  and (_06929_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_06930_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_06931_, _06930_, _06929_);
  and (_06932_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_06933_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and (_06934_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor (_06935_, _06934_, _06933_);
  nor (_06936_, _06935_, _06931_);
  and (_06937_, _06936_, _06932_);
  nor (_06938_, _06937_, _06931_);
  and (_06939_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_06940_, _06939_, _06933_);
  and (_06941_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_06942_, _06941_, _06929_);
  nor (_06943_, _06942_, _06940_);
  not (_06944_, _06943_);
  nor (_06945_, _06944_, _06938_);
  and (_06946_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_06947_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_06948_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_06949_, _06948_, _06947_);
  nor (_06950_, _06948_, _06947_);
  nor (_06951_, _06950_, _06949_);
  and (_06952_, _06951_, _06946_);
  nor (_06953_, _06951_, _06946_);
  nor (_06954_, _06953_, _06952_);
  and (_06955_, _06944_, _06938_);
  nor (_06956_, _06955_, _06945_);
  and (_06957_, _06956_, _06954_);
  nor (_06958_, _06957_, _06945_);
  not (_06959_, _06933_);
  and (_06960_, _06939_, _06959_);
  and (_06961_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_06962_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_06963_, _06962_, _06947_);
  and (_06964_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_06965_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_06966_, _06965_, _06964_);
  nor (_06967_, _06966_, _06963_);
  and (_06968_, _06967_, _06961_);
  nor (_06969_, _06967_, _06961_);
  nor (_06970_, _06969_, _06968_);
  and (_06971_, _06970_, _06960_);
  nor (_06972_, _06970_, _06960_);
  nor (_06973_, _06972_, _06971_);
  not (_06974_, _06973_);
  nor (_06975_, _06974_, _06958_);
  and (_06976_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_06977_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_06978_, _06977_, _06976_);
  nor (_06979_, _06952_, _06949_);
  and (_06980_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_06981_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_06982_, _06981_, _06980_);
  nor (_06983_, _06981_, _06980_);
  nor (_06984_, _06983_, _06982_);
  not (_06985_, _06984_);
  nor (_06986_, _06985_, _06979_);
  and (_06987_, _06985_, _06979_);
  nor (_06988_, _06987_, _06986_);
  and (_06989_, _06988_, _06978_);
  nor (_06990_, _06988_, _06978_);
  nor (_06991_, _06990_, _06989_);
  and (_06992_, _06974_, _06958_);
  nor (_06993_, _06992_, _06975_);
  and (_06994_, _06993_, _06991_);
  nor (_06995_, _06994_, _06975_);
  nor (_06996_, _06968_, _06963_);
  and (_06997_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_06998_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_06999_, _06998_, _06997_);
  nor (_07000_, _06998_, _06997_);
  nor (_07001_, _07000_, _06999_);
  not (_07002_, _07001_);
  nor (_07003_, _07002_, _06996_);
  and (_07004_, _07002_, _06996_);
  nor (_07005_, _07004_, _07003_);
  and (_07006_, _07005_, _06982_);
  nor (_07007_, _07005_, _06982_);
  nor (_07008_, _07007_, _07006_);
  nor (_07009_, _06971_, _06940_);
  and (_07010_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_07011_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_07012_, _07011_, _06962_);
  nor (_07013_, _07011_, _06962_);
  nor (_07014_, _07013_, _07012_);
  and (_07015_, _07014_, _07010_);
  nor (_07016_, _07014_, _07010_);
  nor (_07017_, _07016_, _07015_);
  not (_07018_, _07017_);
  nor (_07019_, _07018_, _07009_);
  and (_07020_, _07018_, _07009_);
  nor (_07021_, _07020_, _07019_);
  and (_07022_, _07021_, _07008_);
  nor (_07023_, _07021_, _07008_);
  nor (_07024_, _07023_, _07022_);
  not (_07025_, _07024_);
  nor (_07026_, _07025_, _06995_);
  nor (_07027_, _06989_, _06986_);
  not (_07028_, _07027_);
  and (_07029_, _07025_, _06995_);
  nor (_07030_, _07029_, _07026_);
  and (_07031_, _07030_, _07028_);
  nor (_07032_, _07031_, _07026_);
  nor (_07033_, _07006_, _07003_);
  not (_07034_, _07033_);
  nor (_07035_, _07022_, _07019_);
  not (_07036_, _07035_);
  and (_07037_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_07038_, _07037_, _06962_);
  and (_07039_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_07040_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_07041_, _07040_, _07039_);
  nor (_07042_, _07041_, _07038_);
  nor (_07043_, _07015_, _07012_);
  and (_07044_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_07045_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_07046_, _07045_, _07044_);
  nor (_07047_, _07045_, _07044_);
  nor (_07048_, _07047_, _07046_);
  not (_07049_, _07048_);
  nor (_07050_, _07049_, _07043_);
  and (_07051_, _07049_, _07043_);
  nor (_07052_, _07051_, _07050_);
  and (_07053_, _07052_, _06999_);
  nor (_07054_, _07052_, _06999_);
  nor (_07055_, _07054_, _07053_);
  and (_07056_, _07055_, _07042_);
  nor (_07057_, _07055_, _07042_);
  nor (_07058_, _07057_, _07056_);
  and (_07059_, _07058_, _07036_);
  nor (_07060_, _07058_, _07036_);
  nor (_07061_, _07060_, _07059_);
  and (_07062_, _07061_, _07034_);
  nor (_07063_, _07061_, _07034_);
  nor (_07064_, _07063_, _07062_);
  not (_07065_, _07064_);
  nor (_07066_, _07065_, _07032_);
  nor (_07067_, _07062_, _07059_);
  nor (_07068_, _07053_, _07050_);
  not (_07069_, _07068_);
  and (_07070_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_07071_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_07072_, _07071_, _07070_);
  nor (_07073_, _07071_, _07070_);
  nor (_07074_, _07073_, _07072_);
  and (_07075_, _07074_, _07038_);
  nor (_07076_, _07074_, _07038_);
  nor (_07077_, _07076_, _07075_);
  and (_07078_, _07077_, _07046_);
  nor (_07079_, _07077_, _07046_);
  nor (_07080_, _07079_, _07078_);
  and (_07081_, _07080_, _07037_);
  nor (_07082_, _07080_, _07037_);
  nor (_07083_, _07082_, _07081_);
  and (_07084_, _07083_, _07056_);
  nor (_07085_, _07083_, _07056_);
  nor (_07086_, _07085_, _07084_);
  and (_07087_, _07086_, _07069_);
  nor (_07088_, _07086_, _07069_);
  nor (_07089_, _07088_, _07087_);
  not (_07090_, _07089_);
  nor (_07091_, _07090_, _07067_);
  and (_07092_, _07090_, _07067_);
  nor (_07093_, _07092_, _07091_);
  and (_07094_, _07093_, _07066_);
  nor (_07095_, _07087_, _07084_);
  nor (_07096_, _07078_, _07075_);
  not (_07097_, _07096_);
  nor (_07098_, _06927_, _06926_);
  nor (_07099_, _07098_, _06928_);
  and (_07100_, _07099_, _07072_);
  nor (_07101_, _07099_, _07072_);
  nor (_07102_, _07101_, _07100_);
  and (_07103_, _07102_, _07081_);
  nor (_07104_, _07102_, _07081_);
  nor (_07105_, _07104_, _07103_);
  and (_07106_, _07105_, _07097_);
  nor (_07107_, _07105_, _07097_);
  nor (_07108_, _07107_, _07106_);
  not (_07109_, _07108_);
  nor (_07110_, _07109_, _07095_);
  and (_07111_, _07109_, _07095_);
  nor (_07112_, _07111_, _07110_);
  and (_07113_, _07112_, _07091_);
  nor (_07114_, _07112_, _07091_);
  nor (_07115_, _07114_, _07113_);
  and (_07116_, _07115_, _07094_);
  nor (_07117_, _07115_, _07094_);
  and (_07118_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_07119_, _07118_, _06933_);
  and (_07120_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_07121_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_07122_, _07121_, _06930_);
  nor (_07123_, _07122_, _07119_);
  and (_07124_, _07123_, _07120_);
  nor (_07125_, _07124_, _07119_);
  not (_07126_, _07125_);
  nor (_07127_, _06936_, _06932_);
  nor (_07128_, _07127_, _06937_);
  and (_07129_, _07128_, _07126_);
  and (_07130_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_07131_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_07132_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_07133_, _07132_, _07131_);
  nor (_07134_, _07132_, _07131_);
  nor (_07135_, _07134_, _07133_);
  and (_07136_, _07135_, _07130_);
  nor (_07137_, _07135_, _07130_);
  nor (_07138_, _07137_, _07136_);
  nor (_07139_, _07128_, _07126_);
  nor (_07140_, _07139_, _07129_);
  and (_07141_, _07140_, _07138_);
  nor (_07142_, _07141_, _07129_);
  nor (_07143_, _06956_, _06954_);
  nor (_07144_, _07143_, _06957_);
  not (_07145_, _07144_);
  nor (_07146_, _07145_, _07142_);
  and (_07147_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_07148_, _07147_, _06977_);
  nor (_07149_, _07136_, _07133_);
  nor (_07150_, _06977_, _06976_);
  nor (_07151_, _07150_, _06978_);
  not (_07152_, _07151_);
  nor (_07153_, _07152_, _07149_);
  and (_07154_, _07152_, _07149_);
  nor (_07155_, _07154_, _07153_);
  and (_07156_, _07155_, _07148_);
  nor (_07157_, _07155_, _07148_);
  nor (_07158_, _07157_, _07156_);
  and (_07159_, _07145_, _07142_);
  nor (_07160_, _07159_, _07146_);
  and (_07161_, _07160_, _07158_);
  nor (_07162_, _07161_, _07146_);
  nor (_07163_, _06993_, _06991_);
  nor (_07164_, _07163_, _06994_);
  not (_07165_, _07164_);
  nor (_07166_, _07165_, _07162_);
  nor (_07167_, _07156_, _07153_);
  not (_07168_, _07167_);
  and (_07169_, _07165_, _07162_);
  nor (_07170_, _07169_, _07166_);
  and (_07171_, _07170_, _07168_);
  nor (_07172_, _07171_, _07166_);
  nor (_07173_, _07030_, _07028_);
  nor (_07174_, _07173_, _07031_);
  not (_07175_, _07174_);
  nor (_07176_, _07175_, _07172_);
  and (_07177_, _07065_, _07032_);
  nor (_07178_, _07177_, _07066_);
  and (_07179_, _07178_, _07176_);
  nor (_07180_, _07093_, _07066_);
  nor (_07181_, _07180_, _07094_);
  and (_07182_, _07181_, _07179_);
  and (_07183_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_07184_, _07183_, _07118_);
  and (_07185_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_07186_, _07183_, _07118_);
  nor (_07187_, _07186_, _07184_);
  and (_07188_, _07187_, _07185_);
  nor (_07189_, _07188_, _07184_);
  not (_07190_, _07189_);
  nor (_07191_, _07123_, _07120_);
  nor (_07192_, _07191_, _07124_);
  and (_07193_, _07192_, _07190_);
  and (_07194_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_07195_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_07196_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_07197_, _07196_, _07195_);
  nor (_07198_, _07196_, _07195_);
  nor (_07199_, _07198_, _07197_);
  and (_07200_, _07199_, _07194_);
  nor (_07201_, _07199_, _07194_);
  nor (_07202_, _07201_, _07200_);
  nor (_07203_, _07192_, _07190_);
  nor (_07204_, _07203_, _07193_);
  and (_07205_, _07204_, _07202_);
  nor (_07206_, _07205_, _07193_);
  not (_07207_, _07206_);
  nor (_07208_, _07140_, _07138_);
  nor (_07209_, _07208_, _07141_);
  and (_07210_, _07209_, _07207_);
  nor (_07211_, _07200_, _07197_);
  and (_07212_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_07213_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_07214_, _07213_, _07212_);
  nor (_07215_, _07214_, _07148_);
  not (_07216_, _07215_);
  nor (_07217_, _07216_, _07211_);
  and (_07218_, _07216_, _07211_);
  nor (_07219_, _07218_, _07217_);
  nor (_07220_, _07209_, _07207_);
  nor (_07221_, _07220_, _07210_);
  and (_07222_, _07221_, _07219_);
  nor (_07223_, _07222_, _07210_);
  nor (_07224_, _07160_, _07158_);
  nor (_07225_, _07224_, _07161_);
  not (_07226_, _07225_);
  nor (_07227_, _07226_, _07223_);
  and (_07228_, _07226_, _07223_);
  nor (_07229_, _07228_, _07227_);
  and (_07230_, _07229_, _07217_);
  nor (_07231_, _07230_, _07227_);
  nor (_07232_, _07170_, _07168_);
  nor (_07233_, _07232_, _07171_);
  not (_07234_, _07233_);
  nor (_07235_, _07234_, _07231_);
  and (_07236_, _07175_, _07172_);
  nor (_07237_, _07236_, _07176_);
  and (_07238_, _07237_, _07235_);
  nor (_07239_, _07178_, _07176_);
  nor (_07240_, _07239_, _07179_);
  and (_07241_, _07240_, _07238_);
  nor (_07242_, _07240_, _07238_);
  nor (_07243_, _07242_, _07241_);
  and (_07244_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_07245_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_07246_, _07245_, _07244_);
  and (_07247_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_07248_, _07245_, _07244_);
  nor (_07249_, _07248_, _07246_);
  and (_07250_, _07249_, _07247_);
  nor (_07251_, _07250_, _07246_);
  not (_07252_, _07251_);
  nor (_07253_, _07187_, _07185_);
  nor (_07254_, _07253_, _07188_);
  and (_07255_, _07254_, _07252_);
  and (_07256_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_07257_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_07258_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_07259_, _07258_, _07257_);
  nor (_07260_, _07258_, _07257_);
  nor (_07261_, _07260_, _07259_);
  and (_07262_, _07261_, _07256_);
  nor (_07263_, _07261_, _07256_);
  nor (_07264_, _07263_, _07262_);
  nor (_07265_, _07254_, _07252_);
  nor (_07266_, _07265_, _07255_);
  and (_07267_, _07266_, _07264_);
  nor (_07268_, _07267_, _07255_);
  not (_07269_, _07268_);
  nor (_07270_, _07204_, _07202_);
  nor (_07271_, _07270_, _07205_);
  and (_07272_, _07271_, _07269_);
  not (_07273_, _07147_);
  nor (_07274_, _07262_, _07259_);
  nor (_07275_, _07274_, _07273_);
  and (_07276_, _07274_, _07273_);
  nor (_07277_, _07276_, _07275_);
  nor (_07278_, _07271_, _07269_);
  nor (_07279_, _07278_, _07272_);
  and (_07280_, _07279_, _07277_);
  nor (_07281_, _07280_, _07272_);
  not (_07282_, _07281_);
  nor (_07283_, _07221_, _07219_);
  nor (_07284_, _07283_, _07222_);
  and (_07285_, _07284_, _07282_);
  nor (_07286_, _07284_, _07282_);
  nor (_07287_, _07286_, _07285_);
  and (_07288_, _07287_, _07275_);
  nor (_07289_, _07288_, _07285_);
  nor (_07290_, _07229_, _07217_);
  nor (_07291_, _07290_, _07230_);
  not (_07292_, _07291_);
  nor (_07293_, _07292_, _07289_);
  and (_07294_, _07234_, _07231_);
  nor (_07295_, _07294_, _07235_);
  and (_07296_, _07295_, _07293_);
  nor (_07297_, _07237_, _07235_);
  nor (_07298_, _07297_, _07238_);
  and (_07299_, _07298_, _07296_);
  nor (_07300_, _07298_, _07296_);
  nor (_07301_, _07300_, _07299_);
  and (_07302_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_07303_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_07304_, _07303_, _07302_);
  and (_07305_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07306_, _07303_, _07302_);
  nor (_07307_, _07306_, _07304_);
  and (_07308_, _07307_, _07305_);
  nor (_07309_, _07308_, _07304_);
  not (_07310_, _07309_);
  nor (_07311_, _07249_, _07247_);
  nor (_07312_, _07311_, _07250_);
  and (_07313_, _07312_, _07310_);
  and (_07314_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_07315_, _07314_, _07258_);
  and (_07316_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_07317_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_07318_, _07317_, _07316_);
  nor (_07319_, _07318_, _07315_);
  nor (_07320_, _07312_, _07310_);
  nor (_07321_, _07320_, _07313_);
  and (_07322_, _07321_, _07319_);
  nor (_07323_, _07322_, _07313_);
  not (_07324_, _07323_);
  nor (_07325_, _07266_, _07264_);
  nor (_07326_, _07325_, _07267_);
  and (_07327_, _07326_, _07324_);
  nor (_07328_, _07326_, _07324_);
  nor (_07329_, _07328_, _07327_);
  and (_07330_, _07329_, _07315_);
  nor (_07331_, _07330_, _07327_);
  not (_07332_, _07331_);
  nor (_07333_, _07279_, _07277_);
  nor (_07334_, _07333_, _07280_);
  and (_07335_, _07334_, _07332_);
  nor (_07336_, _07287_, _07275_);
  nor (_07337_, _07336_, _07288_);
  and (_07338_, _07337_, _07335_);
  and (_07339_, _07292_, _07289_);
  nor (_07340_, _07339_, _07293_);
  and (_07341_, _07340_, _07338_);
  nor (_07342_, _07295_, _07293_);
  nor (_07343_, _07342_, _07296_);
  and (_07344_, _07343_, _07341_);
  nor (_07345_, _07343_, _07341_);
  nor (_07346_, _07345_, _07344_);
  and (_07347_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_07348_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_07349_, _07348_, _07347_);
  and (_07350_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_07351_, _07348_, _07347_);
  nor (_07352_, _07351_, _07349_);
  and (_07353_, _07352_, _07350_);
  nor (_07354_, _07353_, _07349_);
  not (_07355_, _07354_);
  nor (_07356_, _07307_, _07305_);
  nor (_07357_, _07356_, _07308_);
  and (_07358_, _07357_, _07355_);
  nor (_07359_, _07357_, _07355_);
  nor (_07360_, _07359_, _07358_);
  and (_07361_, _07360_, _07314_);
  nor (_07362_, _07361_, _07358_);
  not (_07363_, _07362_);
  nor (_07364_, _07321_, _07319_);
  nor (_07365_, _07364_, _07322_);
  and (_07366_, _07365_, _07363_);
  nor (_07367_, _07329_, _07315_);
  nor (_07368_, _07367_, _07330_);
  and (_07369_, _07368_, _07366_);
  nor (_07370_, _07334_, _07332_);
  nor (_07371_, _07370_, _07335_);
  and (_07372_, _07371_, _07369_);
  nor (_07373_, _07337_, _07335_);
  nor (_07374_, _07373_, _07338_);
  and (_07375_, _07374_, _07372_);
  nor (_07376_, _07340_, _07338_);
  nor (_07377_, _07376_, _07341_);
  and (_07378_, _07377_, _07375_);
  and (_07379_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_07380_, _07379_, _07348_);
  nor (_07381_, _07352_, _07350_);
  nor (_07382_, _07381_, _07353_);
  and (_07383_, _07382_, _07380_);
  nor (_07384_, _07360_, _07314_);
  nor (_07385_, _07384_, _07361_);
  and (_07386_, _07385_, _07383_);
  nor (_07387_, _07365_, _07363_);
  nor (_07388_, _07387_, _07366_);
  and (_07389_, _07388_, _07386_);
  nor (_07390_, _07368_, _07366_);
  nor (_07391_, _07390_, _07369_);
  and (_07392_, _07391_, _07389_);
  nor (_07393_, _07371_, _07369_);
  nor (_07394_, _07393_, _07372_);
  and (_07395_, _07394_, _07392_);
  nor (_07396_, _07374_, _07372_);
  nor (_07397_, _07396_, _07375_);
  and (_07398_, _07397_, _07395_);
  nor (_07399_, _07377_, _07375_);
  nor (_07400_, _07399_, _07378_);
  and (_07401_, _07400_, _07398_);
  nor (_07402_, _07401_, _07378_);
  not (_07403_, _07402_);
  and (_07404_, _07403_, _07346_);
  nor (_07405_, _07404_, _07344_);
  not (_07406_, _07405_);
  and (_07407_, _07406_, _07301_);
  nor (_07408_, _07407_, _07299_);
  not (_07409_, _07408_);
  and (_07410_, _07409_, _07243_);
  nor (_07411_, _07410_, _07241_);
  not (_07412_, _07411_);
  nor (_07413_, _07181_, _07179_);
  nor (_07414_, _07413_, _07182_);
  and (_07415_, _07414_, _07412_);
  nor (_07416_, _07415_, _07182_);
  nor (_07417_, _07416_, _07117_);
  or (_07418_, _07417_, _07116_);
  and (_07419_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_07420_, _07419_);
  nor (_07421_, _07420_, _07071_);
  nor (_07422_, _07421_, _07100_);
  nor (_07423_, _07106_, _07103_);
  nor (_07424_, _07423_, _07422_);
  and (_07425_, _07423_, _07422_);
  nor (_07426_, _07425_, _07424_);
  nor (_07427_, _07113_, _07110_);
  and (_07428_, _07427_, _07426_);
  nor (_07429_, _07427_, _07426_);
  or (_07430_, _07429_, _07428_);
  and (_07431_, _07430_, _07418_);
  and (_07432_, _07426_, _07113_);
  and (_07433_, _07426_, _07110_);
  or (_07434_, _07433_, _07424_);
  or (_07435_, _07434_, _07432_);
  or (_07436_, _07435_, _07431_);
  or (_07437_, _07436_, _06928_);
  or (_07438_, _07437_, _06925_);
  and (_07439_, _07438_, _03501_);
  and (_07440_, _07439_, _06924_);
  not (_07441_, _06889_);
  not (_07442_, _05992_);
  nor (_07443_, _06026_, _07442_);
  or (_07444_, _07443_, _06891_);
  and (_07445_, _07444_, _03500_);
  or (_07446_, _07445_, _07441_);
  or (_07447_, _07446_, _07440_);
  and (_07448_, _07447_, _06890_);
  or (_07449_, _07448_, _05969_);
  and (_07450_, _06171_, _05379_);
  or (_07451_, _06882_, _05970_);
  or (_07452_, _07451_, _07450_);
  and (_07453_, _07452_, _03275_);
  and (_07454_, _07453_, _07449_);
  and (_07455_, _03675_, _03219_);
  nor (_07456_, _06443_, _06883_);
  or (_07457_, _07456_, _06882_);
  and (_07458_, _07457_, _03644_);
  or (_07459_, _07458_, _07455_);
  or (_07460_, _07459_, _07454_);
  not (_07461_, \oc8051_golden_model_1.B [1]);
  nor (_07462_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_07463_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_07464_, _07463_, _07462_);
  and (_07465_, _07464_, _07461_);
  nor (_07466_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_07467_, \oc8051_golden_model_1.B [0]);
  and (_07468_, _07467_, \oc8051_golden_model_1.ACC [7]);
  and (_07469_, _07468_, _07466_);
  and (_07470_, _07469_, _07465_);
  or (_07471_, _07467_, \oc8051_golden_model_1.ACC [7]);
  and (_07472_, _07471_, _07466_);
  and (_07473_, _07472_, _07465_);
  or (_07474_, _07473_, _06061_);
  not (_07475_, \oc8051_golden_model_1.B [2]);
  not (_07476_, \oc8051_golden_model_1.B [3]);
  not (_07477_, \oc8051_golden_model_1.B [4]);
  not (_07478_, \oc8051_golden_model_1.B [5]);
  nor (_07479_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_07480_, _07479_, _07478_);
  and (_07481_, _07480_, _07477_);
  and (_07482_, _07481_, _07476_);
  and (_07483_, _07482_, _07475_);
  not (_07484_, \oc8051_golden_model_1.ACC [6]);
  and (_07485_, \oc8051_golden_model_1.B [0], _07484_);
  nor (_07486_, _07485_, _06061_);
  nor (_07487_, _07486_, _07461_);
  not (_07488_, _07487_);
  and (_07489_, _07488_, _07483_);
  nor (_07490_, _07489_, _07474_);
  nor (_07491_, _07490_, _07470_);
  and (_07492_, _07489_, \oc8051_golden_model_1.B [0]);
  nor (_07493_, _07492_, _07484_);
  and (_07494_, _07493_, _07461_);
  nor (_07495_, _07493_, _07461_);
  nor (_07496_, _07495_, _07494_);
  nor (_07497_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_07498_, _07497_, _07118_);
  nor (_07499_, _07498_, \oc8051_golden_model_1.ACC [4]);
  nor (_07500_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_07501_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_07502_, _07501_, _07467_);
  nor (_07503_, _07502_, _07500_);
  nor (_07504_, _07503_, _07499_);
  not (_07505_, _07504_);
  and (_07506_, _07505_, _07496_);
  nor (_07507_, _07491_, \oc8051_golden_model_1.B [2]);
  nor (_07508_, _07507_, _07494_);
  not (_07509_, _07508_);
  nor (_07510_, _07509_, _07506_);
  and (_07511_, \oc8051_golden_model_1.B [2], _06061_);
  nor (_07512_, _07511_, \oc8051_golden_model_1.B [7]);
  and (_07513_, _07512_, _07464_);
  not (_07514_, _07513_);
  nor (_07515_, _07514_, _07510_);
  nor (_07516_, _07515_, _07491_);
  nor (_07517_, _07516_, _07470_);
  and (_07518_, _07481_, \oc8051_golden_model_1.ACC [7]);
  nor (_07519_, _07518_, _07482_);
  nor (_07520_, _07505_, _07496_);
  nor (_07521_, _07520_, _07506_);
  not (_07522_, _07521_);
  and (_07523_, _07522_, _07515_);
  nor (_07524_, _07515_, _07493_);
  nor (_07525_, _07524_, _07523_);
  and (_07526_, _07525_, _07475_);
  nor (_07527_, _07525_, _07475_);
  nor (_07528_, _07527_, _07526_);
  not (_07529_, _07528_);
  not (_07530_, \oc8051_golden_model_1.ACC [5]);
  nor (_07531_, _07515_, _07530_);
  and (_07532_, _07515_, _07498_);
  or (_07533_, _07532_, _07531_);
  and (_07534_, _07533_, _07461_);
  nor (_07535_, _07533_, _07461_);
  not (_07536_, \oc8051_golden_model_1.ACC [4]);
  and (_07537_, \oc8051_golden_model_1.B [0], _07536_);
  nor (_07538_, _07537_, _07535_);
  nor (_07539_, _07538_, _07534_);
  nor (_07540_, _07539_, _07529_);
  nor (_07541_, _07517_, \oc8051_golden_model_1.B [3]);
  nor (_07542_, _07541_, _07526_);
  not (_07543_, _07542_);
  nor (_07544_, _07543_, _07540_);
  nor (_07545_, _07544_, _07519_);
  nor (_07546_, _07545_, _07517_);
  nor (_07547_, _07546_, _07470_);
  nor (_07548_, _07547_, \oc8051_golden_model_1.B [4]);
  not (_07549_, _07545_);
  and (_07550_, _07539_, _07529_);
  nor (_07551_, _07550_, _07540_);
  nor (_07552_, _07551_, _07549_);
  nor (_07553_, _07545_, _07525_);
  nor (_07554_, _07553_, _07552_);
  and (_07555_, _07554_, _07476_);
  nor (_07556_, _07554_, _07476_);
  nor (_07557_, _07556_, _07555_);
  not (_07558_, _07557_);
  nor (_07559_, _07545_, _07533_);
  nor (_07560_, _07535_, _07534_);
  and (_07561_, _07560_, _07537_);
  nor (_07562_, _07560_, _07537_);
  nor (_07563_, _07562_, _07561_);
  and (_07564_, _07563_, _07545_);
  or (_07565_, _07564_, _07559_);
  nor (_07566_, _07565_, \oc8051_golden_model_1.B [2]);
  and (_07567_, _07565_, \oc8051_golden_model_1.B [2]);
  nor (_07568_, _07545_, _07536_);
  nor (_07569_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_07570_, _07569_, _07244_);
  and (_07571_, _07545_, _07570_);
  or (_07572_, _07571_, _07568_);
  and (_07573_, _07572_, _07461_);
  nor (_07574_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_07575_, _07574_, _07302_);
  nor (_07576_, _07575_, \oc8051_golden_model_1.ACC [2]);
  nor (_07577_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_07578_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_07579_, _07578_, _07467_);
  nor (_07580_, _07579_, _07577_);
  nor (_07581_, _07580_, _07576_);
  not (_07582_, _07581_);
  nor (_07583_, _07572_, _07461_);
  nor (_07584_, _07583_, _07573_);
  and (_07585_, _07584_, _07582_);
  nor (_07586_, _07585_, _07573_);
  nor (_07587_, _07586_, _07567_);
  nor (_07588_, _07587_, _07566_);
  nor (_07589_, _07588_, _07558_);
  or (_07590_, _07589_, _07555_);
  nor (_07591_, _07590_, _07548_);
  and (_07592_, _07480_, \oc8051_golden_model_1.ACC [7]);
  or (_07593_, _07592_, _07481_);
  not (_07594_, _07593_);
  nor (_07595_, _07594_, _07591_);
  nor (_07596_, _07595_, _07547_);
  nor (_07597_, _07596_, _07470_);
  and (_07598_, _07479_, \oc8051_golden_model_1.ACC [7]);
  nor (_07599_, _07598_, _07480_);
  nor (_07600_, _07597_, \oc8051_golden_model_1.B [5]);
  and (_07601_, _07588_, _07558_);
  nor (_07602_, _07601_, _07589_);
  not (_07603_, _07602_);
  and (_07604_, _07603_, _07595_);
  nor (_07605_, _07595_, _07554_);
  nor (_07606_, _07605_, _07604_);
  and (_07607_, _07606_, _07477_);
  nor (_07608_, _07606_, _07477_);
  nor (_07609_, _07608_, _07607_);
  not (_07610_, _07609_);
  nor (_07611_, _07595_, _07565_);
  nor (_07612_, _07567_, _07566_);
  and (_07613_, _07612_, _07586_);
  nor (_07614_, _07612_, _07586_);
  nor (_07615_, _07614_, _07613_);
  not (_07616_, _07615_);
  and (_07617_, _07616_, _07595_);
  nor (_07618_, _07617_, _07611_);
  nor (_07619_, _07618_, \oc8051_golden_model_1.B [3]);
  and (_07620_, _07618_, \oc8051_golden_model_1.B [3]);
  nor (_07621_, _07584_, _07582_);
  nor (_07622_, _07621_, _07585_);
  not (_07623_, _07622_);
  and (_07624_, _07623_, _07595_);
  nor (_07625_, _07595_, _07572_);
  nor (_07626_, _07625_, _07624_);
  and (_07627_, _07626_, _07475_);
  not (_07628_, \oc8051_golden_model_1.ACC [3]);
  nor (_07629_, _07595_, _07628_);
  and (_07630_, _07595_, _07575_);
  or (_07631_, _07630_, _07629_);
  and (_07632_, _07631_, _07461_);
  nor (_07633_, _07631_, _07461_);
  not (_07634_, \oc8051_golden_model_1.ACC [2]);
  and (_07635_, \oc8051_golden_model_1.B [0], _07634_);
  nor (_07636_, _07635_, _07633_);
  nor (_07637_, _07636_, _07632_);
  nor (_07638_, _07626_, _07475_);
  nor (_07639_, _07638_, _07627_);
  not (_07640_, _07639_);
  nor (_07641_, _07640_, _07637_);
  nor (_07642_, _07641_, _07627_);
  nor (_07643_, _07642_, _07620_);
  nor (_07644_, _07643_, _07619_);
  nor (_07645_, _07644_, _07610_);
  or (_07646_, _07645_, _07607_);
  nor (_07647_, _07646_, _07600_);
  nor (_07648_, _07647_, _07599_);
  nor (_07649_, _07648_, _07597_);
  not (_07650_, _07648_);
  and (_07651_, _07644_, _07610_);
  nor (_07652_, _07651_, _07645_);
  nor (_07653_, _07652_, _07650_);
  nor (_07654_, _07648_, _07606_);
  nor (_07655_, _07654_, _07653_);
  and (_07656_, _07655_, _07478_);
  nor (_07657_, _07655_, _07478_);
  nor (_07658_, _07657_, _07656_);
  not (_07659_, _07658_);
  nor (_07660_, _07648_, _07618_);
  nor (_07661_, _07620_, _07619_);
  nor (_07662_, _07661_, _07642_);
  and (_07663_, _07661_, _07642_);
  or (_07664_, _07663_, _07662_);
  and (_07665_, _07664_, _07648_);
  or (_07666_, _07665_, _07660_);
  and (_07667_, _07666_, _07477_);
  nor (_07668_, _07666_, _07477_);
  and (_07669_, _07640_, _07637_);
  nor (_07670_, _07669_, _07641_);
  nor (_07671_, _07670_, _07650_);
  nor (_07672_, _07648_, _07626_);
  nor (_07673_, _07672_, _07671_);
  and (_07674_, _07673_, _07476_);
  nor (_07675_, _07633_, _07632_);
  nor (_07676_, _07675_, _07635_);
  and (_07677_, _07675_, _07635_);
  or (_07678_, _07677_, _07676_);
  nor (_07679_, _07678_, _07650_);
  nor (_07680_, _07648_, _07631_);
  nor (_07681_, _07680_, _07679_);
  and (_07682_, _07681_, _07475_);
  nor (_07683_, _07681_, _07475_);
  nor (_07684_, _07648_, _07634_);
  nor (_07685_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07686_, _07685_, _07347_);
  and (_07687_, _07648_, _07686_);
  or (_07688_, _07687_, _07684_);
  and (_07689_, _07688_, _07461_);
  and (_07690_, \oc8051_golden_model_1.B [0], _03320_);
  not (_07691_, _07690_);
  nor (_07692_, _07688_, _07461_);
  nor (_07693_, _07692_, _07689_);
  and (_07694_, _07693_, _07691_);
  nor (_07695_, _07694_, _07689_);
  nor (_07696_, _07695_, _07683_);
  nor (_07697_, _07696_, _07682_);
  nor (_07698_, _07673_, _07476_);
  nor (_07699_, _07698_, _07674_);
  not (_07700_, _07699_);
  nor (_07701_, _07700_, _07697_);
  nor (_07702_, _07701_, _07674_);
  nor (_07703_, _07702_, _07668_);
  nor (_07704_, _07703_, _07667_);
  nor (_07705_, _07704_, _07659_);
  nor (_07706_, _07705_, _07656_);
  and (_07707_, _06880_, \oc8051_golden_model_1.ACC [7]);
  nor (_07708_, _07707_, _07479_);
  nor (_07709_, _07708_, _07706_);
  not (_07710_, _07479_);
  nor (_07711_, _07649_, _07470_);
  nor (_07712_, _07711_, _07710_);
  nor (_07713_, _07712_, _07709_);
  and (_07714_, _07713_, _07649_);
  nor (_07715_, _07714_, _07470_);
  and (_07716_, _07715_, \oc8051_golden_model_1.B [7]);
  and (_07717_, _07715_, _06880_);
  nor (_07718_, _07717_, _07419_);
  not (_07719_, _07718_);
  not (_07720_, \oc8051_golden_model_1.B [6]);
  and (_07721_, _07704_, _07659_);
  nor (_07722_, _07721_, _07705_);
  nor (_07723_, _07722_, _07713_);
  not (_07724_, _07713_);
  nor (_07725_, _07724_, _07655_);
  nor (_07726_, _07725_, _07723_);
  nor (_07727_, _07726_, _07720_);
  and (_07728_, _07726_, _07720_);
  nor (_07729_, _07668_, _07667_);
  nor (_07730_, _07729_, _07702_);
  and (_07731_, _07729_, _07702_);
  or (_07732_, _07731_, _07730_);
  nor (_07733_, _07732_, _07713_);
  nor (_07734_, _07724_, _07666_);
  nor (_07735_, _07734_, _07733_);
  nor (_07736_, _07735_, _07478_);
  and (_07737_, _07735_, _07478_);
  not (_07738_, _07737_);
  and (_07739_, _07700_, _07697_);
  nor (_07740_, _07739_, _07701_);
  nor (_07741_, _07740_, _07713_);
  nor (_07742_, _07724_, _07673_);
  nor (_07743_, _07742_, _07741_);
  nor (_07744_, _07743_, _07477_);
  and (_07745_, _07713_, _07681_);
  nor (_07746_, _07683_, _07682_);
  and (_07747_, _07746_, _07695_);
  nor (_07748_, _07746_, _07695_);
  nor (_07749_, _07748_, _07747_);
  nor (_07750_, _07749_, _07713_);
  or (_07751_, _07750_, _07745_);
  and (_07752_, _07751_, _07476_);
  nor (_07753_, _07751_, _07476_);
  nor (_07754_, _07753_, _07752_);
  nor (_07755_, _07693_, _07691_);
  nor (_07756_, _07755_, _07694_);
  nor (_07757_, _07756_, _07713_);
  nor (_07758_, _07724_, _07688_);
  nor (_07759_, _07758_, _07757_);
  nor (_07760_, _07759_, _07475_);
  and (_07761_, _07759_, _07475_);
  nor (_07762_, _07761_, _07760_);
  and (_07763_, _07762_, _07754_);
  and (_07764_, _07713_, _03320_);
  and (_07765_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07766_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07767_, _07766_, _07765_);
  nor (_07768_, _07713_, _07767_);
  nor (_07769_, _07768_, _07764_);
  and (_07770_, _07769_, _07461_);
  nor (_07771_, _07769_, _07461_);
  and (_07772_, _07467_, \oc8051_golden_model_1.ACC [0]);
  not (_07773_, _07772_);
  nor (_07774_, _07773_, _07771_);
  nor (_07775_, _07774_, _07770_);
  and (_07776_, _07775_, _07763_);
  and (_07777_, _07760_, _07754_);
  nor (_07778_, _07777_, _07753_);
  not (_07779_, _07778_);
  nor (_07780_, _07779_, _07776_);
  and (_07781_, _07743_, _07477_);
  nor (_07782_, _07781_, _07780_);
  or (_07783_, _07782_, _07744_);
  and (_07784_, _07783_, _07738_);
  nor (_07785_, _07784_, _07736_);
  nor (_07786_, _07785_, _07728_);
  or (_07787_, _07786_, _07727_);
  and (_07788_, _07787_, _07719_);
  nor (_07789_, _07788_, _07716_);
  nor (_07790_, _07737_, _07736_);
  nor (_07791_, _07781_, _07744_);
  and (_07792_, _07791_, _07790_);
  nor (_07793_, _07728_, _07727_);
  and (_07794_, _07793_, _07719_);
  and (_07795_, _07794_, _07792_);
  nor (_07796_, _07771_, _07770_);
  and (_07797_, \oc8051_golden_model_1.B [0], _03397_);
  not (_07798_, _07797_);
  and (_07799_, _07798_, _07796_);
  and (_07800_, _07799_, _07773_);
  and (_07801_, _07800_, _07763_);
  and (_07802_, _07801_, _07795_);
  nor (_07803_, _07802_, _07789_);
  and (_07804_, _07803_, _07714_);
  not (_07805_, _07455_);
  or (_07806_, _07470_, _07805_);
  or (_07807_, _07806_, _07804_);
  and (_07808_, _07807_, _03651_);
  and (_07809_, _07808_, _07460_);
  and (_07810_, _05961_, _05379_);
  or (_07811_, _07810_, _06882_);
  and (_07812_, _07811_, _03649_);
  and (_07813_, _06247_, _05379_);
  or (_07814_, _07813_, _06882_);
  and (_07815_, _07814_, _03650_);
  or (_07816_, _07815_, _03778_);
  or (_07817_, _07816_, _07812_);
  or (_07818_, _07817_, _07809_);
  and (_07819_, _06458_, _05379_);
  or (_07820_, _07819_, _06882_);
  or (_07821_, _07820_, _04589_);
  and (_07822_, _07821_, _04596_);
  and (_07823_, _07822_, _07818_);
  or (_07824_, _06882_, _05397_);
  and (_07825_, _07814_, _03655_);
  and (_07826_, _07825_, _07824_);
  or (_07827_, _07826_, _07823_);
  and (_07828_, _07827_, _04594_);
  and (_07829_, _06899_, _03773_);
  and (_07830_, _07829_, _07824_);
  or (_07831_, _07830_, _03653_);
  or (_07832_, _07831_, _07828_);
  nor (_07833_, _05959_, _06883_);
  or (_07834_, _06882_, _04608_);
  or (_07835_, _07834_, _07833_);
  and (_07836_, _07835_, _04606_);
  and (_07837_, _07836_, _07832_);
  nor (_07838_, _06457_, _06883_);
  or (_07839_, _07838_, _06882_);
  and (_07840_, _07839_, _03786_);
  or (_07841_, _07840_, _03809_);
  or (_07842_, _07841_, _07837_);
  or (_07843_, _06896_, _04260_);
  and (_07844_, _07843_, _03206_);
  and (_07845_, _07844_, _07842_);
  and (_07846_, _06893_, _03205_);
  or (_07847_, _07846_, _03816_);
  or (_07848_, _07847_, _07845_);
  and (_07849_, _05895_, _05379_);
  or (_07850_, _06882_, _03820_);
  or (_07851_, _07850_, _07849_);
  and (_07852_, _07851_, _43227_);
  and (_07853_, _07852_, _07848_);
  or (_07854_, _07853_, _06881_);
  and (_40745_, _07854_, _41991_);
  nor (_07855_, _43227_, _06061_);
  not (_07856_, _05442_);
  and (_07857_, _05903_, \oc8051_golden_model_1.PSW [7]);
  and (_07858_, _07857_, _07856_);
  nor (_07859_, _07858_, _05289_);
  and (_07860_, _07858_, _05289_);
  nor (_07861_, _07860_, _07859_);
  and (_07862_, _07861_, \oc8051_golden_model_1.ACC [7]);
  nor (_07863_, _07861_, \oc8051_golden_model_1.ACC [7]);
  nor (_07864_, _07863_, _07862_);
  nor (_07865_, _07857_, _07856_);
  nor (_07866_, _07865_, _07858_);
  and (_07867_, _07866_, \oc8051_golden_model_1.ACC [6]);
  nor (_07868_, _07866_, _07484_);
  and (_07869_, _07866_, _07484_);
  nor (_07870_, _07869_, _07868_);
  not (_07871_, _05552_);
  not (_07872_, _05840_);
  and (_07873_, _05899_, \oc8051_golden_model_1.PSW [7]);
  and (_07874_, _07873_, _05900_);
  and (_07875_, _07874_, _07872_);
  nor (_07876_, _07875_, _07871_);
  nor (_07877_, _07876_, _07857_);
  and (_07878_, _07877_, \oc8051_golden_model_1.ACC [5]);
  nor (_07879_, _07877_, _07530_);
  and (_07880_, _07877_, _07530_);
  nor (_07881_, _07880_, _07879_);
  nor (_07882_, _07874_, _07872_);
  nor (_07883_, _07882_, _07875_);
  and (_07884_, _07883_, \oc8051_golden_model_1.ACC [4]);
  nor (_07885_, _07883_, _07536_);
  and (_07886_, _07883_, _07536_);
  nor (_07887_, _07886_, _07885_);
  not (_07888_, _04944_);
  not (_07889_, _05130_);
  and (_07890_, _05899_, _07889_);
  and (_07891_, _07890_, \oc8051_golden_model_1.PSW [7]);
  nor (_07892_, _07891_, _07888_);
  nor (_07893_, _07892_, _07874_);
  and (_07894_, _07893_, \oc8051_golden_model_1.ACC [3]);
  nor (_07895_, _07893_, _07628_);
  and (_07896_, _07893_, _07628_);
  nor (_07897_, _07896_, _07895_);
  nor (_07898_, _07873_, _07889_);
  nor (_07899_, _07898_, _07891_);
  and (_07900_, _07899_, \oc8051_golden_model_1.ACC [2]);
  nor (_07901_, _07899_, _07634_);
  and (_07902_, _07899_, _07634_);
  nor (_07903_, _07902_, _07901_);
  and (_07904_, _04491_, \oc8051_golden_model_1.PSW [7]);
  nor (_07905_, _07904_, _05898_);
  nor (_07906_, _07905_, _07873_);
  and (_07907_, _07906_, \oc8051_golden_model_1.ACC [1]);
  and (_07908_, _07906_, _03320_);
  nor (_07909_, _07906_, _03320_);
  nor (_07910_, _07909_, _07908_);
  not (_07911_, \oc8051_golden_model_1.PSW [7]);
  and (_07912_, _04510_, _07911_);
  nor (_07913_, _07912_, _07904_);
  and (_07914_, _07913_, \oc8051_golden_model_1.ACC [0]);
  not (_07915_, _07914_);
  nor (_07916_, _07915_, _07910_);
  nor (_07917_, _07916_, _07907_);
  nor (_07918_, _07917_, _07903_);
  nor (_07919_, _07918_, _07900_);
  nor (_07920_, _07919_, _07897_);
  nor (_07921_, _07920_, _07894_);
  nor (_07922_, _07921_, _07887_);
  nor (_07923_, _07922_, _07884_);
  nor (_07924_, _07923_, _07881_);
  nor (_07925_, _07924_, _07878_);
  nor (_07926_, _07925_, _07870_);
  nor (_07927_, _07926_, _07867_);
  nor (_07928_, _07927_, _07864_);
  and (_07929_, _07927_, _07864_);
  nor (_07930_, _07929_, _07928_);
  and (_07931_, _03666_, _03247_);
  nor (_07932_, _05964_, _04220_);
  nor (_07933_, _07932_, _07931_);
  or (_07934_, _07933_, _07930_);
  nor (_07935_, _06171_, \oc8051_golden_model_1.ACC [7]);
  nand (_07936_, _07935_, _04207_);
  nor (_07937_, _05371_, _06061_);
  and (_07938_, _06247_, _05371_);
  nor (_07939_, _07938_, _07937_);
  or (_07940_, _07939_, _06457_);
  nor (_07941_, _07940_, _04596_);
  and (_07942_, _03675_, _03237_);
  or (_07943_, _06456_, _03772_);
  not (_07944_, _04198_);
  not (_07945_, _04200_);
  nor (_07946_, _05289_, _06061_);
  or (_07947_, _07946_, _07945_);
  and (_07948_, _07947_, _07944_);
  and (_07949_, _05961_, _05371_);
  nor (_07950_, _07949_, _07937_);
  nand (_07951_, _07950_, _03649_);
  and (_07952_, _04197_, _03230_);
  not (_07953_, _07952_);
  and (_07954_, _06171_, \oc8051_golden_model_1.ACC [7]);
  nor (_07955_, _07954_, _07935_);
  or (_07956_, _07955_, _07953_);
  not (_07957_, _05371_);
  nor (_07958_, _07957_, _05289_);
  nor (_07959_, _07958_, _07937_);
  nand (_07960_, _07959_, _07441_);
  and (_07961_, _06846_, \oc8051_golden_model_1.PSW [7]);
  nor (_07962_, _07961_, _06834_);
  and (_07963_, _07961_, _06834_);
  nor (_07964_, _07963_, _07962_);
  and (_07965_, _07964_, \oc8051_golden_model_1.ACC [7]);
  nor (_07966_, _07964_, \oc8051_golden_model_1.ACC [7]);
  nor (_07967_, _07966_, _07965_);
  and (_07968_, _06841_, _06843_);
  and (_07969_, _07968_, \oc8051_golden_model_1.PSW [7]);
  and (_07970_, _07969_, _06842_);
  nor (_07971_, _07970_, _06531_);
  nor (_07972_, _07971_, _07961_);
  nor (_07973_, _07972_, _07484_);
  and (_07974_, _07972_, _07484_);
  nor (_07975_, _07969_, _06842_);
  nor (_07976_, _07975_, _07970_);
  and (_07977_, _07976_, _07530_);
  nor (_07978_, _07976_, _07530_);
  and (_07979_, _06837_, \oc8051_golden_model_1.PSW [7]);
  and (_07980_, _07979_, _06840_);
  nor (_07981_, _07980_, _06843_);
  nor (_07982_, _07981_, _07969_);
  nor (_07983_, _07982_, _07536_);
  nor (_07984_, _07983_, _07978_);
  nor (_07985_, _07984_, _07977_);
  nor (_07986_, _07978_, _07977_);
  and (_07987_, _07982_, _07536_);
  nor (_07988_, _07987_, _07983_);
  and (_07989_, _07988_, _07986_);
  not (_07990_, _07989_);
  and (_07991_, _06837_, _06839_);
  and (_07992_, _07991_, \oc8051_golden_model_1.PSW [7]);
  nor (_07993_, _07992_, _06838_);
  nor (_07994_, _07993_, _07980_);
  nor (_07995_, _07994_, _07628_);
  and (_07996_, _07994_, _07628_);
  nor (_07997_, _07996_, _07995_);
  nor (_07998_, _07979_, _06839_);
  nor (_07999_, _07998_, _07992_);
  nor (_08000_, _07999_, _07634_);
  and (_08001_, _07999_, _07634_);
  nor (_08002_, _08001_, _08000_);
  and (_08003_, _08002_, _07997_);
  and (_08004_, _06836_, \oc8051_golden_model_1.PSW [7]);
  nor (_08005_, _08004_, _06835_);
  nor (_08006_, _08005_, _07979_);
  and (_08007_, _08006_, _03320_);
  nor (_08008_, _08006_, _03320_);
  and (_08009_, _06622_, _07911_);
  nor (_08010_, _08009_, _08004_);
  nor (_08011_, _08010_, _03397_);
  nor (_08012_, _08011_, _08008_);
  or (_08013_, _08012_, _08007_);
  and (_08014_, _08013_, _08003_);
  not (_08015_, _08014_);
  and (_08016_, _08001_, _07997_);
  nor (_08017_, _08016_, _07996_);
  and (_08018_, _08017_, _08015_);
  nor (_08019_, _08008_, _08007_);
  and (_08020_, _08010_, _03397_);
  nor (_08021_, _08011_, _08020_);
  and (_08022_, _08021_, _08019_);
  and (_08023_, _08022_, _08003_);
  nor (_08024_, _08023_, _08018_);
  nor (_08025_, _08024_, _07990_);
  nor (_08026_, _08025_, _07985_);
  nor (_08027_, _08026_, _07974_);
  or (_08028_, _08027_, _07973_);
  or (_08029_, _08028_, _07967_);
  nand (_08030_, _08028_, _07967_);
  and (_08031_, _08030_, _08029_);
  and (_08032_, _04197_, _03276_);
  and (_08033_, _08032_, _08031_);
  and (_08034_, _04563_, _03276_);
  nor (_08035_, _04839_, _03277_);
  or (_08036_, _08035_, _04120_);
  nor (_08037_, _08036_, _08034_);
  not (_08038_, _08037_);
  not (_08039_, _04848_);
  and (_08040_, _04819_, _03997_);
  and (_08041_, _08040_, _08039_);
  not (_08042_, _08041_);
  nand (_08043_, _08042_, _05289_);
  nor (_08044_, _03680_, _03666_);
  nor (_08045_, _08044_, _03261_);
  nor (_08046_, _08045_, _04067_);
  or (_08047_, _04839_, _03261_);
  and (_08048_, _08047_, _08046_);
  not (_08049_, _08048_);
  nand (_08050_, _08049_, _05289_);
  and (_08051_, _03675_, _03945_);
  not (_08052_, _08051_);
  nor (_08053_, _04063_, _06061_);
  and (_08054_, _04063_, _06061_);
  nor (_08055_, _08054_, _08053_);
  nand (_08056_, _08055_, _08048_);
  and (_08057_, _08056_, _08052_);
  and (_08058_, _08057_, _08050_);
  and (_08059_, _08051_, _06171_);
  or (_08060_, _08059_, _08058_);
  and (_08061_, _04515_, _03262_);
  and (_08062_, _08061_, _08060_);
  and (_08063_, _03675_, _03514_);
  and (_08064_, _06185_, _05371_);
  nor (_08065_, _08064_, _07937_);
  nor (_08066_, _08065_, _04515_);
  or (_08067_, _08066_, _08063_);
  or (_08068_, _08067_, _08062_);
  nor (_08069_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_08070_, _08069_, _07628_);
  and (_08071_, _08070_, _07501_);
  and (_08072_, _08071_, \oc8051_golden_model_1.ACC [6]);
  and (_08073_, _08072_, \oc8051_golden_model_1.ACC [7]);
  nor (_08074_, _08072_, \oc8051_golden_model_1.ACC [7]);
  nor (_08075_, _08074_, _08073_);
  and (_08076_, _08070_, \oc8051_golden_model_1.ACC [4]);
  nor (_08077_, _08076_, \oc8051_golden_model_1.ACC [5]);
  nor (_08078_, _08077_, _08071_);
  nor (_08079_, _08071_, \oc8051_golden_model_1.ACC [6]);
  nor (_08080_, _08079_, _08072_);
  nor (_08081_, _08080_, _08078_);
  not (_08082_, _08081_);
  and (_08083_, _08082_, _08075_);
  nor (_08084_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_08085_, _08084_, _08081_);
  nor (_08086_, _08085_, _08075_);
  nor (_08087_, _08086_, _08083_);
  not (_08088_, _08087_);
  nand (_08089_, _08088_, _08063_);
  and (_08090_, _08089_, _03604_);
  and (_08091_, _08090_, _08068_);
  nor (_08092_, _05983_, _06061_);
  and (_08093_, _06042_, _05983_);
  nor (_08094_, _08093_, _08092_);
  nor (_08095_, _08094_, _03516_);
  nor (_08096_, _07959_, _04524_);
  or (_08097_, _08096_, _08042_);
  or (_08098_, _08097_, _08095_);
  or (_08099_, _08098_, _08091_);
  and (_08100_, _08099_, _08043_);
  or (_08101_, _08100_, _04529_);
  not (_08102_, _04529_);
  or (_08103_, _06171_, _08102_);
  and (_08104_, _08103_, _03611_);
  and (_08105_, _08104_, _08101_);
  and (_08106_, _03675_, _03509_);
  nor (_08107_, _06211_, _03611_);
  or (_08108_, _08107_, _08106_);
  or (_08109_, _08108_, _08105_);
  nand (_08110_, _08106_, _07628_);
  and (_08111_, _08110_, _08109_);
  or (_08112_, _08111_, _03511_);
  and (_08113_, _06038_, _05983_);
  nor (_08114_, _08113_, _08092_);
  nand (_08115_, _08114_, _03511_);
  and (_08116_, _08115_, _03505_);
  and (_08117_, _08116_, _08112_);
  and (_08118_, _08093_, _06216_);
  nor (_08119_, _08118_, _08092_);
  nor (_08120_, _08119_, _03505_);
  or (_08121_, _08120_, _06919_);
  or (_08122_, _08121_, _08117_);
  nor (_08123_, _07397_, _07395_);
  nor (_08124_, _08123_, _07398_);
  or (_08125_, _08124_, _06925_);
  and (_08126_, _08125_, _08122_);
  or (_08127_, _08126_, _08038_);
  not (_08128_, _08032_);
  not (_08129_, _07864_);
  nor (_08130_, _07885_, _07879_);
  nor (_08131_, _08130_, _07880_);
  and (_08132_, _07887_, _07881_);
  not (_08133_, _08132_);
  and (_08134_, _07903_, _07897_);
  nor (_08135_, _07913_, _03397_);
  nor (_08136_, _08135_, _07909_);
  or (_08137_, _08136_, _07908_);
  and (_08138_, _08137_, _08134_);
  not (_08139_, _08138_);
  and (_08140_, _07902_, _07897_);
  nor (_08141_, _08140_, _07896_);
  and (_08142_, _08141_, _08139_);
  and (_08143_, _07913_, _03397_);
  nor (_08144_, _08135_, _08143_);
  and (_08145_, _08144_, _07910_);
  and (_08146_, _08145_, _08134_);
  nor (_08147_, _08146_, _08142_);
  nor (_08148_, _08147_, _08133_);
  nor (_08149_, _08148_, _08131_);
  nor (_08150_, _08149_, _07869_);
  or (_08151_, _08150_, _07868_);
  and (_08152_, _08151_, _08129_);
  nor (_08153_, _08151_, _08129_);
  or (_08154_, _08153_, _08152_);
  or (_08155_, _08154_, _08037_);
  and (_08156_, _08155_, _08128_);
  and (_08157_, _08156_, _08127_);
  or (_08158_, _08157_, _03635_);
  or (_08159_, _08158_, _08033_);
  and (_08160_, _03675_, _03276_);
  not (_08161_, _08160_);
  and (_08162_, _05363_, \oc8051_golden_model_1.P0INREG [6]);
  and (_08163_, _05383_, \oc8051_golden_model_1.P1INREG [6]);
  not (_08164_, _08163_);
  and (_08165_, _05386_, \oc8051_golden_model_1.P2INREG [6]);
  and (_08166_, _05388_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_08167_, _08166_, _08165_);
  and (_08168_, _08167_, _08164_);
  nand (_08169_, _08168_, _05477_);
  nor (_08170_, _08169_, _08162_);
  and (_08171_, _08170_, _05470_);
  and (_08172_, _08171_, _05460_);
  and (_08173_, _08172_, _05443_);
  not (_08174_, _08173_);
  not (_08175_, _05612_);
  and (_08176_, _08175_, _05642_);
  nor (_08177_, _05615_, _05613_);
  and (_08178_, _08177_, _05624_);
  and (_08179_, _05386_, \oc8051_golden_model_1.P2INREG [3]);
  and (_08180_, _05388_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_08181_, _08180_, _08179_);
  and (_08182_, _05363_, \oc8051_golden_model_1.P0INREG [3]);
  and (_08183_, _05383_, \oc8051_golden_model_1.P1INREG [3]);
  nor (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _08181_);
  and (_08186_, _08185_, _08178_);
  and (_08187_, _08186_, _08176_);
  and (_08188_, _05621_, _05632_);
  and (_08189_, _08188_, _05611_);
  and (_08190_, _08189_, _08187_);
  and (_08191_, _08190_, _05602_);
  not (_08192_, _08191_);
  and (_08193_, _05383_, \oc8051_golden_model_1.P1INREG [2]);
  not (_08194_, _08193_);
  not (_08195_, _05766_);
  and (_08196_, _05386_, \oc8051_golden_model_1.P2INREG [2]);
  and (_08197_, _05388_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_08198_, _08197_, _08196_);
  and (_08199_, _08198_, _08195_);
  and (_08200_, _08199_, _08194_);
  and (_08201_, _05784_, _05781_);
  and (_08202_, _05363_, \oc8051_golden_model_1.P0INREG [2]);
  not (_08203_, _08202_);
  and (_08204_, _08203_, _05787_);
  and (_08205_, _08204_, _08201_);
  and (_08206_, _08205_, _08200_);
  and (_08207_, _08206_, _05764_);
  and (_08208_, _08207_, _05746_);
  not (_08209_, _08208_);
  and (_08210_, _05383_, \oc8051_golden_model_1.P1INREG [1]);
  not (_08211_, _08210_);
  and (_08212_, _05386_, \oc8051_golden_model_1.P2INREG [1]);
  and (_08213_, _05388_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_08214_, _08213_, _08212_);
  and (_08215_, _08214_, _05659_);
  and (_08216_, _08215_, _08211_);
  and (_08217_, _05363_, \oc8051_golden_model_1.P0INREG [1]);
  not (_08218_, _08217_);
  and (_08219_, _08218_, _05675_);
  and (_08220_, _08219_, _08216_);
  and (_08221_, _08220_, _05657_);
  and (_08222_, _08221_, _05696_);
  and (_08223_, _08222_, _05651_);
  not (_08224_, _08223_);
  and (_08225_, _05383_, \oc8051_golden_model_1.P1INREG [0]);
  not (_08226_, _08225_);
  not (_08227_, _05721_);
  and (_08228_, _05386_, \oc8051_golden_model_1.P2INREG [0]);
  and (_08229_, _05388_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_08230_, _08229_, _08228_);
  and (_08231_, _08230_, _08227_);
  and (_08232_, _08231_, _08226_);
  and (_08233_, _05363_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_08234_, _08233_, _05739_);
  and (_08235_, _08234_, _05737_);
  and (_08236_, _08235_, _08232_);
  and (_08237_, _08236_, _05718_);
  and (_08238_, _08237_, _05700_);
  nor (_08239_, _08238_, _07911_);
  and (_08240_, _08239_, _08224_);
  and (_08241_, _08240_, _08209_);
  and (_08242_, _08241_, _08192_);
  and (_08243_, _05363_, \oc8051_golden_model_1.P0INREG [5]);
  not (_08244_, _08243_);
  and (_08245_, _05383_, \oc8051_golden_model_1.P1INREG [5]);
  not (_08246_, _08245_);
  and (_08247_, _05386_, \oc8051_golden_model_1.P2INREG [5]);
  and (_08248_, _05388_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_08249_, _08248_, _08247_);
  and (_08250_, _08249_, _08246_);
  and (_08251_, _08250_, _05587_);
  and (_08252_, _08251_, _08244_);
  and (_08253_, _08252_, _05580_);
  and (_08254_, _08253_, _05570_);
  and (_08255_, _08254_, _05553_);
  and (_08256_, _05383_, \oc8051_golden_model_1.P1INREG [4]);
  not (_08257_, _08256_);
  and (_08258_, _05386_, \oc8051_golden_model_1.P2INREG [4]);
  and (_08259_, _05388_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_08260_, _08259_, _08258_);
  and (_08261_, _08260_, _05849_);
  and (_08262_, _08261_, _08257_);
  and (_08263_, _05363_, \oc8051_golden_model_1.P0INREG [4]);
  not (_08264_, _08263_);
  and (_08265_, _08264_, _05865_);
  and (_08266_, _08265_, _08262_);
  and (_08267_, _08266_, _05847_);
  and (_08268_, _08267_, _05886_);
  and (_08269_, _08268_, _05841_);
  nor (_08270_, _08269_, _08255_);
  and (_08271_, _08270_, _08242_);
  and (_08272_, _08271_, _08174_);
  nor (_08273_, _08272_, _06211_);
  and (_08274_, _08272_, _06211_);
  nor (_08275_, _08274_, _08273_);
  and (_08276_, _08275_, \oc8051_golden_model_1.ACC [7]);
  nor (_08277_, _08275_, \oc8051_golden_model_1.ACC [7]);
  nor (_08278_, _08277_, _08276_);
  nor (_08279_, _08271_, _08174_);
  nor (_08280_, _08279_, _08272_);
  nor (_08281_, _08280_, _07484_);
  and (_08282_, _08280_, _07484_);
  not (_08283_, _08255_);
  not (_08284_, _08269_);
  and (_08285_, _08242_, _08284_);
  nor (_08286_, _08285_, _08283_);
  nor (_08287_, _08286_, _08271_);
  nor (_08288_, _08287_, _07530_);
  and (_08289_, _08287_, _07530_);
  nor (_08290_, _08289_, _08288_);
  nor (_08291_, _08242_, _08284_);
  nor (_08292_, _08291_, _08285_);
  nor (_08293_, _08292_, _07536_);
  and (_08294_, _08292_, _07536_);
  nor (_08295_, _08294_, _08293_);
  and (_08296_, _08295_, _08290_);
  nor (_08297_, _08241_, _08192_);
  nor (_08298_, _08297_, _08242_);
  nor (_08299_, _08298_, _07628_);
  and (_08300_, _08298_, _07628_);
  nor (_08301_, _08300_, _08299_);
  nor (_08302_, _08240_, _08209_);
  nor (_08303_, _08302_, _08241_);
  nor (_08304_, _08303_, _07634_);
  and (_08305_, _08303_, _07634_);
  nor (_08306_, _08305_, _08304_);
  and (_08307_, _08306_, _08301_);
  nor (_08308_, _08239_, _08224_);
  nor (_08309_, _08308_, _08240_);
  nor (_08310_, _08309_, _03320_);
  and (_08311_, _08309_, _03320_);
  and (_08312_, _08238_, _07911_);
  nor (_08313_, _08312_, _08239_);
  and (_08314_, _08313_, _03397_);
  nor (_08315_, _08314_, _08311_);
  or (_08316_, _08315_, _08310_);
  and (_08317_, _08316_, _08307_);
  and (_08318_, _08304_, _08301_);
  or (_08319_, _08318_, _08299_);
  nor (_08320_, _08319_, _08317_);
  not (_08321_, _08320_);
  and (_08322_, _08321_, _08296_);
  nor (_08323_, _08293_, _08288_);
  or (_08324_, _08323_, _08289_);
  not (_08325_, _08324_);
  nor (_08326_, _08325_, _08322_);
  nor (_08327_, _08326_, _08282_);
  nor (_08328_, _08327_, _08281_);
  nor (_08329_, _08328_, _08278_);
  and (_08330_, _08328_, _08278_);
  or (_08331_, _08330_, _08329_);
  or (_08332_, _08331_, _03640_);
  and (_08333_, _08332_, _08161_);
  and (_08334_, _08333_, _08159_);
  and (_08335_, _05295_, \oc8051_golden_model_1.PSW [7]);
  and (_08336_, _08335_, _05302_);
  and (_08337_, _08336_, _05374_);
  and (_08338_, _08337_, _05056_);
  nor (_08339_, _08338_, _04559_);
  and (_08340_, _08337_, _03557_);
  nor (_08341_, _08340_, _08339_);
  and (_08342_, _08341_, \oc8051_golden_model_1.ACC [7]);
  nor (_08343_, _08341_, \oc8051_golden_model_1.ACC [7]);
  nor (_08344_, _08343_, _08342_);
  not (_08345_, _08344_);
  nor (_08346_, _08337_, _05056_);
  nor (_08347_, _08346_, _08338_);
  nor (_08348_, _08347_, _07484_);
  and (_08349_, _08347_, _07484_);
  and (_08350_, _08336_, _05327_);
  nor (_08351_, _08350_, _05334_);
  nor (_08352_, _08351_, _08337_);
  nor (_08353_, _08352_, _07530_);
  and (_08354_, _08352_, _07530_);
  nor (_08355_, _08354_, _08353_);
  nor (_08356_, _08336_, _05327_);
  nor (_08357_, _08356_, _08350_);
  nor (_08358_, _08357_, _07536_);
  and (_08359_, _08357_, _07536_);
  nor (_08360_, _08359_, _08358_);
  and (_08361_, _08360_, _08355_);
  not (_08362_, _08361_);
  nor (_08363_, _06025_, _03558_);
  nor (_08364_, _08363_, _08336_);
  and (_08365_, _08364_, _07628_);
  nor (_08366_, _08364_, _07628_);
  nor (_08367_, _08366_, _08365_);
  nor (_08368_, _08335_, _03899_);
  nor (_08369_, _08368_, _06025_);
  nor (_08370_, _08369_, _07634_);
  and (_08371_, _08369_, _07634_);
  nor (_08372_, _08371_, _08370_);
  and (_08373_, _08372_, _08367_);
  not (_08374_, _08373_);
  nor (_08375_, _04042_, _07911_);
  and (_08376_, _04042_, _07911_);
  nor (_08377_, _08376_, _08375_);
  and (_08378_, _08377_, _03397_);
  nor (_08379_, _08377_, _03397_);
  nor (_08380_, _08379_, _08378_);
  nor (_08381_, _04434_, _03320_);
  and (_08382_, _04434_, _03320_);
  nor (_08383_, _08382_, _08381_);
  and (_08384_, \oc8051_golden_model_1.PSW [7], _03397_);
  and (_08385_, _07911_, \oc8051_golden_model_1.ACC [0]);
  nor (_08386_, _08385_, _04042_);
  nor (_08387_, _08386_, _08384_);
  and (_08388_, _08387_, _08383_);
  nor (_08389_, _08387_, _08383_);
  nor (_08390_, _08389_, _08388_);
  nand (_08391_, _08390_, _08380_);
  nor (_08392_, _08391_, _08374_);
  nor (_08393_, _08375_, _04435_);
  nor (_08394_, _08393_, _08335_);
  and (_08395_, _08394_, _03320_);
  nor (_08396_, _08394_, _03320_);
  nor (_08397_, _08379_, _08396_);
  nor (_08398_, _08397_, _08395_);
  nor (_08399_, _08398_, _08374_);
  and (_08400_, _08371_, _08367_);
  nor (_08401_, _08400_, _08365_);
  not (_08402_, _08401_);
  nor (_08403_, _08402_, _08399_);
  nor (_08404_, _08403_, _08392_);
  nor (_08405_, _08404_, _08362_);
  not (_08406_, _08405_);
  nor (_08407_, _08358_, _08353_);
  or (_08408_, _08407_, _08354_);
  and (_08409_, _08408_, _08406_);
  nor (_08410_, _08409_, _08349_);
  or (_08411_, _08410_, _08348_);
  and (_08412_, _08411_, _08345_);
  nor (_08413_, _08411_, _08345_);
  or (_08414_, _08413_, _08412_);
  and (_08415_, _08414_, _08160_);
  or (_08416_, _08415_, _03371_);
  or (_08417_, _08416_, _08334_);
  or (_08418_, _03463_, _03285_);
  and (_08419_, _08418_, _03501_);
  and (_08420_, _08419_, _08417_);
  not (_08421_, _05983_);
  nor (_08422_, _06026_, _08421_);
  nor (_08423_, _08422_, _08092_);
  nor (_08424_, _08423_, _03501_);
  or (_08425_, _08424_, _07441_);
  or (_08426_, _08425_, _08420_);
  and (_08427_, _08426_, _07960_);
  or (_08428_, _08427_, _05969_);
  and (_08429_, _06171_, _05371_);
  nor (_08430_, _08429_, _07937_);
  nand (_08431_, _08430_, _05969_);
  and (_08432_, _08431_, _03275_);
  and (_08433_, _08432_, _08428_);
  nor (_08434_, _06443_, _07957_);
  nor (_08435_, _08434_, _07937_);
  nor (_08436_, _08435_, _03275_);
  or (_08437_, _08436_, _07455_);
  or (_08438_, _08437_, _08433_);
  or (_08439_, _07473_, _07805_);
  and (_08440_, _08439_, _08438_);
  or (_08441_, _08440_, _03313_);
  or (_08442_, _03463_, _03314_);
  and (_08443_, _08442_, _08441_);
  or (_08444_, _08443_, _03650_);
  and (_08445_, _03675_, _03226_);
  not (_08446_, _08445_);
  nand (_08447_, _07939_, _03650_);
  and (_08448_, _08447_, _08446_);
  and (_08449_, _08448_, _08444_);
  nand (_08450_, _08445_, _03463_);
  or (_08451_, _03983_, _03961_);
  not (_08452_, _08451_);
  not (_08453_, _03230_);
  nor (_08454_, _03587_, _03584_);
  or (_08455_, _08454_, _08453_);
  and (_08456_, _08455_, _08452_);
  nand (_08457_, _08456_, _08450_);
  or (_08458_, _08457_, _08449_);
  and (_08459_, _05289_, _06061_);
  nor (_08460_, _08459_, _07946_);
  or (_08461_, _08456_, _08460_);
  and (_08462_, _03589_, _03230_);
  nor (_08463_, _08462_, _04188_);
  and (_08464_, _08463_, _08461_);
  and (_08465_, _08464_, _08458_);
  not (_08466_, _08460_);
  nor (_08467_, _08463_, _08466_);
  or (_08468_, _08467_, _07952_);
  or (_08469_, _08468_, _08465_);
  and (_08470_, _08469_, _07956_);
  or (_08471_, _08470_, _03776_);
  and (_08472_, _03675_, _03230_);
  not (_08473_, _08472_);
  or (_08474_, _06458_, _03777_);
  and (_08475_, _08474_, _08473_);
  and (_08476_, _08475_, _08471_);
  and (_08477_, _03463_, \oc8051_golden_model_1.ACC [7]);
  nor (_08478_, _03463_, \oc8051_golden_model_1.ACC [7]);
  nor (_08479_, _08478_, _08477_);
  and (_08480_, _08472_, _08479_);
  or (_08481_, _08480_, _03649_);
  or (_08482_, _08481_, _08476_);
  and (_08483_, _08482_, _07951_);
  or (_08484_, _08483_, _03778_);
  or (_08485_, _07937_, _04589_);
  and (_08486_, _03574_, _03237_);
  nor (_08487_, _08486_, _04357_);
  and (_08488_, _08487_, _08485_);
  and (_08489_, _08488_, _08484_);
  not (_08490_, _08487_);
  and (_08491_, _08490_, _07946_);
  or (_08492_, _08491_, _04200_);
  or (_08493_, _08492_, _08489_);
  and (_08494_, _08493_, _07948_);
  and (_08495_, _07954_, _04198_);
  or (_08496_, _08495_, _03771_);
  or (_08497_, _08496_, _08494_);
  and (_08498_, _08497_, _07943_);
  or (_08499_, _08498_, _07942_);
  not (_08500_, _07942_);
  or (_08501_, _08477_, _08500_);
  and (_08502_, _08501_, _04596_);
  and (_08503_, _08502_, _08499_);
  or (_08504_, _08503_, _07941_);
  and (_08505_, _03584_, _03235_);
  nor (_08506_, _08505_, _03954_);
  and (_08507_, _08506_, _08504_);
  nor (_08508_, _05080_, _04204_);
  nor (_08509_, _08506_, _08459_);
  or (_08510_, _08509_, _08508_);
  or (_08511_, _08510_, _08507_);
  and (_08512_, _03568_, _03235_);
  nor (_08513_, _04206_, _08512_);
  and (_08514_, _03570_, _03235_);
  nor (_08515_, _08459_, _08514_);
  or (_08516_, _08515_, _08513_);
  and (_08517_, _08516_, _08511_);
  not (_08518_, _08514_);
  nor (_08519_, _08459_, _08518_);
  or (_08520_, _08519_, _04207_);
  or (_08521_, _08520_, _08517_);
  and (_08522_, _08521_, _07936_);
  or (_08523_, _08522_, _03784_);
  and (_08524_, _03675_, _03235_);
  not (_08525_, _08524_);
  nand (_08526_, _06457_, _03784_);
  and (_08527_, _08526_, _08525_);
  and (_08528_, _08527_, _08523_);
  nor (_08529_, _08525_, _08478_);
  or (_08530_, _08529_, _08528_);
  and (_08531_, _08530_, _04608_);
  not (_08532_, _07933_);
  nor (_08533_, _05959_, _07957_);
  nor (_08534_, _08533_, _07937_);
  nor (_08535_, _08534_, _04608_);
  or (_08536_, _08535_, _08532_);
  or (_08537_, _08536_, _08531_);
  and (_08538_, _08537_, _07934_);
  and (_08539_, _04197_, _03247_);
  or (_08540_, _08539_, _08538_);
  not (_08541_, _08539_);
  and (_08542_, _07972_, \oc8051_golden_model_1.ACC [6]);
  nor (_08543_, _07973_, _07974_);
  and (_08544_, _07976_, \oc8051_golden_model_1.ACC [5]);
  and (_08545_, _07982_, \oc8051_golden_model_1.ACC [4]);
  and (_08546_, _07994_, \oc8051_golden_model_1.ACC [3]);
  and (_08547_, _07999_, \oc8051_golden_model_1.ACC [2]);
  and (_08548_, _08006_, \oc8051_golden_model_1.ACC [1]);
  and (_08549_, _08010_, \oc8051_golden_model_1.ACC [0]);
  not (_08550_, _08549_);
  nor (_08551_, _08550_, _08019_);
  nor (_08552_, _08551_, _08548_);
  nor (_08553_, _08552_, _08002_);
  nor (_08554_, _08553_, _08547_);
  nor (_08555_, _08554_, _07997_);
  nor (_08556_, _08555_, _08546_);
  nor (_08557_, _08556_, _07988_);
  nor (_08558_, _08557_, _08545_);
  nor (_08559_, _08558_, _07986_);
  nor (_08560_, _08559_, _08544_);
  nor (_08561_, _08560_, _08543_);
  nor (_08562_, _08561_, _08542_);
  nor (_08563_, _08562_, _07967_);
  and (_08564_, _08562_, _07967_);
  nor (_08565_, _08564_, _08563_);
  or (_08566_, _08565_, _08541_);
  and (_08567_, _08566_, _03783_);
  and (_08568_, _08567_, _08540_);
  and (_08569_, _03675_, _03247_);
  nor (_08570_, _08569_, _03782_);
  not (_08571_, _08570_);
  and (_08572_, _08280_, \oc8051_golden_model_1.ACC [6]);
  nor (_08573_, _08281_, _08282_);
  and (_08574_, _08287_, \oc8051_golden_model_1.ACC [5]);
  and (_08575_, _08292_, \oc8051_golden_model_1.ACC [4]);
  and (_08576_, _08298_, \oc8051_golden_model_1.ACC [3]);
  and (_08577_, _08303_, \oc8051_golden_model_1.ACC [2]);
  and (_08578_, _08309_, \oc8051_golden_model_1.ACC [1]);
  nor (_08579_, _08310_, _08311_);
  and (_08580_, _08313_, \oc8051_golden_model_1.ACC [0]);
  not (_08581_, _08580_);
  nor (_08582_, _08581_, _08579_);
  nor (_08583_, _08582_, _08578_);
  nor (_08584_, _08583_, _08306_);
  nor (_08585_, _08584_, _08577_);
  nor (_08586_, _08585_, _08301_);
  nor (_08587_, _08586_, _08576_);
  nor (_08588_, _08587_, _08295_);
  nor (_08589_, _08588_, _08575_);
  nor (_08590_, _08589_, _08290_);
  nor (_08591_, _08590_, _08574_);
  nor (_08592_, _08591_, _08573_);
  nor (_08593_, _08592_, _08572_);
  nor (_08594_, _08593_, _08278_);
  and (_08595_, _08593_, _08278_);
  nor (_08596_, _08595_, _08594_);
  or (_08597_, _08596_, _08569_);
  and (_08598_, _08597_, _08571_);
  or (_08599_, _08598_, _08568_);
  and (_08600_, _03648_, _03247_);
  not (_08601_, _08600_);
  not (_08602_, _08569_);
  and (_08603_, _08347_, \oc8051_golden_model_1.ACC [6]);
  nor (_08604_, _08348_, _08349_);
  and (_08605_, _08352_, \oc8051_golden_model_1.ACC [5]);
  and (_08606_, _08357_, \oc8051_golden_model_1.ACC [4]);
  and (_08607_, _08364_, \oc8051_golden_model_1.ACC [3]);
  and (_08608_, _08369_, \oc8051_golden_model_1.ACC [2]);
  and (_08609_, _08394_, \oc8051_golden_model_1.ACC [1]);
  nor (_08610_, _08396_, _08395_);
  and (_08611_, _08377_, \oc8051_golden_model_1.ACC [0]);
  not (_08612_, _08611_);
  nor (_08613_, _08612_, _08610_);
  nor (_08614_, _08613_, _08609_);
  nor (_08615_, _08614_, _08372_);
  nor (_08616_, _08615_, _08608_);
  nor (_08617_, _08616_, _08367_);
  nor (_08618_, _08617_, _08607_);
  nor (_08619_, _08618_, _08360_);
  nor (_08620_, _08619_, _08606_);
  nor (_08621_, _08620_, _08355_);
  nor (_08622_, _08621_, _08605_);
  nor (_08623_, _08622_, _08604_);
  nor (_08624_, _08623_, _08603_);
  nor (_08625_, _08624_, _08344_);
  and (_08626_, _08624_, _08344_);
  nor (_08627_, _08626_, _08625_);
  or (_08628_, _08627_, _08602_);
  and (_08629_, _08628_, _08601_);
  and (_08630_, _08629_, _08599_);
  and (_08631_, _08600_, \oc8051_golden_model_1.ACC [6]);
  and (_08632_, _04563_, _03245_);
  not (_08633_, _03245_);
  nor (_08634_, _04839_, _08633_);
  or (_08635_, _08634_, _08632_);
  or (_08636_, _08635_, _08631_);
  or (_08637_, _08636_, _08630_);
  and (_08638_, _03666_, _03245_);
  not (_08639_, _08638_);
  not (_08640_, _08635_);
  nor (_08641_, _05442_, _07484_);
  and (_08642_, _05442_, _07484_);
  nor (_08643_, _08642_, _08641_);
  nor (_08644_, _05552_, _07530_);
  and (_08645_, _05552_, _07530_);
  nor (_08646_, _05840_, _07536_);
  and (_08647_, _05840_, _07536_);
  nor (_08648_, _08647_, _08646_);
  and (_08649_, _04944_, _07628_);
  not (_08650_, _08649_);
  nor (_08651_, _04944_, _07628_);
  not (_08652_, _08651_);
  nor (_08653_, _05130_, _07634_);
  and (_08654_, _05130_, _07634_);
  nor (_08655_, _08654_, _08653_);
  not (_08656_, _08655_);
  and (_08657_, _05898_, \oc8051_golden_model_1.ACC [1]);
  and (_08658_, _04699_, _03320_);
  nor (_08659_, _08658_, _08657_);
  and (_08660_, _04491_, \oc8051_golden_model_1.ACC [0]);
  and (_08661_, _08660_, _08659_);
  nor (_08662_, _08661_, _08657_);
  nor (_08663_, _08662_, _08656_);
  nor (_08664_, _08663_, _08653_);
  nand (_08665_, _08664_, _08652_);
  and (_08666_, _08665_, _08650_);
  and (_08667_, _08666_, _08648_);
  nor (_08668_, _08667_, _08646_);
  nor (_08669_, _08668_, _08645_);
  or (_08670_, _08669_, _08644_);
  and (_08671_, _08670_, _08643_);
  nor (_08672_, _08671_, _08641_);
  nor (_08673_, _08672_, _08460_);
  and (_08674_, _08672_, _08460_);
  or (_08675_, _08674_, _08673_);
  or (_08676_, _08675_, _08640_);
  and (_08677_, _08676_, _08639_);
  and (_08678_, _08677_, _08637_);
  and (_08679_, _04197_, _03245_);
  and (_08680_, _08675_, _08638_);
  or (_08681_, _08680_, _08679_);
  or (_08682_, _08681_, _08678_);
  and (_08683_, _06531_, \oc8051_golden_model_1.ACC [6]);
  nor (_08684_, _06531_, \oc8051_golden_model_1.ACC [6]);
  nor (_08685_, _08683_, _08684_);
  and (_08686_, _06842_, \oc8051_golden_model_1.ACC [5]);
  and (_08687_, _06761_, _07530_);
  or (_08688_, _08687_, _08686_);
  and (_08689_, _06843_, \oc8051_golden_model_1.ACC [4]);
  and (_08690_, _06806_, _07536_);
  nor (_08691_, _08689_, _08690_);
  and (_08692_, _06838_, \oc8051_golden_model_1.ACC [3]);
  and (_08693_, _06668_, _07628_);
  and (_08694_, _06839_, \oc8051_golden_model_1.ACC [2]);
  and (_08695_, _06714_, _07634_);
  nor (_08696_, _08694_, _08695_);
  not (_08697_, _08696_);
  and (_08698_, _06835_, \oc8051_golden_model_1.ACC [1]);
  and (_08699_, _06577_, _03320_);
  nor (_08700_, _08698_, _08699_);
  and (_08701_, _06836_, \oc8051_golden_model_1.ACC [0]);
  and (_08702_, _08701_, _08700_);
  nor (_08703_, _08702_, _08698_);
  nor (_08704_, _08703_, _08697_);
  nor (_08705_, _08704_, _08694_);
  nor (_08706_, _08705_, _08693_);
  or (_08707_, _08706_, _08692_);
  and (_08708_, _08707_, _08691_);
  nor (_08709_, _08708_, _08689_);
  nor (_08710_, _08709_, _08688_);
  or (_08711_, _08710_, _08686_);
  and (_08712_, _08711_, _08685_);
  nor (_08713_, _08712_, _08683_);
  nor (_08714_, _08713_, _07955_);
  and (_08715_, _08713_, _07955_);
  nor (_08716_, _08715_, _08714_);
  nand (_08717_, _08716_, _08679_);
  and (_08718_, _08717_, _03525_);
  and (_08719_, _08718_, _08682_);
  and (_08720_, _03675_, _03245_);
  nor (_08721_, _08720_, _03524_);
  not (_08722_, _08721_);
  and (_08723_, _06211_, _06061_);
  nor (_08724_, _06211_, _06061_);
  nor (_08725_, _08724_, _08723_);
  nor (_08726_, _08173_, _07484_);
  and (_08727_, _08173_, \oc8051_golden_model_1.ACC [6]);
  nor (_08728_, _08173_, \oc8051_golden_model_1.ACC [6]);
  nor (_08729_, _08728_, _08727_);
  nor (_08730_, _08255_, _07530_);
  nor (_08731_, _08255_, \oc8051_golden_model_1.ACC [5]);
  and (_08732_, _08255_, \oc8051_golden_model_1.ACC [5]);
  nor (_08733_, _08732_, _08731_);
  nor (_08734_, _08269_, _07536_);
  and (_08735_, _08269_, \oc8051_golden_model_1.ACC [4]);
  nor (_08736_, _08269_, \oc8051_golden_model_1.ACC [4]);
  nor (_08737_, _08736_, _08735_);
  not (_08738_, _08737_);
  nor (_08739_, _08208_, _07634_);
  and (_08740_, _08208_, \oc8051_golden_model_1.ACC [2]);
  nor (_08741_, _08208_, \oc8051_golden_model_1.ACC [2]);
  nor (_08742_, _08741_, _08740_);
  nor (_08743_, _08223_, _03320_);
  nor (_08744_, _08223_, \oc8051_golden_model_1.ACC [1]);
  and (_08745_, _08223_, \oc8051_golden_model_1.ACC [1]);
  nor (_08746_, _08745_, _08744_);
  nor (_08747_, _08238_, _03397_);
  not (_08748_, _08747_);
  nor (_08749_, _08748_, _08746_);
  nor (_08750_, _08749_, _08743_);
  nor (_08751_, _08750_, _08742_);
  nor (_08752_, _08751_, _08739_);
  nor (_08753_, _08752_, _08191_);
  or (_08754_, _08753_, \oc8051_golden_model_1.ACC [3]);
  nand (_08755_, _08752_, _08191_);
  and (_08756_, _08755_, _08754_);
  and (_08757_, _08756_, _08738_);
  nor (_08758_, _08757_, _08734_);
  nor (_08759_, _08758_, _08733_);
  nor (_08760_, _08759_, _08730_);
  nor (_08761_, _08760_, _08729_);
  nor (_08762_, _08761_, _08726_);
  nor (_08763_, _08762_, _08725_);
  and (_08764_, _08762_, _08725_);
  or (_08765_, _08764_, _08763_);
  or (_08766_, _08765_, _08720_);
  and (_08767_, _08766_, _08722_);
  or (_08768_, _08767_, _08719_);
  and (_08769_, _03648_, _03245_);
  not (_08770_, _08769_);
  not (_08771_, _08720_);
  nor (_08772_, _03556_, _07484_);
  and (_08773_, _03556_, _07484_);
  or (_08774_, _08773_, _08772_);
  not (_08775_, _08774_);
  nor (_08776_, _03853_, _07530_);
  and (_08777_, _03853_, _07530_);
  nor (_08778_, _04308_, _07536_);
  and (_08779_, _04308_, _07536_);
  nor (_08780_, _08779_, _08778_);
  nor (_08781_, _03494_, _07628_);
  and (_08782_, _03494_, _07628_);
  nor (_08783_, _03898_, _07634_);
  and (_08784_, _03898_, _07634_);
  nor (_08785_, _08784_, _08783_);
  not (_08786_, _08785_);
  nor (_08787_, _04042_, _03397_);
  and (_08788_, _08787_, _08383_);
  nor (_08789_, _08788_, _08381_);
  nor (_08790_, _08789_, _08786_);
  nor (_08791_, _08790_, _08783_);
  nor (_08792_, _08791_, _08782_);
  or (_08793_, _08792_, _08781_);
  and (_08794_, _08793_, _08780_);
  nor (_08795_, _08794_, _08778_);
  nor (_08796_, _08795_, _08777_);
  or (_08797_, _08796_, _08776_);
  and (_08798_, _08797_, _08775_);
  nor (_08799_, _08798_, _08772_);
  nor (_08800_, _08799_, _08479_);
  and (_08801_, _08799_, _08479_);
  or (_08802_, _08801_, _08800_);
  or (_08803_, _08802_, _08771_);
  and (_08804_, _08803_, _08770_);
  and (_08805_, _08804_, _08768_);
  and (_08806_, _08769_, \oc8051_golden_model_1.ACC [6]);
  or (_08807_, _08806_, _03809_);
  or (_08808_, _08807_, _08805_);
  and (_08809_, _03675_, _03066_);
  not (_08810_, _08809_);
  nand (_08811_, _08065_, _03809_);
  and (_08812_, _08811_, _08810_);
  and (_08813_, _08812_, _08808_);
  and (_08814_, _03648_, _03066_);
  nor (_08815_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08816_, _08815_, _07577_);
  and (_08817_, _08816_, _07500_);
  and (_08818_, _08817_, _07484_);
  nor (_08819_, _08818_, _06061_);
  and (_08820_, _08818_, _06061_);
  nor (_08821_, _08820_, _08819_);
  nor (_08822_, _08821_, _08810_);
  or (_08823_, _08822_, _08814_);
  or (_08824_, _08823_, _08813_);
  nand (_08825_, _08814_, _07911_);
  and (_08826_, _08825_, _03206_);
  and (_08827_, _08826_, _08824_);
  nor (_08828_, _08114_, _03206_);
  or (_08829_, _08828_, _03816_);
  or (_08830_, _08829_, _08827_);
  and (_08831_, _03675_, _03241_);
  not (_08832_, _08831_);
  and (_08833_, _05895_, _05371_);
  nor (_08834_, _08833_, _07937_);
  nand (_08835_, _08834_, _03816_);
  and (_08836_, _08835_, _08832_);
  and (_08837_, _08836_, _08830_);
  and (_08838_, _03648_, _03241_);
  and (_08839_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08840_, _08839_, _07578_);
  nor (_08841_, _08840_, _07536_);
  and (_08842_, _08841_, \oc8051_golden_model_1.ACC [5]);
  and (_08843_, _08842_, \oc8051_golden_model_1.ACC [6]);
  nor (_08844_, _08843_, \oc8051_golden_model_1.ACC [7]);
  and (_08845_, _08843_, \oc8051_golden_model_1.ACC [7]);
  nor (_08846_, _08845_, _08844_);
  and (_08847_, _08846_, _08831_);
  or (_08848_, _08847_, _08838_);
  or (_08849_, _08848_, _08837_);
  nand (_08850_, _08838_, _03397_);
  and (_08851_, _08850_, _43227_);
  and (_08852_, _08851_, _08849_);
  or (_08853_, _08852_, _07855_);
  and (_40746_, _08853_, _41991_);
  not (_08854_, \oc8051_golden_model_1.DPL [7]);
  nor (_08855_, _43227_, _08854_);
  nor (_08856_, _05319_, _08854_);
  not (_08857_, _05319_);
  nor (_08858_, _06457_, _08857_);
  or (_08859_, _08858_, _08856_);
  and (_08860_, _08859_, _03786_);
  not (_08861_, _03651_);
  nor (_08862_, _08857_, _05289_);
  or (_08863_, _08862_, _08856_);
  or (_08864_, _08863_, _06889_);
  not (_08865_, _03656_);
  and (_08866_, _06185_, _05319_);
  or (_08867_, _08866_, _08856_);
  or (_08868_, _08867_, _04515_);
  and (_08869_, _05319_, \oc8051_golden_model_1.ACC [7]);
  or (_08870_, _08869_, _08856_);
  and (_08871_, _08870_, _04499_);
  nor (_08872_, _04499_, _08854_);
  or (_08873_, _08872_, _03599_);
  or (_08874_, _08873_, _08871_);
  and (_08875_, _08874_, _04524_);
  and (_08876_, _08875_, _08868_);
  and (_08877_, _08863_, _03597_);
  or (_08878_, _08877_, _03603_);
  or (_08879_, _08878_, _08876_);
  nor (_08880_, _03284_, _03264_);
  not (_08881_, _08880_);
  or (_08882_, _08870_, _03611_);
  and (_08883_, _08882_, _08881_);
  and (_08884_, _08883_, _08879_);
  and (_08885_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_08886_, _08885_, \oc8051_golden_model_1.DPL [2]);
  and (_08887_, _08886_, \oc8051_golden_model_1.DPL [3]);
  and (_08888_, _08887_, \oc8051_golden_model_1.DPL [4]);
  and (_08889_, _08888_, \oc8051_golden_model_1.DPL [5]);
  and (_08890_, _08889_, \oc8051_golden_model_1.DPL [6]);
  nor (_08891_, _08890_, \oc8051_golden_model_1.DPL [7]);
  and (_08892_, _08890_, \oc8051_golden_model_1.DPL [7]);
  nor (_08893_, _08892_, _08891_);
  and (_08894_, _08893_, _08880_);
  or (_08895_, _08894_, _08884_);
  and (_08896_, _08895_, _08865_);
  nor (_08897_, _05958_, _08865_);
  or (_08898_, _08897_, _07441_);
  or (_08899_, _08898_, _08896_);
  and (_08900_, _08899_, _08864_);
  or (_08901_, _08900_, _05969_);
  and (_08902_, _06171_, _05319_);
  or (_08903_, _08856_, _05970_);
  or (_08904_, _08903_, _08902_);
  and (_08905_, _08904_, _03275_);
  and (_08906_, _08905_, _08901_);
  nor (_08907_, _06443_, _08857_);
  or (_08908_, _08907_, _08856_);
  and (_08909_, _08908_, _03644_);
  or (_08910_, _08909_, _08906_);
  or (_08911_, _08910_, _08861_);
  and (_08912_, _05961_, _05319_);
  or (_08913_, _08856_, _04591_);
  or (_08914_, _08913_, _08912_);
  and (_08915_, _06247_, _05319_);
  or (_08916_, _08915_, _08856_);
  or (_08917_, _08916_, _04582_);
  and (_08918_, _08917_, _04589_);
  and (_08919_, _08918_, _08914_);
  and (_08920_, _08919_, _08911_);
  and (_08922_, _06458_, _05319_);
  or (_08923_, _08922_, _08856_);
  and (_08924_, _08923_, _03778_);
  or (_08925_, _08924_, _08920_);
  and (_08926_, _08925_, _04596_);
  or (_08927_, _08856_, _05397_);
  and (_08928_, _08916_, _03655_);
  and (_08929_, _08928_, _08927_);
  or (_08930_, _08929_, _08926_);
  and (_08931_, _08930_, _04594_);
  and (_08933_, _08870_, _03773_);
  and (_08934_, _08933_, _08927_);
  or (_08935_, _08934_, _03653_);
  or (_08936_, _08935_, _08931_);
  nor (_08937_, _05959_, _08857_);
  or (_08938_, _08856_, _04608_);
  or (_08939_, _08938_, _08937_);
  and (_08940_, _08939_, _04606_);
  and (_08941_, _08940_, _08936_);
  or (_08942_, _08941_, _08860_);
  and (_08944_, _08942_, _04260_);
  and (_08945_, _08867_, _03809_);
  or (_08946_, _08945_, _03816_);
  or (_08947_, _08946_, _08944_);
  and (_08948_, _05895_, _05319_);
  or (_08949_, _08856_, _03820_);
  or (_08950_, _08949_, _08948_);
  and (_08951_, _08950_, _43227_);
  and (_08952_, _08951_, _08947_);
  or (_08953_, _08952_, _08855_);
  and (_40747_, _08953_, _41991_);
  not (_08955_, \oc8051_golden_model_1.DPH [7]);
  nor (_08956_, _43227_, _08955_);
  nor (_08957_, _05297_, _08955_);
  not (_08958_, _05297_);
  nor (_08959_, _06457_, _08958_);
  or (_08960_, _08959_, _08957_);
  and (_08961_, _08960_, _03786_);
  nor (_08962_, _08958_, _05289_);
  or (_08963_, _08962_, _08957_);
  or (_08965_, _08963_, _06889_);
  and (_08966_, _06185_, _05297_);
  or (_08967_, _08966_, _08957_);
  or (_08968_, _08967_, _04515_);
  and (_08969_, _05297_, \oc8051_golden_model_1.ACC [7]);
  or (_08970_, _08969_, _08957_);
  and (_08971_, _08970_, _04499_);
  nor (_08972_, _04499_, _08955_);
  or (_08973_, _08972_, _03599_);
  or (_08974_, _08973_, _08971_);
  and (_08976_, _08974_, _04524_);
  and (_08977_, _08976_, _08968_);
  and (_08978_, _08963_, _03597_);
  or (_08979_, _08978_, _03603_);
  or (_08980_, _08979_, _08977_);
  or (_08981_, _08970_, _03611_);
  and (_08982_, _08981_, _08881_);
  and (_08983_, _08982_, _08980_);
  and (_08984_, \oc8051_golden_model_1.DPH [1], \oc8051_golden_model_1.DPH [0]);
  and (_08985_, _08984_, _08892_);
  and (_08987_, _08985_, \oc8051_golden_model_1.DPH [2]);
  and (_08988_, _08987_, \oc8051_golden_model_1.DPH [3]);
  and (_08989_, _08988_, \oc8051_golden_model_1.DPH [4]);
  and (_08990_, _08989_, \oc8051_golden_model_1.DPH [5]);
  nand (_08991_, _08990_, \oc8051_golden_model_1.DPH [6]);
  or (_08992_, _08991_, _08955_);
  nand (_08993_, _08991_, _08955_);
  and (_08994_, _08993_, _08880_);
  and (_08995_, _08994_, _08992_);
  or (_08996_, _08995_, _08983_);
  and (_08997_, _08996_, _08865_);
  and (_08998_, _03656_, _03463_);
  or (_08999_, _08998_, _07441_);
  or (_09000_, _08999_, _08997_);
  and (_09001_, _09000_, _08965_);
  or (_09002_, _09001_, _05969_);
  and (_09003_, _06171_, _05297_);
  or (_09004_, _08957_, _05970_);
  or (_09005_, _09004_, _09003_);
  and (_09006_, _09005_, _03275_);
  and (_09007_, _09006_, _09002_);
  nor (_09008_, _06443_, _08958_);
  or (_09009_, _09008_, _08957_);
  and (_09010_, _09009_, _03644_);
  or (_09011_, _09010_, _09007_);
  or (_09012_, _09011_, _08861_);
  and (_09013_, _05961_, _05297_);
  or (_09014_, _08957_, _04591_);
  or (_09015_, _09014_, _09013_);
  and (_09016_, _06247_, _05297_);
  or (_09017_, _09016_, _08957_);
  or (_09018_, _09017_, _04582_);
  and (_09019_, _09018_, _04589_);
  and (_09020_, _09019_, _09015_);
  and (_09021_, _09020_, _09012_);
  and (_09022_, _06458_, _05297_);
  or (_09023_, _09022_, _08957_);
  and (_09024_, _09023_, _03778_);
  or (_09025_, _09024_, _09021_);
  and (_09026_, _09025_, _04596_);
  or (_09027_, _08957_, _05397_);
  and (_09028_, _09017_, _03655_);
  and (_09029_, _09028_, _09027_);
  or (_09030_, _09029_, _09026_);
  and (_09031_, _09030_, _04594_);
  and (_09032_, _08970_, _03773_);
  and (_09033_, _09032_, _09027_);
  or (_09034_, _09033_, _03653_);
  or (_09035_, _09034_, _09031_);
  nor (_09036_, _05959_, _08958_);
  or (_09037_, _08957_, _04608_);
  or (_09038_, _09037_, _09036_);
  and (_09039_, _09038_, _04606_);
  and (_09040_, _09039_, _09035_);
  or (_09041_, _09040_, _08961_);
  and (_09042_, _09041_, _04260_);
  and (_09043_, _08967_, _03809_);
  or (_09044_, _09043_, _03816_);
  or (_09045_, _09044_, _09042_);
  and (_09046_, _05895_, _05297_);
  or (_09047_, _08957_, _03820_);
  or (_09048_, _09047_, _09046_);
  and (_09049_, _09048_, _43227_);
  and (_09050_, _09049_, _09045_);
  or (_09051_, _09050_, _08956_);
  and (_40748_, _09051_, _41991_);
  not (_09052_, \oc8051_golden_model_1.IE [7]);
  nor (_09053_, _05337_, _09052_);
  not (_09054_, _05337_);
  nor (_09055_, _09054_, _05289_);
  nor (_09056_, _09055_, _09053_);
  and (_09057_, _09056_, _07441_);
  nor (_09058_, _05979_, _09052_);
  and (_09059_, _06038_, _05979_);
  nor (_09060_, _09059_, _09058_);
  nor (_09061_, _09060_, _03512_);
  and (_09062_, _05337_, \oc8051_golden_model_1.ACC [7]);
  nor (_09063_, _09062_, _09053_);
  nor (_09064_, _09063_, _04500_);
  nor (_09065_, _04499_, _09052_);
  or (_09066_, _09065_, _09064_);
  and (_09067_, _09066_, _04515_);
  and (_09068_, _06185_, _05337_);
  nor (_09069_, _09068_, _09053_);
  nor (_09070_, _09069_, _04515_);
  or (_09071_, _09070_, _09067_);
  and (_09072_, _09071_, _03516_);
  and (_09073_, _06042_, _05979_);
  nor (_09074_, _09073_, _09058_);
  nor (_09075_, _09074_, _03516_);
  or (_09076_, _09075_, _03597_);
  or (_09077_, _09076_, _09072_);
  nand (_09078_, _09056_, _03597_);
  and (_09079_, _09078_, _09077_);
  and (_09080_, _09079_, _03611_);
  nor (_09081_, _09063_, _03611_);
  or (_09082_, _09081_, _09080_);
  and (_09083_, _09082_, _03512_);
  nor (_09084_, _09083_, _09061_);
  nor (_09085_, _09084_, _03504_);
  nor (_09086_, _09058_, _06216_);
  or (_09087_, _09074_, _03505_);
  nor (_09088_, _09087_, _09086_);
  nor (_09089_, _09088_, _09085_);
  nor (_09090_, _09089_, _03500_);
  not (_09091_, _05979_);
  nor (_09092_, _06026_, _09091_);
  nor (_09093_, _09092_, _09058_);
  nor (_09094_, _09093_, _03501_);
  nor (_09095_, _09094_, _07441_);
  not (_09096_, _09095_);
  nor (_09097_, _09096_, _09090_);
  nor (_09098_, _09097_, _09057_);
  nor (_09099_, _09098_, _05969_);
  and (_09100_, _06171_, _05337_);
  nor (_09101_, _09053_, _05970_);
  not (_09102_, _09101_);
  nor (_09103_, _09102_, _09100_);
  nor (_09104_, _09103_, _03644_);
  not (_09105_, _09104_);
  nor (_09106_, _09105_, _09099_);
  nor (_09107_, _06443_, _09054_);
  nor (_09108_, _09107_, _09053_);
  nor (_09109_, _09108_, _03275_);
  or (_09110_, _09109_, _08861_);
  or (_09111_, _09110_, _09106_);
  and (_09112_, _05961_, _05337_);
  or (_09113_, _09053_, _04591_);
  or (_09114_, _09113_, _09112_);
  and (_09115_, _06247_, _05337_);
  nor (_09116_, _09115_, _09053_);
  and (_09117_, _09116_, _03650_);
  nor (_09118_, _09117_, _03778_);
  and (_09119_, _09118_, _09114_);
  and (_09120_, _09119_, _09111_);
  and (_09121_, _06458_, _05337_);
  nor (_09122_, _09121_, _09053_);
  nor (_09123_, _09122_, _04589_);
  nor (_09124_, _09123_, _09120_);
  nor (_09125_, _09124_, _03655_);
  nor (_09126_, _09053_, _05397_);
  not (_09127_, _09126_);
  nor (_09128_, _09116_, _04596_);
  and (_09129_, _09128_, _09127_);
  nor (_09130_, _09129_, _09125_);
  nor (_09131_, _09130_, _03773_);
  nor (_09132_, _09063_, _04594_);
  and (_09133_, _09132_, _09127_);
  or (_09134_, _09133_, _09131_);
  and (_09135_, _09134_, _04608_);
  nor (_09136_, _05959_, _09054_);
  nor (_09137_, _09136_, _09053_);
  nor (_09138_, _09137_, _04608_);
  or (_09139_, _09138_, _09135_);
  and (_09140_, _09139_, _04606_);
  nor (_09141_, _06457_, _09054_);
  nor (_09142_, _09141_, _09053_);
  nor (_09143_, _09142_, _04606_);
  or (_09144_, _09143_, _09140_);
  and (_09145_, _09144_, _04260_);
  nor (_09146_, _09069_, _04260_);
  or (_09147_, _09146_, _09145_);
  and (_09148_, _09147_, _03206_);
  nor (_09149_, _09060_, _03206_);
  or (_09150_, _09149_, _09148_);
  and (_09151_, _09150_, _03820_);
  and (_09152_, _05895_, _05337_);
  nor (_09153_, _09152_, _09053_);
  nor (_09154_, _09153_, _03820_);
  or (_09155_, _09154_, _09151_);
  or (_09156_, _09155_, _43231_);
  or (_09157_, _43227_, \oc8051_golden_model_1.IE [7]);
  and (_09158_, _09157_, _41991_);
  and (_40750_, _09158_, _09156_);
  not (_09159_, \oc8051_golden_model_1.IP [7]);
  nor (_09160_, _05376_, _09159_);
  not (_09161_, _05376_);
  nor (_09162_, _09161_, _05289_);
  nor (_09163_, _09162_, _09160_);
  and (_09164_, _09163_, _07441_);
  nor (_09165_, _05989_, _09159_);
  and (_09166_, _06038_, _05989_);
  nor (_09167_, _09166_, _09165_);
  nor (_09168_, _09167_, _03512_);
  and (_09169_, _05376_, \oc8051_golden_model_1.ACC [7]);
  nor (_09170_, _09169_, _09160_);
  nor (_09171_, _09170_, _04500_);
  nor (_09172_, _04499_, _09159_);
  or (_09173_, _09172_, _09171_);
  and (_09174_, _09173_, _04515_);
  and (_09175_, _06185_, _05376_);
  nor (_09176_, _09175_, _09160_);
  nor (_09177_, _09176_, _04515_);
  or (_09178_, _09177_, _09174_);
  and (_09179_, _09178_, _03516_);
  and (_09180_, _06042_, _05989_);
  nor (_09181_, _09180_, _09165_);
  nor (_09182_, _09181_, _03516_);
  or (_09183_, _09182_, _03597_);
  or (_09184_, _09183_, _09179_);
  nand (_09185_, _09163_, _03597_);
  and (_09186_, _09185_, _09184_);
  and (_09187_, _09186_, _03611_);
  nor (_09188_, _09170_, _03611_);
  or (_09189_, _09188_, _09187_);
  and (_09190_, _09189_, _03512_);
  nor (_09191_, _09190_, _09168_);
  nor (_09192_, _09191_, _03504_);
  nor (_09193_, _09165_, _06216_);
  or (_09194_, _09181_, _03505_);
  nor (_09195_, _09194_, _09193_);
  nor (_09196_, _09195_, _09192_);
  nor (_09197_, _09196_, _03500_);
  not (_09198_, _05989_);
  nor (_09199_, _06026_, _09198_);
  nor (_09200_, _09199_, _09165_);
  nor (_09201_, _09200_, _03501_);
  nor (_09202_, _09201_, _07441_);
  not (_09203_, _09202_);
  nor (_09204_, _09203_, _09197_);
  nor (_09205_, _09204_, _09164_);
  nor (_09206_, _09205_, _05969_);
  and (_09207_, _06171_, _05376_);
  nor (_09208_, _09160_, _05970_);
  not (_09209_, _09208_);
  nor (_09210_, _09209_, _09207_);
  nor (_09211_, _09210_, _03644_);
  not (_09212_, _09211_);
  nor (_09213_, _09212_, _09206_);
  nor (_09214_, _06443_, _09161_);
  nor (_09215_, _09214_, _09160_);
  nor (_09216_, _09215_, _03275_);
  or (_09217_, _09216_, _08861_);
  or (_09218_, _09217_, _09213_);
  and (_09219_, _05961_, _05376_);
  or (_09220_, _09160_, _04591_);
  or (_09221_, _09220_, _09219_);
  and (_09222_, _06247_, _05376_);
  nor (_09223_, _09222_, _09160_);
  and (_09224_, _09223_, _03650_);
  nor (_09225_, _09224_, _03778_);
  and (_09226_, _09225_, _09221_);
  and (_09227_, _09226_, _09218_);
  and (_09228_, _06458_, _05376_);
  nor (_09229_, _09228_, _09160_);
  nor (_09230_, _09229_, _04589_);
  nor (_09231_, _09230_, _09227_);
  nor (_09232_, _09231_, _03655_);
  nor (_09233_, _09160_, _05397_);
  not (_09234_, _09233_);
  nor (_09235_, _09223_, _04596_);
  and (_09236_, _09235_, _09234_);
  nor (_09237_, _09236_, _09232_);
  nor (_09238_, _09237_, _03773_);
  nor (_09239_, _09170_, _04594_);
  and (_09240_, _09239_, _09234_);
  or (_09241_, _09240_, _09238_);
  and (_09242_, _09241_, _04608_);
  nor (_09243_, _05959_, _09161_);
  nor (_09244_, _09243_, _09160_);
  nor (_09245_, _09244_, _04608_);
  or (_09246_, _09245_, _09242_);
  and (_09247_, _09246_, _04606_);
  nor (_09248_, _06457_, _09161_);
  nor (_09249_, _09248_, _09160_);
  nor (_09250_, _09249_, _04606_);
  or (_09251_, _09250_, _09247_);
  and (_09252_, _09251_, _04260_);
  nor (_09253_, _09176_, _04260_);
  or (_09254_, _09253_, _09252_);
  and (_09255_, _09254_, _03206_);
  nor (_09256_, _09167_, _03206_);
  or (_09257_, _09256_, _09255_);
  and (_09258_, _09257_, _03820_);
  and (_09259_, _05895_, _05376_);
  nor (_09260_, _09259_, _09160_);
  nor (_09261_, _09260_, _03820_);
  or (_09262_, _09261_, _09258_);
  or (_09263_, _09262_, _43231_);
  or (_09264_, _43227_, \oc8051_golden_model_1.IP [7]);
  and (_09265_, _09264_, _41991_);
  and (_40751_, _09265_, _09263_);
  not (_09266_, \oc8051_golden_model_1.P0 [7]);
  nor (_09267_, _05363_, _09266_);
  not (_09268_, _05363_);
  nor (_09269_, _09268_, _05289_);
  or (_09270_, _09269_, _09267_);
  or (_09271_, _09270_, _06889_);
  nor (_09272_, _05294_, _09266_);
  and (_09273_, _06038_, _05294_);
  or (_09274_, _09273_, _09272_);
  and (_09275_, _09274_, _03511_);
  and (_09276_, _06185_, _05363_);
  or (_09277_, _09276_, _09267_);
  or (_09278_, _09277_, _04515_);
  and (_09279_, _05363_, \oc8051_golden_model_1.ACC [7]);
  or (_09280_, _09279_, _09267_);
  and (_09281_, _09280_, _04499_);
  nor (_09282_, _04499_, _09266_);
  or (_09283_, _09282_, _03599_);
  or (_09284_, _09283_, _09281_);
  and (_09285_, _09284_, _03516_);
  and (_09286_, _09285_, _09278_);
  and (_09287_, _06042_, _05294_);
  or (_09288_, _09287_, _09272_);
  and (_09289_, _09288_, _03515_);
  or (_09290_, _09289_, _03597_);
  or (_09291_, _09290_, _09286_);
  or (_09292_, _09270_, _04524_);
  and (_09293_, _09292_, _09291_);
  or (_09294_, _09293_, _03603_);
  or (_09295_, _09280_, _03611_);
  and (_09296_, _09295_, _03512_);
  and (_09297_, _09296_, _09294_);
  or (_09298_, _09297_, _09275_);
  and (_09299_, _09298_, _03505_);
  or (_09300_, _09272_, _06216_);
  and (_09301_, _09300_, _03504_);
  and (_09302_, _09301_, _09288_);
  or (_09303_, _09302_, _09299_);
  and (_09304_, _09303_, _03501_);
  or (_09305_, _06038_, _06025_);
  and (_09306_, _09305_, _05294_);
  or (_09307_, _09306_, _09272_);
  and (_09308_, _09307_, _03500_);
  or (_09309_, _09308_, _07441_);
  or (_09310_, _09309_, _09304_);
  and (_09311_, _09310_, _09271_);
  or (_09312_, _09311_, _05969_);
  and (_09313_, _06171_, _05363_);
  or (_09314_, _09267_, _05970_);
  or (_09315_, _09314_, _09313_);
  and (_09316_, _09315_, _03275_);
  and (_09317_, _09316_, _09312_);
  and (_09318_, _06356_, \oc8051_golden_model_1.P0 [7]);
  and (_09319_, _06361_, \oc8051_golden_model_1.P2 [7]);
  or (_09320_, _09319_, _06351_);
  or (_09321_, _09320_, _09318_);
  and (_09322_, _06378_, \oc8051_golden_model_1.P1 [7]);
  and (_09323_, _06382_, \oc8051_golden_model_1.P3 [7]);
  or (_09324_, _09323_, _09322_);
  or (_09325_, _09324_, _06373_);
  or (_09326_, _09325_, _06369_);
  nor (_09327_, _09326_, _09321_);
  and (_09328_, _09327_, _06407_);
  nand (_09329_, _09328_, _06440_);
  or (_09330_, _09329_, _06248_);
  and (_09331_, _09330_, _05363_);
  or (_09332_, _09331_, _09267_);
  and (_09333_, _09332_, _03644_);
  or (_09334_, _09333_, _08861_);
  or (_09335_, _09334_, _09317_);
  and (_09336_, _05961_, _05363_);
  or (_09337_, _09267_, _04591_);
  or (_09338_, _09337_, _09336_);
  and (_09339_, _06247_, _05363_);
  or (_09340_, _09339_, _09267_);
  or (_09341_, _09340_, _04582_);
  and (_09342_, _09341_, _04589_);
  and (_09343_, _09342_, _09338_);
  and (_09344_, _09343_, _09335_);
  and (_09345_, _06458_, _05363_);
  or (_09346_, _09345_, _09267_);
  and (_09347_, _09346_, _03778_);
  or (_09348_, _09347_, _09344_);
  and (_09349_, _09348_, _04596_);
  or (_09350_, _09267_, _05397_);
  and (_09351_, _09340_, _03655_);
  and (_09352_, _09351_, _09350_);
  or (_09353_, _09352_, _09349_);
  and (_09354_, _09353_, _04594_);
  and (_09355_, _09280_, _03773_);
  and (_09356_, _09355_, _09350_);
  or (_09357_, _09356_, _03653_);
  or (_09358_, _09357_, _09354_);
  nor (_09359_, _05959_, _09268_);
  or (_09360_, _09267_, _04608_);
  or (_09361_, _09360_, _09359_);
  and (_09362_, _09361_, _04606_);
  and (_09363_, _09362_, _09358_);
  nor (_09364_, _06457_, _09268_);
  or (_09365_, _09364_, _09267_);
  and (_09366_, _09365_, _03786_);
  or (_09367_, _09366_, _03809_);
  or (_09368_, _09367_, _09363_);
  or (_09369_, _09277_, _04260_);
  and (_09370_, _09369_, _03206_);
  and (_09371_, _09370_, _09368_);
  and (_09372_, _09274_, _03205_);
  or (_09373_, _09372_, _03816_);
  or (_09374_, _09373_, _09371_);
  and (_09375_, _05895_, _05363_);
  or (_09376_, _09267_, _03820_);
  or (_09377_, _09376_, _09375_);
  and (_09378_, _09377_, _43227_);
  and (_09379_, _09378_, _09374_);
  nor (_09380_, _43227_, _09266_);
  or (_09381_, _09380_, rst);
  or (_40752_, _09381_, _09379_);
  not (_09382_, \oc8051_golden_model_1.P1 [7]);
  nor (_09383_, _43227_, _09382_);
  or (_09384_, _09383_, rst);
  nor (_09385_, _05383_, _09382_);
  not (_09386_, _05383_);
  nor (_09387_, _09386_, _05289_);
  or (_09388_, _09387_, _09385_);
  or (_09389_, _09388_, _06889_);
  nor (_09390_, _06013_, _09382_);
  and (_09391_, _06038_, _06013_);
  or (_09392_, _09391_, _09390_);
  and (_09393_, _09392_, _03511_);
  and (_09394_, _06185_, _05383_);
  or (_09395_, _09394_, _09385_);
  or (_09396_, _09395_, _04515_);
  and (_09397_, _05383_, \oc8051_golden_model_1.ACC [7]);
  or (_09398_, _09397_, _09385_);
  and (_09399_, _09398_, _04499_);
  nor (_09400_, _04499_, _09382_);
  or (_09401_, _09400_, _03599_);
  or (_09402_, _09401_, _09399_);
  and (_09403_, _09402_, _03516_);
  and (_09404_, _09403_, _09396_);
  and (_09405_, _06042_, _06013_);
  or (_09406_, _09405_, _09390_);
  and (_09407_, _09406_, _03515_);
  or (_09408_, _09407_, _03597_);
  or (_09409_, _09408_, _09404_);
  or (_09410_, _09388_, _04524_);
  and (_09411_, _09410_, _09409_);
  or (_09412_, _09411_, _03603_);
  or (_09413_, _09398_, _03611_);
  and (_09414_, _09413_, _03512_);
  and (_09415_, _09414_, _09412_);
  or (_09416_, _09415_, _09393_);
  and (_09417_, _09416_, _03505_);
  and (_09418_, _06217_, _06013_);
  or (_09419_, _09418_, _09390_);
  and (_09420_, _09419_, _03504_);
  or (_09421_, _09420_, _09417_);
  and (_09422_, _09421_, _03501_);
  and (_09423_, _09305_, _06013_);
  or (_09424_, _09423_, _09390_);
  and (_09425_, _09424_, _03500_);
  or (_09426_, _09425_, _07441_);
  or (_09427_, _09426_, _09422_);
  and (_09428_, _09427_, _09389_);
  or (_09429_, _09428_, _05969_);
  and (_09430_, _06171_, _05383_);
  or (_09431_, _09385_, _05970_);
  or (_09432_, _09431_, _09430_);
  and (_09433_, _09432_, _03275_);
  and (_09434_, _09433_, _09429_);
  and (_09435_, _09330_, _05383_);
  or (_09436_, _09435_, _09385_);
  and (_09437_, _09436_, _03644_);
  or (_09438_, _09437_, _08861_);
  or (_09439_, _09438_, _09434_);
  and (_09440_, _05961_, _05383_);
  or (_09441_, _09385_, _04591_);
  or (_09442_, _09441_, _09440_);
  and (_09443_, _06247_, _05383_);
  or (_09444_, _09443_, _09385_);
  or (_09445_, _09444_, _04582_);
  and (_09446_, _09445_, _04589_);
  and (_09447_, _09446_, _09442_);
  and (_09448_, _09447_, _09439_);
  and (_09449_, _06458_, _05383_);
  or (_09450_, _09449_, _09385_);
  and (_09451_, _09450_, _03778_);
  or (_09452_, _09451_, _09448_);
  and (_09453_, _09452_, _04596_);
  or (_09454_, _09385_, _05397_);
  and (_09455_, _09444_, _03655_);
  and (_09456_, _09455_, _09454_);
  or (_09457_, _09456_, _09453_);
  and (_09458_, _09457_, _04594_);
  and (_09459_, _09398_, _03773_);
  and (_09460_, _09459_, _09454_);
  or (_09461_, _09460_, _03653_);
  or (_09462_, _09461_, _09458_);
  nor (_09463_, _05959_, _09386_);
  or (_09464_, _09385_, _04608_);
  or (_09465_, _09464_, _09463_);
  and (_09466_, _09465_, _04606_);
  and (_09467_, _09466_, _09462_);
  nor (_09468_, _06457_, _09386_);
  or (_09469_, _09468_, _09385_);
  and (_09470_, _09469_, _03786_);
  or (_09471_, _09470_, _03809_);
  or (_09472_, _09471_, _09467_);
  or (_09473_, _09395_, _04260_);
  and (_09474_, _09473_, _03206_);
  and (_09475_, _09474_, _09472_);
  and (_09476_, _09392_, _03205_);
  or (_09477_, _09476_, _03816_);
  or (_09478_, _09477_, _09475_);
  and (_09479_, _05895_, _05383_);
  or (_09480_, _09385_, _03820_);
  or (_09481_, _09480_, _09479_);
  and (_09482_, _09481_, _43227_);
  and (_09483_, _09482_, _09478_);
  or (_40753_, _09483_, _09384_);
  not (_09484_, \oc8051_golden_model_1.P2 [7]);
  nor (_09485_, _05386_, _09484_);
  not (_09486_, _05386_);
  nor (_09487_, _09486_, _05289_);
  or (_09488_, _09487_, _09485_);
  or (_09489_, _09488_, _06889_);
  nor (_09490_, _06009_, _09484_);
  and (_09491_, _06038_, _06009_);
  or (_09492_, _09491_, _09490_);
  and (_09493_, _09492_, _03511_);
  and (_09494_, _06185_, _05386_);
  or (_09495_, _09494_, _09485_);
  or (_09496_, _09495_, _04515_);
  and (_09497_, _05386_, \oc8051_golden_model_1.ACC [7]);
  or (_09498_, _09497_, _09485_);
  and (_09499_, _09498_, _04499_);
  nor (_09500_, _04499_, _09484_);
  or (_09501_, _09500_, _03599_);
  or (_09502_, _09501_, _09499_);
  and (_09503_, _09502_, _03516_);
  and (_09504_, _09503_, _09496_);
  and (_09505_, _06042_, _06009_);
  or (_09506_, _09505_, _09490_);
  and (_09507_, _09506_, _03515_);
  or (_09508_, _09507_, _03597_);
  or (_09509_, _09508_, _09504_);
  or (_09510_, _09488_, _04524_);
  and (_09511_, _09510_, _09509_);
  or (_09512_, _09511_, _03603_);
  or (_09513_, _09498_, _03611_);
  and (_09514_, _09513_, _03512_);
  and (_09515_, _09514_, _09512_);
  or (_09516_, _09515_, _09493_);
  and (_09517_, _09516_, _03505_);
  and (_09518_, _06217_, _06009_);
  or (_09519_, _09518_, _09490_);
  and (_09520_, _09519_, _03504_);
  or (_09521_, _09520_, _09517_);
  and (_09522_, _09521_, _03501_);
  and (_09523_, _09305_, _06009_);
  or (_09524_, _09523_, _09490_);
  and (_09525_, _09524_, _03500_);
  or (_09526_, _09525_, _07441_);
  or (_09527_, _09526_, _09522_);
  and (_09528_, _09527_, _09489_);
  or (_09529_, _09528_, _05969_);
  and (_09530_, _06171_, _05386_);
  or (_09531_, _09485_, _05970_);
  or (_09533_, _09531_, _09530_);
  and (_09534_, _09533_, _03275_);
  and (_09535_, _09534_, _09529_);
  and (_09536_, _09330_, _05386_);
  or (_09537_, _09536_, _09485_);
  and (_09538_, _09537_, _03644_);
  or (_09539_, _09538_, _08861_);
  or (_09540_, _09539_, _09535_);
  and (_09541_, _05961_, _05386_);
  or (_09542_, _09485_, _04591_);
  or (_09543_, _09542_, _09541_);
  and (_09544_, _06247_, _05386_);
  or (_09545_, _09544_, _09485_);
  or (_09546_, _09545_, _04582_);
  and (_09547_, _09546_, _04589_);
  and (_09548_, _09547_, _09543_);
  and (_09549_, _09548_, _09540_);
  and (_09550_, _06458_, _05386_);
  or (_09551_, _09550_, _09485_);
  and (_09552_, _09551_, _03778_);
  or (_09554_, _09552_, _09549_);
  and (_09555_, _09554_, _04596_);
  or (_09556_, _09485_, _05397_);
  and (_09557_, _09545_, _03655_);
  and (_09558_, _09557_, _09556_);
  or (_09559_, _09558_, _09555_);
  and (_09560_, _09559_, _04594_);
  and (_09561_, _09498_, _03773_);
  and (_09562_, _09561_, _09556_);
  or (_09563_, _09562_, _03653_);
  or (_09564_, _09563_, _09560_);
  nor (_09565_, _05959_, _09486_);
  or (_09566_, _09485_, _04608_);
  or (_09567_, _09566_, _09565_);
  and (_09568_, _09567_, _04606_);
  and (_09569_, _09568_, _09564_);
  nor (_09570_, _06457_, _09486_);
  or (_09571_, _09570_, _09485_);
  and (_09572_, _09571_, _03786_);
  or (_09573_, _09572_, _03809_);
  or (_09574_, _09573_, _09569_);
  or (_09575_, _09495_, _04260_);
  and (_09576_, _09575_, _03206_);
  and (_09577_, _09576_, _09574_);
  and (_09578_, _09492_, _03205_);
  or (_09579_, _09578_, _03816_);
  or (_09580_, _09579_, _09577_);
  and (_09581_, _05895_, _05386_);
  or (_09582_, _09485_, _03820_);
  or (_09583_, _09582_, _09581_);
  and (_09584_, _09583_, _43227_);
  and (_09585_, _09584_, _09580_);
  nor (_09586_, _43227_, _09484_);
  or (_09587_, _09586_, rst);
  or (_40754_, _09587_, _09585_);
  not (_09588_, \oc8051_golden_model_1.P3 [7]);
  nor (_09589_, _43227_, _09588_);
  or (_09590_, _09589_, rst);
  nor (_09591_, _05388_, _09588_);
  not (_09592_, _05388_);
  nor (_09593_, _09592_, _05289_);
  or (_09594_, _09593_, _09591_);
  or (_09595_, _09594_, _06889_);
  nor (_09596_, _06016_, _09588_);
  and (_09597_, _06038_, _06016_);
  or (_09598_, _09597_, _09596_);
  and (_09599_, _09598_, _03511_);
  and (_09600_, _06185_, _05388_);
  or (_09601_, _09600_, _09591_);
  or (_09602_, _09601_, _04515_);
  and (_09603_, _05388_, \oc8051_golden_model_1.ACC [7]);
  or (_09604_, _09603_, _09591_);
  and (_09605_, _09604_, _04499_);
  nor (_09606_, _04499_, _09588_);
  or (_09607_, _09606_, _03599_);
  or (_09608_, _09607_, _09605_);
  and (_09609_, _09608_, _03516_);
  and (_09610_, _09609_, _09602_);
  and (_09611_, _06042_, _06016_);
  or (_09612_, _09611_, _09596_);
  and (_09613_, _09612_, _03515_);
  or (_09614_, _09613_, _03597_);
  or (_09615_, _09614_, _09610_);
  or (_09616_, _09594_, _04524_);
  and (_09617_, _09616_, _09615_);
  or (_09618_, _09617_, _03603_);
  or (_09619_, _09604_, _03611_);
  and (_09620_, _09619_, _03512_);
  and (_09621_, _09620_, _09618_);
  or (_09622_, _09621_, _09599_);
  and (_09623_, _09622_, _03505_);
  and (_09624_, _06217_, _06016_);
  or (_09625_, _09624_, _09596_);
  and (_09626_, _09625_, _03504_);
  or (_09627_, _09626_, _09623_);
  and (_09628_, _09627_, _03501_);
  and (_09629_, _09305_, _06016_);
  or (_09630_, _09629_, _09596_);
  and (_09631_, _09630_, _03500_);
  or (_09632_, _09631_, _07441_);
  or (_09633_, _09632_, _09628_);
  and (_09634_, _09633_, _09595_);
  or (_09635_, _09634_, _05969_);
  and (_09636_, _06171_, _05388_);
  or (_09637_, _09591_, _05970_);
  or (_09638_, _09637_, _09636_);
  and (_09639_, _09638_, _03275_);
  and (_09640_, _09639_, _09635_);
  and (_09641_, _09330_, _05388_);
  or (_09642_, _09641_, _09591_);
  and (_09643_, _09642_, _03644_);
  or (_09644_, _09643_, _08861_);
  or (_09645_, _09644_, _09640_);
  and (_09646_, _05961_, _05388_);
  or (_09647_, _09591_, _04591_);
  or (_09648_, _09647_, _09646_);
  and (_09649_, _06247_, _05388_);
  or (_09650_, _09649_, _09591_);
  or (_09651_, _09650_, _04582_);
  and (_09652_, _09651_, _04589_);
  and (_09653_, _09652_, _09648_);
  and (_09654_, _09653_, _09645_);
  and (_09655_, _06458_, _05388_);
  or (_09656_, _09655_, _09591_);
  and (_09657_, _09656_, _03778_);
  or (_09658_, _09657_, _09654_);
  and (_09659_, _09658_, _04596_);
  or (_09660_, _09591_, _05397_);
  and (_09661_, _09650_, _03655_);
  and (_09662_, _09661_, _09660_);
  or (_09663_, _09662_, _09659_);
  and (_09664_, _09663_, _04594_);
  and (_09665_, _09604_, _03773_);
  and (_09666_, _09665_, _09660_);
  or (_09667_, _09666_, _03653_);
  or (_09668_, _09667_, _09664_);
  nor (_09669_, _05959_, _09592_);
  or (_09670_, _09591_, _04608_);
  or (_09671_, _09670_, _09669_);
  and (_09672_, _09671_, _04606_);
  and (_09673_, _09672_, _09668_);
  nor (_09674_, _06457_, _09592_);
  or (_09675_, _09674_, _09591_);
  and (_09676_, _09675_, _03786_);
  or (_09677_, _09676_, _03809_);
  or (_09678_, _09677_, _09673_);
  or (_09679_, _09601_, _04260_);
  and (_09680_, _09679_, _03206_);
  and (_09681_, _09680_, _09678_);
  and (_09682_, _09598_, _03205_);
  or (_09683_, _09682_, _03816_);
  or (_09684_, _09683_, _09681_);
  and (_09685_, _05895_, _05388_);
  or (_09686_, _09591_, _03820_);
  or (_09687_, _09686_, _09685_);
  and (_09688_, _09687_, _43227_);
  and (_09689_, _09688_, _09684_);
  or (_40756_, _09689_, _09590_);
  not (_09690_, _08814_);
  not (_09691_, _08477_);
  nor (_09692_, _08799_, _08478_);
  nor (_09693_, _09692_, _08771_);
  nand (_09694_, _09693_, _09691_);
  nor (_09695_, _08672_, _08459_);
  nand (_09696_, _03245_, _03134_);
  or (_09697_, _09696_, _09695_);
  or (_09698_, _09697_, _07946_);
  and (_09699_, _07875_, _07871_);
  and (_09700_, _09699_, _05906_);
  nor (_09701_, _07861_, _06061_);
  or (_09702_, _09701_, _07928_);
  or (_09703_, _09702_, _09700_);
  or (_09704_, _09703_, _07933_);
  nor (_09705_, _05368_, _07911_);
  and (_09706_, _06458_, _05368_);
  or (_09707_, _09706_, _09705_);
  and (_09708_, _09707_, _03778_);
  not (_09709_, _05368_);
  nor (_09710_, _06443_, _09709_);
  or (_09711_, _09710_, _09705_);
  and (_09712_, _09711_, _03644_);
  nor (_09713_, _09709_, _05289_);
  or (_09714_, _09713_, _09705_);
  or (_09715_, _09714_, _06889_);
  and (_09716_, _08285_, _08283_);
  nand (_09717_, _09716_, _08174_);
  nor (_09718_, _09717_, _06211_);
  and (_09719_, _08281_, _08278_);
  nor (_09720_, _09719_, _08276_);
  not (_09721_, _09720_);
  and (_09722_, _08573_, _08278_);
  not (_09723_, _09722_);
  nor (_09724_, _09723_, _08326_);
  nor (_09725_, _09724_, _09721_);
  or (_09726_, _09725_, _09718_);
  and (_09727_, _09726_, _03635_);
  not (_09728_, _03629_);
  not (_09729_, _03630_);
  not (_09730_, _05318_);
  and (_09731_, _05989_, \oc8051_golden_model_1.IP [2]);
  and (_09732_, _05983_, \oc8051_golden_model_1.ACC [2]);
  nor (_09733_, _09732_, _09731_);
  and (_09734_, _05976_, \oc8051_golden_model_1.SCON [2]);
  and (_09735_, _05979_, \oc8051_golden_model_1.IE [2]);
  nor (_09736_, _09735_, _09734_);
  and (_09737_, _06000_, \oc8051_golden_model_1.PSW [2]);
  and (_09738_, _05992_, \oc8051_golden_model_1.B [2]);
  nor (_09739_, _09738_, _09737_);
  and (_09740_, _09739_, _09736_);
  and (_09741_, _09740_, _09733_);
  and (_09742_, _05997_, \oc8051_golden_model_1.TCON [2]);
  and (_09743_, _05294_, \oc8051_golden_model_1.P0INREG [2]);
  nor (_09744_, _09743_, _09742_);
  and (_09745_, _06016_, \oc8051_golden_model_1.P3INREG [2]);
  not (_09746_, _09745_);
  and (_09747_, _06013_, \oc8051_golden_model_1.P1INREG [2]);
  and (_09748_, _06009_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_09749_, _09748_, _09747_);
  and (_09750_, _09749_, _09746_);
  and (_09751_, _09750_, _09744_);
  and (_09752_, _09751_, _09741_);
  and (_09753_, _09752_, _05746_);
  nor (_09754_, _09753_, _09730_);
  not (_09755_, _05314_);
  and (_09756_, _05997_, \oc8051_golden_model_1.TCON [1]);
  and (_09757_, _05992_, \oc8051_golden_model_1.B [1]);
  nor (_09758_, _09757_, _09756_);
  and (_09759_, _05989_, \oc8051_golden_model_1.IP [1]);
  not (_09760_, _09759_);
  and (_09761_, _06000_, \oc8051_golden_model_1.PSW [1]);
  and (_09762_, _05983_, \oc8051_golden_model_1.ACC [1]);
  nor (_09763_, _09762_, _09761_);
  and (_09764_, _09763_, _09760_);
  and (_09765_, _09764_, _09758_);
  and (_09766_, _05976_, \oc8051_golden_model_1.SCON [1]);
  and (_09767_, _05979_, \oc8051_golden_model_1.IE [1]);
  nor (_09768_, _09767_, _09766_);
  and (_09769_, _05294_, \oc8051_golden_model_1.P0INREG [1]);
  and (_09770_, _06009_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_09771_, _09770_, _09769_);
  and (_09772_, _06013_, \oc8051_golden_model_1.P1INREG [1]);
  and (_09773_, _06016_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_09774_, _09773_, _09772_);
  and (_09775_, _09774_, _09771_);
  and (_09776_, _09775_, _09768_);
  and (_09777_, _09776_, _09765_);
  and (_09778_, _09777_, _05651_);
  nor (_09779_, _09778_, _09755_);
  nor (_09780_, _09779_, _09754_);
  and (_09781_, _05301_, _03899_);
  not (_09782_, _09781_);
  and (_09783_, _05976_, \oc8051_golden_model_1.SCON [4]);
  and (_09784_, _05979_, \oc8051_golden_model_1.IE [4]);
  nor (_09785_, _09784_, _09783_);
  and (_09786_, _05997_, \oc8051_golden_model_1.TCON [4]);
  and (_09787_, _06016_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_09788_, _09787_, _09786_);
  and (_09789_, _09788_, _09785_);
  and (_09790_, _06000_, \oc8051_golden_model_1.PSW [4]);
  and (_09791_, _05992_, \oc8051_golden_model_1.B [4]);
  nor (_09792_, _09791_, _09790_);
  and (_09793_, _05989_, \oc8051_golden_model_1.IP [4]);
  and (_09794_, _05983_, \oc8051_golden_model_1.ACC [4]);
  nor (_09795_, _09794_, _09793_);
  and (_09796_, _09795_, _09792_);
  and (_09797_, _06013_, \oc8051_golden_model_1.P1INREG [4]);
  and (_09798_, _06009_, \oc8051_golden_model_1.P2INREG [4]);
  and (_09799_, _05294_, \oc8051_golden_model_1.P0INREG [4]);
  or (_09800_, _09799_, _09798_);
  nor (_09801_, _09800_, _09797_);
  and (_09802_, _09801_, _09796_);
  and (_09803_, _09802_, _09789_);
  and (_09804_, _09803_, _05841_);
  nor (_09805_, _09804_, _09782_);
  nor (_09806_, _06023_, _06041_);
  nor (_09807_, _09806_, _09805_);
  and (_09808_, _09807_, _09780_);
  not (_09809_, _05332_);
  and (_09810_, _05997_, \oc8051_golden_model_1.TCON [0]);
  and (_09811_, _05992_, \oc8051_golden_model_1.B [0]);
  nor (_09812_, _09811_, _09810_);
  and (_09813_, _06000_, \oc8051_golden_model_1.PSW [0]);
  not (_09814_, _09813_);
  and (_09815_, _05989_, \oc8051_golden_model_1.IP [0]);
  and (_09816_, _05983_, \oc8051_golden_model_1.ACC [0]);
  nor (_09817_, _09816_, _09815_);
  and (_09818_, _09817_, _09814_);
  and (_09819_, _09818_, _09812_);
  and (_09820_, _05976_, \oc8051_golden_model_1.SCON [0]);
  and (_09821_, _05979_, \oc8051_golden_model_1.IE [0]);
  nor (_09822_, _09821_, _09820_);
  and (_09823_, _05294_, \oc8051_golden_model_1.P0INREG [0]);
  and (_09824_, _06009_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_09825_, _09824_, _09823_);
  and (_09826_, _06013_, \oc8051_golden_model_1.P1INREG [0]);
  and (_09827_, _06016_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_09828_, _09827_, _09826_);
  and (_09829_, _09828_, _09825_);
  and (_09830_, _09829_, _09822_);
  and (_09831_, _09830_, _09819_);
  and (_09832_, _09831_, _05700_);
  nor (_09833_, _09832_, _09809_);
  and (_09834_, _05317_, _03899_);
  not (_09835_, _09834_);
  and (_09836_, _05997_, \oc8051_golden_model_1.TCON [6]);
  and (_09837_, _05992_, \oc8051_golden_model_1.B [6]);
  nor (_09838_, _09837_, _09836_);
  and (_09839_, _06000_, \oc8051_golden_model_1.PSW [6]);
  not (_09840_, _09839_);
  and (_09841_, _05989_, \oc8051_golden_model_1.IP [6]);
  and (_09842_, _05983_, \oc8051_golden_model_1.ACC [6]);
  nor (_09843_, _09842_, _09841_);
  and (_09844_, _09843_, _09840_);
  and (_09845_, _09844_, _09838_);
  and (_09846_, _05976_, \oc8051_golden_model_1.SCON [6]);
  and (_09847_, _05979_, \oc8051_golden_model_1.IE [6]);
  nor (_09848_, _09847_, _09846_);
  and (_09849_, _05294_, \oc8051_golden_model_1.P0INREG [6]);
  and (_09850_, _06013_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_09851_, _09850_, _09849_);
  and (_09852_, _06009_, \oc8051_golden_model_1.P2INREG [6]);
  and (_09853_, _06016_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_09854_, _09853_, _09852_);
  and (_09855_, _09854_, _09851_);
  and (_09856_, _09855_, _09848_);
  and (_09857_, _09856_, _09845_);
  and (_09858_, _09857_, _05443_);
  nor (_09859_, _09858_, _09835_);
  nor (_09860_, _09859_, _09833_);
  not (_09861_, _05296_);
  and (_09862_, _05997_, \oc8051_golden_model_1.TCON [3]);
  and (_09863_, _05983_, \oc8051_golden_model_1.ACC [3]);
  nor (_09864_, _09863_, _09862_);
  and (_09865_, _05989_, \oc8051_golden_model_1.IP [3]);
  not (_09866_, _09865_);
  and (_09867_, _06000_, \oc8051_golden_model_1.PSW [3]);
  and (_09868_, _05992_, \oc8051_golden_model_1.B [3]);
  nor (_09869_, _09868_, _09867_);
  and (_09870_, _09869_, _09866_);
  and (_09871_, _09870_, _09864_);
  and (_09872_, _05976_, \oc8051_golden_model_1.SCON [3]);
  and (_09873_, _05979_, \oc8051_golden_model_1.IE [3]);
  nor (_09874_, _09873_, _09872_);
  and (_09875_, _05294_, \oc8051_golden_model_1.P0INREG [3]);
  and (_09876_, _06009_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_09877_, _09876_, _09875_);
  and (_09878_, _06013_, \oc8051_golden_model_1.P1INREG [3]);
  and (_09879_, _06016_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_09880_, _09879_, _09878_);
  and (_09881_, _09880_, _09877_);
  and (_09882_, _09881_, _09874_);
  and (_09883_, _09882_, _09871_);
  and (_09884_, _09883_, _05602_);
  nor (_09885_, _09884_, _09861_);
  and (_09886_, _05313_, _03899_);
  not (_09887_, _09886_);
  and (_09888_, _05989_, \oc8051_golden_model_1.IP [5]);
  and (_09889_, _05983_, \oc8051_golden_model_1.ACC [5]);
  nor (_09890_, _09889_, _09888_);
  and (_09891_, _05976_, \oc8051_golden_model_1.SCON [5]);
  and (_09892_, _05979_, \oc8051_golden_model_1.IE [5]);
  nor (_09893_, _09892_, _09891_);
  and (_09894_, _06000_, \oc8051_golden_model_1.PSW [5]);
  and (_09895_, _05992_, \oc8051_golden_model_1.B [5]);
  nor (_09896_, _09895_, _09894_);
  and (_09897_, _09896_, _09893_);
  and (_09898_, _09897_, _09890_);
  and (_09899_, _05997_, \oc8051_golden_model_1.TCON [5]);
  and (_09900_, _06016_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_09901_, _09900_, _09899_);
  and (_09902_, _06009_, \oc8051_golden_model_1.P2INREG [5]);
  not (_09903_, _09902_);
  and (_09904_, _05294_, \oc8051_golden_model_1.P0INREG [5]);
  and (_09905_, _06013_, \oc8051_golden_model_1.P1INREG [5]);
  nor (_09906_, _09905_, _09904_);
  and (_09907_, _09906_, _09903_);
  and (_09908_, _09907_, _09901_);
  and (_09909_, _09908_, _09898_);
  and (_09910_, _09909_, _05553_);
  nor (_09911_, _09910_, _09887_);
  nor (_09912_, _09911_, _09885_);
  and (_09913_, _09912_, _09860_);
  and (_09914_, _09913_, _09808_);
  nor (_09915_, _09914_, _09729_);
  not (_09916_, _03676_);
  nor (_09917_, _08191_, \oc8051_golden_model_1.ACC [3]);
  and (_09918_, _08191_, \oc8051_golden_model_1.ACC [3]);
  nor (_09919_, _09918_, _09917_);
  and (_09920_, _09919_, _08742_);
  not (_09921_, _08746_);
  and (_09922_, _08238_, \oc8051_golden_model_1.ACC [0]);
  nor (_09923_, _09922_, _09921_);
  or (_09924_, _09923_, _08744_);
  and (_09925_, _09924_, _09920_);
  and (_09926_, _09919_, _08741_);
  or (_09927_, _09926_, _09917_);
  or (_09928_, _09927_, _09925_);
  and (_09929_, _08733_, _08737_);
  not (_09930_, _08725_);
  and (_09931_, _08729_, _09930_);
  and (_09932_, _09931_, _09929_);
  and (_09933_, _09932_, _09928_);
  nor (_09934_, _08736_, _08731_);
  nor (_09935_, _09934_, _08732_);
  and (_09936_, _09931_, _09935_);
  nor (_09937_, _06211_, \oc8051_golden_model_1.ACC [7]);
  and (_09938_, _08728_, _09930_);
  or (_09939_, _09938_, _09937_);
  or (_09940_, _09939_, _09936_);
  or (_09941_, _09940_, _09933_);
  nor (_09942_, _08238_, \oc8051_golden_model_1.ACC [0]);
  nor (_09943_, _09922_, _09942_);
  and (_09944_, _09943_, _08746_);
  and (_09945_, _09944_, _09920_);
  and (_09946_, _09932_, _09945_);
  nor (_09947_, _09946_, _04046_);
  and (_09948_, _09947_, _09941_);
  and (_09949_, _06185_, _05368_);
  nor (_09950_, _09949_, _09705_);
  nand (_09951_, _09950_, _03599_);
  not (_09952_, _08063_);
  and (_09953_, _05368_, \oc8051_golden_model_1.ACC [7]);
  or (_09954_, _09953_, _09705_);
  and (_09955_, _09954_, _04499_);
  nor (_09956_, _04499_, _07911_);
  or (_09957_, _09956_, _03599_);
  or (_09958_, _09957_, _09955_);
  and (_09959_, _09958_, _09952_);
  and (_09960_, _09959_, _09951_);
  nor (_09961_, _08073_, \oc8051_golden_model_1.PSW [7]);
  not (_09962_, _09961_);
  nor (_09963_, _09962_, _08083_);
  nor (_09964_, _09963_, _09952_);
  nor (_09965_, _03284_, _03255_);
  not (_09966_, _09965_);
  nand (_09967_, _09966_, _03604_);
  or (_09968_, _09967_, _09964_);
  or (_09969_, _09968_, _09960_);
  nor (_09970_, _06000_, _07911_);
  and (_09971_, _06042_, _06000_);
  or (_09972_, _09971_, _09970_);
  or (_09973_, _09972_, _03516_);
  or (_09974_, _09714_, _04524_);
  and (_09975_, _09974_, _09973_);
  and (_09976_, _09975_, _09969_);
  or (_09977_, _09976_, _03603_);
  or (_09978_, _09954_, _03611_);
  nor (_09979_, _03284_, _03259_);
  nor (_09980_, _09979_, _03511_);
  and (_09981_, _09980_, _09978_);
  and (_09982_, _09981_, _09977_);
  and (_09983_, _06038_, _06000_);
  nor (_09984_, _09983_, _09970_);
  nor (_09985_, _09984_, _03512_);
  or (_09986_, _09985_, _09982_);
  nor (_09987_, _05964_, _03252_);
  nor (_09988_, _09987_, _03667_);
  and (_09989_, _09988_, _09986_);
  and (_09990_, _04944_, _03558_);
  and (_09991_, _05130_, _03899_);
  nor (_09992_, _09991_, _09990_);
  nor (_09993_, _04944_, _03558_);
  nor (_09994_, _05130_, _03899_);
  nor (_09995_, _09994_, _09993_);
  and (_09996_, _09995_, _09992_);
  and (_09997_, _04699_, _04435_);
  and (_09998_, _05898_, _04434_);
  and (_09999_, _04491_, _04042_);
  or (_10000_, _09999_, _09997_);
  nor (_10001_, _10000_, _09998_);
  or (_10002_, _10001_, _09997_);
  and (_10003_, _10002_, _09996_);
  not (_10004_, _09991_);
  nor (_10005_, _09993_, _10004_);
  or (_10006_, _10005_, _09990_);
  or (_10007_, _10006_, _10003_);
  and (_10008_, _05289_, _03463_);
  not (_10009_, _10008_);
  and (_10010_, _10009_, _05290_);
  and (_10011_, _05442_, _03556_);
  nor (_10012_, _05442_, _03556_);
  or (_10013_, _10012_, _10011_);
  and (_10014_, _10013_, _10010_);
  and (_10015_, _05552_, _05334_);
  nor (_10016_, _05552_, _05334_);
  nor (_10017_, _10016_, _10015_);
  and (_10018_, _05840_, _04308_);
  nor (_10019_, _05840_, _04308_);
  or (_10020_, _10019_, _10018_);
  and (_10021_, _10020_, _10017_);
  and (_10022_, _10021_, _10014_);
  and (_10023_, _10022_, _10007_);
  and (_10024_, _05840_, _05327_);
  and (_10025_, _10017_, _10024_);
  or (_10026_, _10025_, _10015_);
  and (_10027_, _10026_, _10014_);
  and (_10028_, _05442_, _05056_);
  and (_10029_, _10028_, _05290_);
  or (_10030_, _10029_, _10008_);
  or (_10031_, _10030_, _10027_);
  or (_10032_, _10031_, _10023_);
  and (_10033_, _04510_, _04192_);
  not (_10034_, _10033_);
  and (_10035_, _10001_, _09996_);
  and (_10036_, _10035_, _10034_);
  and (_10037_, _10036_, _10022_);
  nor (_10038_, _10037_, _09988_);
  and (_10039_, _10038_, _10032_);
  or (_10040_, _10039_, _09989_);
  and (_10041_, _04197_, _03503_);
  not (_10042_, _10041_);
  and (_10043_, _10042_, _10040_);
  and (_10044_, _06577_, _04435_);
  or (_10045_, _06577_, _04435_);
  and (_10046_, _06836_, _04042_);
  nor (_10047_, _10046_, _10044_);
  and (_10048_, _10047_, _10045_);
  or (_10049_, _10048_, _10044_);
  or (_10050_, _06838_, _03494_);
  or (_10051_, _06668_, _03558_);
  and (_10052_, _10051_, _10050_);
  and (_10053_, _06714_, _03899_);
  and (_10054_, _06839_, _03898_);
  nor (_10055_, _10054_, _10053_);
  and (_10056_, _10055_, _10052_);
  and (_10057_, _10056_, _10049_);
  nand (_10058_, _10052_, _10053_);
  nand (_10059_, _10058_, _10050_);
  or (_10060_, _10059_, _10057_);
  and (_10061_, _06806_, _05327_);
  and (_10062_, _06761_, _05334_);
  not (_10063_, _10062_);
  or (_10064_, _06761_, _05334_);
  nand (_10065_, _10064_, _10063_);
  nor (_10066_, _10065_, _10061_);
  and (_10067_, _06843_, _04308_);
  not (_10068_, _10067_);
  nand (_10069_, _06531_, _03556_);
  nor (_10070_, _06531_, _03556_);
  nor (_10071_, _06171_, _04559_);
  or (_10072_, _10071_, _06228_);
  nor (_10073_, _10072_, _10070_);
  and (_10074_, _10073_, _10069_);
  and (_10075_, _10074_, _10068_);
  and (_10076_, _10075_, _10066_);
  and (_10077_, _10076_, _10060_);
  or (_10078_, _10061_, _10062_);
  and (_10079_, _10074_, _10078_);
  and (_10080_, _10079_, _10064_);
  not (_10081_, _06228_);
  and (_10082_, _10070_, _10081_);
  or (_10083_, _10082_, _10071_);
  or (_10084_, _10083_, _10080_);
  or (_10085_, _10084_, _10077_);
  and (_10086_, _06622_, _04192_);
  nand (_10087_, _10056_, _10048_);
  nor (_10088_, _10087_, _10086_);
  and (_10089_, _10088_, _10076_);
  nor (_10090_, _10089_, _10042_);
  and (_10091_, _10090_, _10085_);
  or (_10092_, _10091_, _10043_);
  and (_10093_, _10092_, _04046_);
  or (_10094_, _10093_, _09948_);
  and (_10095_, _10094_, _09916_);
  nor (_10096_, _03284_, _03252_);
  nor (_10097_, _08781_, _08782_);
  nor (_10098_, _10097_, _08785_);
  nor (_10099_, _04434_, \oc8051_golden_model_1.ACC [1]);
  and (_10100_, _04434_, \oc8051_golden_model_1.ACC [1]);
  and (_10101_, _04042_, \oc8051_golden_model_1.ACC [0]);
  nor (_10102_, _10101_, _10100_);
  or (_10103_, _10102_, _10099_);
  and (_10104_, _10103_, _10098_);
  nand (_10105_, _03494_, \oc8051_golden_model_1.ACC [3]);
  nor (_10106_, _03494_, \oc8051_golden_model_1.ACC [3]);
  nor (_10107_, _03898_, \oc8051_golden_model_1.ACC [2]);
  or (_10108_, _10107_, _10106_);
  and (_10109_, _10108_, _10105_);
  or (_10110_, _10109_, _10104_);
  or (_10111_, _08776_, _08777_);
  not (_10112_, _10111_);
  nor (_10113_, _10112_, _08780_);
  nor (_10114_, _08775_, _08479_);
  and (_10115_, _10114_, _10113_);
  and (_10116_, _10115_, _10110_);
  nand (_10117_, _03853_, \oc8051_golden_model_1.ACC [5]);
  nor (_10118_, _03853_, \oc8051_golden_model_1.ACC [5]);
  nor (_10119_, _04308_, \oc8051_golden_model_1.ACC [4]);
  or (_10120_, _10119_, _10118_);
  and (_10121_, _10120_, _10117_);
  and (_10122_, _10121_, _10114_);
  and (_10123_, _03463_, _06061_);
  or (_10124_, _03556_, \oc8051_golden_model_1.ACC [6]);
  nor (_10125_, _10124_, _08479_);
  or (_10126_, _10125_, _10123_);
  or (_10127_, _10126_, _10122_);
  or (_10128_, _10127_, _10116_);
  and (_10129_, _04042_, _03397_);
  nor (_10130_, _10129_, _08787_);
  nor (_10131_, _10130_, _08383_);
  and (_10132_, _10131_, _10098_);
  and (_10133_, _10132_, _10115_);
  nor (_10134_, _10133_, _09916_);
  and (_10135_, _10134_, _10128_);
  or (_10136_, _10135_, _10096_);
  or (_10137_, _10136_, _10095_);
  nand (_10138_, _10096_, \oc8051_golden_model_1.PSW [7]);
  and (_10139_, _10138_, _03505_);
  and (_10140_, _10139_, _10137_);
  or (_10141_, _09970_, _06216_);
  and (_10142_, _09972_, _03504_);
  and (_10143_, _10142_, _10141_);
  nor (_10144_, _10143_, _10140_);
  nor (_10145_, _10144_, _03621_);
  and (_10146_, _05294_, \oc8051_golden_model_1.P0 [2]);
  and (_10147_, _06016_, \oc8051_golden_model_1.P3 [2]);
  nor (_10148_, _10147_, _10146_);
  not (_10149_, _09742_);
  and (_10150_, _06013_, \oc8051_golden_model_1.P1 [2]);
  and (_10151_, _06009_, \oc8051_golden_model_1.P2 [2]);
  nor (_10152_, _10151_, _10150_);
  and (_10153_, _10152_, _10149_);
  and (_10154_, _10153_, _10148_);
  and (_10155_, _10154_, _09741_);
  and (_10156_, _10155_, _05746_);
  nor (_10157_, _10156_, _09730_);
  and (_10158_, _06009_, \oc8051_golden_model_1.P2 [1]);
  and (_10159_, _06016_, \oc8051_golden_model_1.P3 [1]);
  nor (_10160_, _10159_, _10158_);
  and (_10161_, _05294_, \oc8051_golden_model_1.P0 [1]);
  and (_10162_, _06013_, \oc8051_golden_model_1.P1 [1]);
  nor (_10163_, _10162_, _10161_);
  and (_10164_, _10163_, _10160_);
  and (_10165_, _10164_, _09768_);
  and (_10166_, _10165_, _09765_);
  and (_10167_, _10166_, _05651_);
  nor (_10168_, _10167_, _09755_);
  nor (_10169_, _10168_, _10157_);
  and (_10170_, _05294_, \oc8051_golden_model_1.P0 [4]);
  and (_10171_, _06013_, \oc8051_golden_model_1.P1 [4]);
  nor (_10172_, _10171_, _10170_);
  and (_10173_, _06016_, \oc8051_golden_model_1.P3 [4]);
  and (_10174_, _06009_, \oc8051_golden_model_1.P2 [4]);
  or (_10175_, _10174_, _10173_);
  nor (_10176_, _10175_, _09786_);
  and (_10177_, _10176_, _09796_);
  and (_10178_, _10177_, _09785_);
  and (_10179_, _10178_, _10172_);
  and (_10180_, _10179_, _05841_);
  nor (_10181_, _09782_, _10180_);
  nor (_10182_, _10181_, _06215_);
  and (_10183_, _10182_, _10169_);
  and (_10184_, _06009_, \oc8051_golden_model_1.P2 [0]);
  and (_10185_, _06016_, \oc8051_golden_model_1.P3 [0]);
  nor (_10186_, _10185_, _10184_);
  and (_10187_, _05294_, \oc8051_golden_model_1.P0 [0]);
  and (_10188_, _06013_, \oc8051_golden_model_1.P1 [0]);
  nor (_10189_, _10188_, _10187_);
  and (_10190_, _10189_, _10186_);
  and (_10191_, _10190_, _09822_);
  and (_10192_, _10191_, _09819_);
  and (_10193_, _10192_, _05700_);
  nor (_10194_, _10193_, _09809_);
  and (_10195_, _06009_, \oc8051_golden_model_1.P2 [6]);
  and (_10196_, _06016_, \oc8051_golden_model_1.P3 [6]);
  nor (_10197_, _10196_, _10195_);
  and (_10198_, _05294_, \oc8051_golden_model_1.P0 [6]);
  and (_10199_, _06013_, \oc8051_golden_model_1.P1 [6]);
  nor (_10200_, _10199_, _10198_);
  and (_10201_, _10200_, _10197_);
  and (_10202_, _10201_, _09848_);
  and (_10203_, _10202_, _09845_);
  and (_10204_, _10203_, _05443_);
  nor (_10205_, _09835_, _10204_);
  nor (_10206_, _10205_, _10194_);
  and (_10207_, _06009_, \oc8051_golden_model_1.P2 [3]);
  and (_10208_, _06016_, \oc8051_golden_model_1.P3 [3]);
  nor (_10209_, _10208_, _10207_);
  and (_10210_, _05294_, \oc8051_golden_model_1.P0 [3]);
  and (_10211_, _06013_, \oc8051_golden_model_1.P1 [3]);
  nor (_10212_, _10211_, _10210_);
  and (_10213_, _10212_, _10209_);
  and (_10214_, _10213_, _09874_);
  and (_10215_, _10214_, _09871_);
  and (_10216_, _10215_, _05602_);
  nor (_10217_, _10216_, _09861_);
  and (_10218_, _05294_, \oc8051_golden_model_1.P0 [5]);
  and (_10219_, _06016_, \oc8051_golden_model_1.P3 [5]);
  nor (_10220_, _10219_, _10218_);
  not (_10221_, _09899_);
  and (_10222_, _06013_, \oc8051_golden_model_1.P1 [5]);
  and (_10223_, _06009_, \oc8051_golden_model_1.P2 [5]);
  nor (_10224_, _10223_, _10222_);
  and (_10225_, _10224_, _10221_);
  and (_10226_, _10225_, _10220_);
  and (_10227_, _10226_, _09898_);
  and (_10228_, _10227_, _05553_);
  nor (_10229_, _09887_, _10228_);
  nor (_10230_, _10229_, _10217_);
  and (_10231_, _10230_, _10206_);
  and (_10232_, _10231_, _10183_);
  and (_10233_, _03621_, \oc8051_golden_model_1.PSW [7]);
  and (_10234_, _10233_, _10232_);
  or (_10235_, _10234_, _10145_);
  nor (_10236_, _06919_, _03630_);
  and (_10237_, _10236_, _10235_);
  or (_10238_, _10237_, _09915_);
  and (_10239_, _10238_, _09728_);
  nor (_10240_, _08454_, _03277_);
  nor (_10241_, _10240_, _08034_);
  nor (_10242_, _05080_, _03277_);
  not (_10243_, _10242_);
  and (_10244_, _10243_, _10241_);
  not (_10245_, _10244_);
  or (_10246_, _10232_, \oc8051_golden_model_1.PSW [7]);
  and (_10247_, _10246_, _03629_);
  or (_10248_, _10247_, _10245_);
  or (_10249_, _10248_, _10239_);
  and (_10250_, _03570_, _03276_);
  not (_10251_, _10250_);
  and (_10252_, _07868_, _07864_);
  nor (_10253_, _10252_, _07862_);
  not (_10254_, _10253_);
  and (_10255_, _07870_, _07864_);
  not (_10256_, _10255_);
  nor (_10257_, _10256_, _08149_);
  nor (_10258_, _10257_, _10254_);
  or (_10259_, _10258_, _09700_);
  or (_10260_, _10259_, _10244_);
  and (_10261_, _10260_, _10251_);
  and (_10262_, _10261_, _10249_);
  and (_10263_, _10259_, _10250_);
  or (_10264_, _10263_, _08032_);
  or (_10265_, _10264_, _10262_);
  and (_10266_, _07973_, _07967_);
  nor (_10267_, _10266_, _07965_);
  not (_10268_, _10267_);
  and (_10269_, _08543_, _07967_);
  not (_10270_, _10269_);
  nor (_10271_, _10270_, _08026_);
  nor (_10272_, _10271_, _10268_);
  and (_10273_, _07970_, _06531_);
  and (_10274_, _10273_, _06171_);
  or (_10275_, _08128_, _10274_);
  or (_10276_, _10275_, _10272_);
  and (_10277_, _10276_, _03640_);
  and (_10278_, _10277_, _10265_);
  or (_10279_, _10278_, _09727_);
  and (_10280_, _10279_, _08161_);
  and (_10281_, _08336_, _05378_);
  and (_10282_, _08348_, _08344_);
  nor (_10283_, _10282_, _08342_);
  not (_10284_, _10283_);
  and (_10285_, _08604_, _08344_);
  not (_10286_, _10285_);
  nor (_10287_, _10286_, _08409_);
  nor (_10288_, _10287_, _10284_);
  or (_10289_, _10288_, _10281_);
  and (_10290_, _10289_, _08160_);
  or (_10291_, _10290_, _07441_);
  or (_10292_, _10291_, _10280_);
  and (_10293_, _10292_, _09715_);
  or (_10294_, _10293_, _05969_);
  and (_10295_, _06171_, _05368_);
  or (_10296_, _09705_, _05970_);
  or (_10297_, _10296_, _10295_);
  and (_10298_, _10297_, _03275_);
  and (_10299_, _10298_, _10294_);
  or (_10300_, _10299_, _09712_);
  nor (_10301_, _07455_, _03562_);
  and (_10302_, _10301_, _10300_);
  nor (_10303_, _10232_, _07911_);
  and (_10304_, _10303_, _03562_);
  or (_10305_, _10304_, _03650_);
  or (_10306_, _10305_, _10302_);
  and (_10307_, _06247_, _05368_);
  or (_10308_, _10307_, _09705_);
  or (_10309_, _10308_, _04582_);
  and (_10310_, _10309_, _10306_);
  or (_10311_, _10310_, _03561_);
  nand (_10312_, _10232_, _07911_);
  or (_10313_, _10312_, _04181_);
  and (_10314_, _10313_, _10311_);
  or (_10315_, _10314_, _03649_);
  and (_10316_, _05961_, _05368_);
  or (_10317_, _10316_, _09705_);
  or (_10318_, _10317_, _04591_);
  and (_10319_, _10318_, _04589_);
  and (_10320_, _10319_, _10315_);
  or (_10321_, _10320_, _09708_);
  and (_10322_, _10321_, _04596_);
  or (_10323_, _09705_, _05397_);
  and (_10324_, _10308_, _03655_);
  and (_10325_, _10324_, _10323_);
  or (_10326_, _10325_, _10322_);
  and (_10327_, _10326_, _04594_);
  and (_10328_, _09954_, _03773_);
  and (_10329_, _10328_, _10323_);
  or (_10330_, _10329_, _03653_);
  or (_10331_, _10330_, _10327_);
  nor (_10332_, _05959_, _09709_);
  or (_10333_, _09705_, _04608_);
  or (_10334_, _10333_, _10332_);
  and (_10335_, _10334_, _04606_);
  and (_10336_, _10335_, _10331_);
  nor (_10337_, _06457_, _09709_);
  or (_10338_, _10337_, _09705_);
  and (_10339_, _10338_, _03786_);
  or (_10340_, _10339_, _08532_);
  or (_10341_, _10340_, _10336_);
  and (_10342_, _10341_, _09704_);
  or (_10343_, _10342_, _08539_);
  nor (_10344_, _07964_, _06061_);
  or (_10345_, _10344_, _08563_);
  or (_10346_, _08541_, _10274_);
  or (_10347_, _10346_, _10345_);
  and (_10348_, _10347_, _03783_);
  and (_10349_, _10348_, _10343_);
  nor (_10350_, _08275_, _06061_);
  or (_10351_, _10350_, _08594_);
  or (_10352_, _10351_, _09718_);
  and (_10353_, _10352_, _03782_);
  or (_10354_, _10353_, _10349_);
  or (_10355_, _10354_, _08569_);
  nor (_10356_, _08341_, _06061_);
  nor (_10357_, _10356_, _08625_);
  nor (_10358_, _10281_, _08602_);
  nand (_10359_, _10358_, _10357_);
  and (_10360_, _10359_, _08601_);
  and (_10361_, _10360_, _10355_);
  not (_10362_, _09696_);
  and (_10363_, _08600_, \oc8051_golden_model_1.ACC [7]);
  or (_10364_, _10363_, _10362_);
  or (_10365_, _10364_, _10361_);
  and (_10366_, _10365_, _09698_);
  or (_10367_, _10366_, _08679_);
  and (_10368_, _08712_, _07955_);
  not (_10369_, _08679_);
  nor (_10370_, _08683_, _07954_);
  nor (_10371_, _10370_, _07935_);
  or (_10372_, _10371_, _10369_);
  or (_10373_, _10372_, _10368_);
  and (_10374_, _10373_, _03525_);
  and (_10375_, _10374_, _10367_);
  not (_10376_, _08723_);
  not (_10377_, _08724_);
  and (_10378_, _08762_, _10377_);
  nor (_10379_, _10378_, _03525_);
  and (_10380_, _10379_, _10376_);
  or (_10381_, _10380_, _08720_);
  or (_10382_, _10381_, _10375_);
  and (_10383_, _10382_, _09694_);
  and (_10384_, _10383_, _04260_);
  nor (_10385_, _09950_, _04260_);
  or (_10386_, _10385_, _10384_);
  and (_10387_, _10386_, _09690_);
  and (_10388_, _08814_, \oc8051_golden_model_1.ACC [0]);
  or (_10389_, _10388_, _10387_);
  and (_10390_, _10389_, _03206_);
  nor (_10391_, _09984_, _03206_);
  or (_10392_, _10391_, _10390_);
  and (_10393_, _10392_, _03820_);
  and (_10394_, _05895_, _05368_);
  nor (_10395_, _10394_, _09705_);
  nor (_10396_, _10395_, _03820_);
  or (_10397_, _10396_, _10393_);
  or (_10398_, _10397_, _43231_);
  or (_10399_, _43227_, \oc8051_golden_model_1.PSW [7]);
  and (_10400_, _10399_, _41991_);
  and (_40757_, _10400_, _10398_);
  not (_10401_, \oc8051_golden_model_1.PCON [7]);
  nor (_10402_, _05323_, _10401_);
  not (_10403_, _05323_);
  nor (_10404_, _06457_, _10403_);
  nor (_10405_, _10404_, _10402_);
  nor (_10406_, _10405_, _04606_);
  and (_10407_, _06247_, _05323_);
  nor (_10408_, _10407_, _10402_);
  and (_10409_, _10408_, _03650_);
  nor (_10410_, _10403_, _05289_);
  nor (_10411_, _10410_, _10402_);
  and (_10412_, _10411_, _07441_);
  and (_10413_, _05323_, \oc8051_golden_model_1.ACC [7]);
  nor (_10414_, _10413_, _10402_);
  nor (_10415_, _10414_, _04500_);
  nor (_10416_, _04499_, _10401_);
  or (_10417_, _10416_, _10415_);
  and (_10418_, _10417_, _04515_);
  and (_10419_, _06185_, _05323_);
  nor (_10420_, _10419_, _10402_);
  nor (_10421_, _10420_, _04515_);
  or (_10422_, _10421_, _10418_);
  and (_10423_, _10422_, _04524_);
  nor (_10424_, _10411_, _04524_);
  nor (_10425_, _10424_, _10423_);
  nor (_10426_, _10425_, _03603_);
  nor (_10427_, _10414_, _03611_);
  nor (_10428_, _10427_, _07441_);
  not (_10429_, _10428_);
  nor (_10430_, _10429_, _10426_);
  nor (_10431_, _10430_, _10412_);
  nor (_10432_, _10431_, _05969_);
  and (_10433_, _06171_, _05323_);
  nor (_10434_, _10402_, _05970_);
  not (_10435_, _10434_);
  nor (_10436_, _10435_, _10433_);
  or (_10437_, _10436_, _03644_);
  nor (_10438_, _10437_, _10432_);
  nor (_10439_, _06443_, _10403_);
  nor (_10440_, _10439_, _10402_);
  nor (_10441_, _10440_, _03275_);
  or (_10442_, _10441_, _03650_);
  nor (_10443_, _10442_, _10438_);
  nor (_10444_, _10443_, _10409_);
  or (_10445_, _10444_, _03649_);
  and (_10446_, _05961_, _05323_);
  or (_10447_, _10446_, _10402_);
  or (_10448_, _10447_, _04591_);
  and (_10449_, _10448_, _04589_);
  and (_10450_, _10449_, _10445_);
  and (_10451_, _06458_, _05323_);
  nor (_10452_, _10451_, _10402_);
  nor (_10453_, _10452_, _04589_);
  nor (_10454_, _10453_, _10450_);
  nor (_10455_, _10454_, _03655_);
  nor (_10456_, _10402_, _05397_);
  not (_10457_, _10456_);
  nor (_10458_, _10408_, _04596_);
  and (_10459_, _10458_, _10457_);
  nor (_10460_, _10459_, _10455_);
  nor (_10461_, _10460_, _03773_);
  nor (_10462_, _10414_, _04594_);
  and (_10463_, _10462_, _10457_);
  or (_10464_, _10463_, _10461_);
  and (_10465_, _10464_, _04608_);
  nor (_10466_, _05959_, _10403_);
  nor (_10467_, _10466_, _10402_);
  nor (_10468_, _10467_, _04608_);
  or (_10469_, _10468_, _10465_);
  and (_10470_, _10469_, _04606_);
  nor (_10471_, _10470_, _10406_);
  nor (_10472_, _10471_, _03809_);
  nor (_10473_, _10420_, _04260_);
  or (_10474_, _10473_, _03816_);
  nor (_10475_, _10474_, _10472_);
  and (_10476_, _05895_, _05323_);
  or (_10477_, _10402_, _03820_);
  nor (_10478_, _10477_, _10476_);
  nor (_10479_, _10478_, _10475_);
  or (_10480_, _10479_, _43231_);
  or (_10481_, _43227_, \oc8051_golden_model_1.PCON [7]);
  and (_10482_, _10481_, _41991_);
  and (_40758_, _10482_, _10480_);
  not (_10483_, \oc8051_golden_model_1.SBUF [7]);
  nor (_10484_, _05330_, _10483_);
  not (_10485_, _05330_);
  nor (_10486_, _06457_, _10485_);
  nor (_10487_, _10486_, _10484_);
  nor (_10488_, _10487_, _04606_);
  and (_10489_, _06247_, _05330_);
  nor (_10490_, _10489_, _10484_);
  and (_10491_, _10490_, _03650_);
  nor (_10492_, _10485_, _05289_);
  nor (_10493_, _10492_, _10484_);
  and (_10494_, _10493_, _07441_);
  and (_10495_, _05330_, \oc8051_golden_model_1.ACC [7]);
  nor (_10496_, _10495_, _10484_);
  nor (_10497_, _10496_, _03611_);
  nor (_10498_, _10496_, _04500_);
  nor (_10499_, _04499_, _10483_);
  or (_10500_, _10499_, _10498_);
  and (_10501_, _10500_, _04515_);
  and (_10502_, _06185_, _05330_);
  nor (_10503_, _10502_, _10484_);
  nor (_10504_, _10503_, _04515_);
  or (_10505_, _10504_, _10501_);
  and (_10506_, _10505_, _04524_);
  nor (_10507_, _10493_, _04524_);
  nor (_10508_, _10507_, _10506_);
  nor (_10509_, _10508_, _03603_);
  or (_10510_, _10509_, _07441_);
  nor (_10511_, _10510_, _10497_);
  nor (_10512_, _10511_, _10494_);
  nor (_10513_, _10512_, _05969_);
  and (_10514_, _06171_, _05330_);
  nor (_10515_, _10484_, _05970_);
  not (_10516_, _10515_);
  nor (_10517_, _10516_, _10514_);
  or (_10518_, _10517_, _03644_);
  nor (_10519_, _10518_, _10513_);
  nor (_10520_, _06443_, _10485_);
  nor (_10521_, _10520_, _10484_);
  nor (_10522_, _10521_, _03275_);
  or (_10523_, _10522_, _03650_);
  nor (_10524_, _10523_, _10519_);
  nor (_10525_, _10524_, _10491_);
  or (_10526_, _10525_, _03649_);
  and (_10527_, _05961_, _05330_);
  or (_10528_, _10527_, _10484_);
  or (_10529_, _10528_, _04591_);
  and (_10530_, _10529_, _04589_);
  and (_10531_, _10530_, _10526_);
  and (_10532_, _06458_, _05330_);
  nor (_10533_, _10532_, _10484_);
  nor (_10534_, _10533_, _04589_);
  nor (_10535_, _10534_, _10531_);
  nor (_10536_, _10535_, _03655_);
  nor (_10537_, _10484_, _05397_);
  not (_10538_, _10537_);
  nor (_10539_, _10490_, _04596_);
  and (_10540_, _10539_, _10538_);
  nor (_10541_, _10540_, _10536_);
  nor (_10542_, _10541_, _03773_);
  nor (_10543_, _10496_, _04594_);
  and (_10544_, _10543_, _10538_);
  or (_10545_, _10544_, _10542_);
  and (_10546_, _10545_, _04608_);
  nor (_10547_, _05959_, _10485_);
  nor (_10548_, _10547_, _10484_);
  nor (_10549_, _10548_, _04608_);
  or (_10550_, _10549_, _10546_);
  and (_10551_, _10550_, _04606_);
  nor (_10552_, _10551_, _10488_);
  nor (_10553_, _10552_, _03809_);
  nor (_10554_, _10503_, _04260_);
  or (_10555_, _10554_, _03816_);
  nor (_10556_, _10555_, _10553_);
  and (_10557_, _05895_, _05330_);
  or (_10558_, _10484_, _03820_);
  nor (_10559_, _10558_, _10557_);
  nor (_10560_, _10559_, _10556_);
  or (_10561_, _10560_, _43231_);
  or (_10562_, _43227_, \oc8051_golden_model_1.SBUF [7]);
  and (_10563_, _10562_, _41991_);
  and (_40759_, _10563_, _10561_);
  not (_10564_, \oc8051_golden_model_1.SCON [7]);
  nor (_10565_, _05345_, _10564_);
  not (_10566_, _05345_);
  nor (_10567_, _10566_, _05289_);
  nor (_10568_, _10567_, _10565_);
  and (_10569_, _10568_, _07441_);
  nor (_10570_, _05976_, _10564_);
  and (_10571_, _06038_, _05976_);
  nor (_10572_, _10571_, _10570_);
  nor (_10573_, _10572_, _03512_);
  and (_10574_, _05345_, \oc8051_golden_model_1.ACC [7]);
  nor (_10575_, _10574_, _10565_);
  nor (_10576_, _10575_, _04500_);
  nor (_10577_, _04499_, _10564_);
  or (_10578_, _10577_, _10576_);
  and (_10579_, _10578_, _04515_);
  and (_10580_, _06185_, _05345_);
  nor (_10581_, _10580_, _10565_);
  nor (_10582_, _10581_, _04515_);
  or (_10583_, _10582_, _10579_);
  and (_10584_, _10583_, _03516_);
  and (_10585_, _06042_, _05976_);
  nor (_10586_, _10585_, _10570_);
  nor (_10587_, _10586_, _03516_);
  or (_10588_, _10587_, _03597_);
  or (_10589_, _10588_, _10584_);
  nand (_10590_, _10568_, _03597_);
  and (_10591_, _10590_, _10589_);
  and (_10592_, _10591_, _03611_);
  nor (_10593_, _10575_, _03611_);
  or (_10594_, _10593_, _10592_);
  and (_10595_, _10594_, _03512_);
  nor (_10596_, _10595_, _10573_);
  nor (_10597_, _10596_, _03504_);
  nor (_10598_, _10570_, _06216_);
  or (_10599_, _10586_, _03505_);
  nor (_10600_, _10599_, _10598_);
  nor (_10601_, _10600_, _10597_);
  nor (_10602_, _10601_, _03500_);
  not (_10603_, _05976_);
  nor (_10604_, _06026_, _10603_);
  nor (_10605_, _10604_, _10570_);
  nor (_10606_, _10605_, _03501_);
  nor (_10607_, _10606_, _07441_);
  not (_10608_, _10607_);
  nor (_10609_, _10608_, _10602_);
  nor (_10610_, _10609_, _10569_);
  nor (_10611_, _10610_, _05969_);
  and (_10612_, _06171_, _05345_);
  nor (_10613_, _10565_, _05970_);
  not (_10614_, _10613_);
  nor (_10615_, _10614_, _10612_);
  nor (_10616_, _10615_, _03644_);
  not (_10617_, _10616_);
  nor (_10618_, _10617_, _10611_);
  nor (_10619_, _06443_, _10566_);
  nor (_10620_, _10619_, _10565_);
  nor (_10621_, _10620_, _03275_);
  or (_10622_, _10621_, _08861_);
  or (_10623_, _10622_, _10618_);
  and (_10624_, _05961_, _05345_);
  or (_10625_, _10565_, _04591_);
  or (_10626_, _10625_, _10624_);
  and (_10627_, _06247_, _05345_);
  nor (_10628_, _10627_, _10565_);
  and (_10629_, _10628_, _03650_);
  nor (_10630_, _10629_, _03778_);
  and (_10631_, _10630_, _10626_);
  and (_10632_, _10631_, _10623_);
  and (_10633_, _06458_, _05345_);
  nor (_10634_, _10633_, _10565_);
  nor (_10635_, _10634_, _04589_);
  nor (_10636_, _10635_, _10632_);
  nor (_10637_, _10636_, _03655_);
  nor (_10638_, _10565_, _05397_);
  not (_10639_, _10638_);
  nor (_10640_, _10628_, _04596_);
  and (_10641_, _10640_, _10639_);
  nor (_10642_, _10641_, _10637_);
  nor (_10643_, _10642_, _03773_);
  nor (_10644_, _10575_, _04594_);
  and (_10645_, _10644_, _10639_);
  nor (_10646_, _10645_, _03653_);
  not (_10647_, _10646_);
  nor (_10648_, _10647_, _10643_);
  nor (_10649_, _05959_, _10566_);
  or (_10650_, _10565_, _04608_);
  nor (_10651_, _10650_, _10649_);
  or (_10652_, _10651_, _03786_);
  nor (_10653_, _10652_, _10648_);
  nor (_10654_, _06457_, _10566_);
  nor (_10655_, _10654_, _10565_);
  nor (_10656_, _10655_, _04606_);
  or (_10657_, _10656_, _10653_);
  and (_10658_, _10657_, _04260_);
  nor (_10659_, _10581_, _04260_);
  or (_10660_, _10659_, _10658_);
  and (_10661_, _10660_, _03206_);
  nor (_10662_, _10572_, _03206_);
  or (_10663_, _10662_, _10661_);
  and (_10664_, _10663_, _03820_);
  and (_10665_, _05895_, _05345_);
  nor (_10666_, _10665_, _10565_);
  nor (_10667_, _10666_, _03820_);
  or (_10668_, _10667_, _10664_);
  or (_10669_, _10668_, _43231_);
  or (_10670_, _43227_, \oc8051_golden_model_1.SCON [7]);
  and (_10671_, _10670_, _41991_);
  and (_40760_, _10671_, _10669_);
  and (_10672_, _04952_, \oc8051_golden_model_1.SP [4]);
  and (_10673_, _10672_, \oc8051_golden_model_1.SP [5]);
  and (_10674_, _10673_, \oc8051_golden_model_1.SP [6]);
  nor (_10675_, _10674_, \oc8051_golden_model_1.SP [7]);
  and (_10676_, _10674_, \oc8051_golden_model_1.SP [7]);
  nor (_10677_, _10676_, _10675_);
  nor (_10679_, _10677_, _04625_);
  not (_10680_, _03792_);
  not (_10681_, \oc8051_golden_model_1.SP [7]);
  nor (_10682_, _05315_, _10681_);
  and (_10683_, _06458_, _05315_);
  nor (_10684_, _10683_, _10682_);
  nor (_10685_, _10684_, _04589_);
  not (_10686_, _05315_);
  nor (_10687_, _10686_, _05289_);
  nor (_10688_, _10687_, _10682_);
  nor (_10690_, _10688_, _06889_);
  or (_10691_, _10690_, _05969_);
  nor (_10692_, _04499_, _10681_);
  and (_10693_, _05315_, \oc8051_golden_model_1.ACC [7]);
  nor (_10694_, _10693_, _10682_);
  nor (_10695_, _10694_, _04500_);
  or (_10696_, _10695_, _10692_);
  and (_10697_, _10696_, _04868_);
  and (_10698_, _10677_, _03947_);
  nor (_10699_, _10698_, _10697_);
  nor (_10701_, _10699_, _03599_);
  and (_10702_, _06185_, _05315_);
  nor (_10703_, _10702_, _10682_);
  nor (_10704_, _10703_, _04515_);
  or (_10705_, _10704_, _10701_);
  and (_10706_, _10705_, _03257_);
  not (_10707_, _10677_);
  nor (_10708_, _10707_, _03257_);
  or (_10709_, _10708_, _10706_);
  and (_10710_, _10709_, _04524_);
  not (_10712_, \oc8051_golden_model_1.SP [6]);
  not (_10713_, \oc8051_golden_model_1.SP [5]);
  not (_10714_, \oc8051_golden_model_1.SP [4]);
  and (_10715_, _06074_, _10714_);
  and (_10716_, _10715_, _10713_);
  and (_10717_, _10716_, _10712_);
  and (_10718_, _10717_, _04079_);
  nor (_10719_, _10718_, _10681_);
  and (_10720_, _10718_, _10681_);
  nor (_10721_, _10720_, _10719_);
  nor (_10723_, _10721_, _04524_);
  or (_10724_, _10723_, _10710_);
  and (_10725_, _10724_, _03611_);
  nor (_10726_, _10694_, _03611_);
  or (_10727_, _10726_, _10725_);
  and (_10728_, _10727_, _04650_);
  not (_10729_, _04856_);
  and (_10730_, _10674_, \oc8051_golden_model_1.SP [0]);
  nor (_10731_, _10730_, _10681_);
  and (_10732_, _10730_, _10681_);
  nor (_10734_, _10732_, _10731_);
  nor (_10735_, _10734_, _04650_);
  nor (_10736_, _10735_, _10729_);
  not (_10737_, _10736_);
  nor (_10738_, _10737_, _10728_);
  nor (_10739_, _10677_, _04856_);
  or (_10740_, _10739_, _07441_);
  nor (_10741_, _10740_, _10738_);
  nor (_10742_, _10741_, _10691_);
  and (_10743_, _06171_, _05315_);
  nor (_10745_, _10682_, _05970_);
  not (_10746_, _10745_);
  nor (_10747_, _10746_, _10743_);
  nor (_10748_, _10747_, _03644_);
  not (_10749_, _10748_);
  nor (_10750_, _10749_, _10742_);
  nor (_10751_, _06443_, _10686_);
  nor (_10752_, _10751_, _10682_);
  nor (_10753_, _10752_, _03275_);
  or (_10754_, _10753_, _03650_);
  or (_10755_, _10754_, _10750_);
  and (_10756_, _06247_, _05315_);
  nor (_10757_, _10756_, _10682_);
  nand (_10758_, _10757_, _03650_);
  and (_10759_, _10758_, _10755_);
  nor (_10760_, _10759_, _03227_);
  and (_10761_, _10707_, _03227_);
  nor (_10762_, _10761_, _10760_);
  nor (_10763_, _10762_, _03649_);
  and (_10764_, _05961_, _05315_);
  or (_10765_, _10682_, _04591_);
  nor (_10766_, _10765_, _10764_);
  or (_10767_, _10766_, _03778_);
  nor (_10768_, _10767_, _10763_);
  nor (_10769_, _10768_, _10685_);
  nor (_10770_, _10769_, _03655_);
  nor (_10771_, _10682_, _05397_);
  not (_10772_, _10771_);
  nor (_10773_, _10757_, _04596_);
  and (_10774_, _10773_, _10772_);
  nor (_10775_, _10774_, _10770_);
  nor (_10776_, _03773_, _03238_);
  not (_10777_, _10776_);
  nor (_10778_, _10777_, _10775_);
  and (_10779_, _10677_, _03238_);
  or (_10780_, _10771_, _04594_);
  nor (_10781_, _10780_, _10694_);
  nor (_10782_, _10781_, _10779_);
  and (_10783_, _10782_, _04608_);
  not (_10784_, _10783_);
  nor (_10785_, _10784_, _10778_);
  nor (_10786_, _05959_, _10686_);
  nor (_10787_, _10786_, _10682_);
  and (_10788_, _10787_, _03653_);
  nor (_10789_, _10788_, _10785_);
  and (_10790_, _10789_, _04606_);
  nor (_10791_, _06457_, _10686_);
  nor (_10792_, _10791_, _10682_);
  nor (_10793_, _10792_, _04606_);
  or (_10794_, _10793_, _10790_);
  and (_10795_, _10794_, _10680_);
  nor (_10796_, _03792_, _03248_);
  nor (_10797_, _10717_, \oc8051_golden_model_1.SP [7]);
  and (_10798_, _10717_, \oc8051_golden_model_1.SP [7]);
  nor (_10799_, _10798_, _10797_);
  nor (_10800_, _10799_, _03248_);
  nor (_10801_, _10800_, _10796_);
  nor (_10802_, _10801_, _10795_);
  and (_10803_, _10707_, _03248_);
  nor (_10804_, _10803_, _10802_);
  and (_10805_, _10804_, _03522_);
  and (_10806_, _10799_, _03521_);
  or (_10807_, _10806_, _10805_);
  and (_10808_, _10807_, _04260_);
  nor (_10809_, _10703_, _04260_);
  nor (_10810_, _10809_, _05047_);
  not (_10811_, _10810_);
  nor (_10812_, _10811_, _10808_);
  nor (_10813_, _10812_, _10679_);
  and (_10814_, _10813_, _03820_);
  and (_10815_, _05895_, _05315_);
  nor (_10816_, _10815_, _10682_);
  nor (_10817_, _10816_, _03820_);
  or (_10818_, _10817_, _10814_);
  or (_10819_, _10818_, _43231_);
  or (_10820_, _43227_, \oc8051_golden_model_1.SP [7]);
  and (_10821_, _10820_, _41991_);
  and (_40762_, _10821_, _10819_);
  not (_10822_, \oc8051_golden_model_1.TCON [7]);
  nor (_10823_, _05353_, _10822_);
  not (_10824_, _05353_);
  nor (_10825_, _10824_, _05289_);
  nor (_10826_, _10825_, _10823_);
  and (_10827_, _10826_, _07441_);
  nor (_10828_, _05997_, _10822_);
  and (_10829_, _06038_, _05997_);
  nor (_10830_, _10829_, _10828_);
  nor (_10831_, _10830_, _03512_);
  and (_10832_, _05353_, \oc8051_golden_model_1.ACC [7]);
  nor (_10833_, _10832_, _10823_);
  nor (_10834_, _10833_, _04500_);
  nor (_10835_, _04499_, _10822_);
  or (_10836_, _10835_, _10834_);
  and (_10837_, _10836_, _04515_);
  and (_10838_, _06185_, _05353_);
  nor (_10839_, _10838_, _10823_);
  nor (_10840_, _10839_, _04515_);
  or (_10841_, _10840_, _10837_);
  and (_10842_, _10841_, _03516_);
  and (_10843_, _06042_, _05997_);
  nor (_10844_, _10843_, _10828_);
  nor (_10845_, _10844_, _03516_);
  or (_10846_, _10845_, _03597_);
  or (_10847_, _10846_, _10842_);
  nand (_10848_, _10826_, _03597_);
  and (_10849_, _10848_, _10847_);
  and (_10850_, _10849_, _03611_);
  nor (_10851_, _10833_, _03611_);
  or (_10852_, _10851_, _10850_);
  and (_10853_, _10852_, _03512_);
  nor (_10854_, _10853_, _10831_);
  nor (_10855_, _10854_, _03504_);
  and (_10856_, _06217_, _05997_);
  nor (_10857_, _10856_, _10828_);
  nor (_10858_, _10857_, _03505_);
  nor (_10859_, _10858_, _10855_);
  nor (_10860_, _10859_, _03500_);
  not (_10861_, _05997_);
  nor (_10862_, _06026_, _10861_);
  nor (_10863_, _10862_, _10828_);
  nor (_10864_, _10863_, _03501_);
  nor (_10865_, _10864_, _07441_);
  not (_10866_, _10865_);
  nor (_10867_, _10866_, _10860_);
  nor (_10868_, _10867_, _10827_);
  nor (_10869_, _10868_, _05969_);
  and (_10870_, _06171_, _05353_);
  nor (_10871_, _10823_, _05970_);
  not (_10872_, _10871_);
  nor (_10873_, _10872_, _10870_);
  nor (_10874_, _10873_, _03644_);
  not (_10875_, _10874_);
  nor (_10876_, _10875_, _10869_);
  nor (_10877_, _06443_, _10824_);
  nor (_10878_, _10877_, _10823_);
  nor (_10879_, _10878_, _03275_);
  or (_10880_, _10879_, _08861_);
  or (_10881_, _10880_, _10876_);
  and (_10882_, _05961_, _05353_);
  or (_10883_, _10823_, _04591_);
  or (_10884_, _10883_, _10882_);
  and (_10885_, _06247_, _05353_);
  nor (_10886_, _10885_, _10823_);
  and (_10887_, _10886_, _03650_);
  nor (_10888_, _10887_, _03778_);
  and (_10889_, _10888_, _10884_);
  and (_10890_, _10889_, _10881_);
  and (_10891_, _06458_, _05353_);
  nor (_10892_, _10891_, _10823_);
  nor (_10893_, _10892_, _04589_);
  nor (_10894_, _10893_, _10890_);
  nor (_10895_, _10894_, _03655_);
  nor (_10896_, _10823_, _05397_);
  not (_10897_, _10896_);
  nor (_10898_, _10886_, _04596_);
  and (_10899_, _10898_, _10897_);
  nor (_10900_, _10899_, _10895_);
  nor (_10901_, _10900_, _03773_);
  nor (_10902_, _10833_, _04594_);
  and (_10903_, _10902_, _10897_);
  or (_10904_, _10903_, _10901_);
  and (_10905_, _10904_, _04608_);
  nor (_10906_, _05959_, _10824_);
  nor (_10907_, _10906_, _10823_);
  nor (_10908_, _10907_, _04608_);
  or (_10909_, _10908_, _10905_);
  and (_10910_, _10909_, _04606_);
  nor (_10911_, _06457_, _10824_);
  nor (_10912_, _10911_, _10823_);
  nor (_10913_, _10912_, _04606_);
  or (_10914_, _10913_, _10910_);
  and (_10915_, _10914_, _04260_);
  nor (_10916_, _10839_, _04260_);
  or (_10917_, _10916_, _10915_);
  and (_10918_, _10917_, _03206_);
  nor (_10919_, _10830_, _03206_);
  or (_10920_, _10919_, _10918_);
  and (_10921_, _10920_, _03820_);
  and (_10922_, _05895_, _05353_);
  nor (_10923_, _10922_, _10823_);
  nor (_10924_, _10923_, _03820_);
  or (_10925_, _10924_, _10921_);
  or (_10926_, _10925_, _43231_);
  or (_10927_, _43227_, \oc8051_golden_model_1.TCON [7]);
  and (_10928_, _10927_, _41991_);
  and (_40763_, _10928_, _10926_);
  not (_10929_, \oc8051_golden_model_1.TH0 [7]);
  nor (_10930_, _05304_, _10929_);
  not (_10931_, _05304_);
  nor (_10932_, _06457_, _10931_);
  nor (_10933_, _10932_, _10930_);
  nor (_10934_, _10933_, _04606_);
  and (_10935_, _06247_, _05304_);
  nor (_10936_, _10935_, _10930_);
  and (_10937_, _10936_, _03650_);
  nor (_10938_, _10931_, _05289_);
  nor (_10939_, _10938_, _10930_);
  and (_10940_, _10939_, _07441_);
  and (_10941_, _05304_, \oc8051_golden_model_1.ACC [7]);
  nor (_10942_, _10941_, _10930_);
  nor (_10943_, _10942_, _04500_);
  nor (_10944_, _04499_, _10929_);
  or (_10945_, _10944_, _10943_);
  and (_10946_, _10945_, _04515_);
  and (_10947_, _06185_, _05304_);
  nor (_10948_, _10947_, _10930_);
  nor (_10949_, _10948_, _04515_);
  or (_10950_, _10949_, _10946_);
  and (_10951_, _10950_, _04524_);
  nor (_10952_, _10939_, _04524_);
  nor (_10953_, _10952_, _10951_);
  nor (_10954_, _10953_, _03603_);
  nor (_10955_, _10942_, _03611_);
  nor (_10956_, _10955_, _07441_);
  not (_10957_, _10956_);
  nor (_10958_, _10957_, _10954_);
  nor (_10959_, _10958_, _10940_);
  nor (_10960_, _10959_, _05969_);
  and (_10961_, _06171_, _05304_);
  nor (_10962_, _10930_, _05970_);
  not (_10963_, _10962_);
  nor (_10964_, _10963_, _10961_);
  or (_10965_, _10964_, _03644_);
  nor (_10966_, _10965_, _10960_);
  nor (_10967_, _06443_, _10931_);
  nor (_10968_, _10967_, _10930_);
  nor (_10969_, _10968_, _03275_);
  or (_10970_, _10969_, _03650_);
  nor (_10971_, _10970_, _10966_);
  nor (_10972_, _10971_, _10937_);
  or (_10973_, _10972_, _03649_);
  and (_10974_, _05961_, _05304_);
  or (_10975_, _10974_, _10930_);
  or (_10976_, _10975_, _04591_);
  and (_10977_, _10976_, _04589_);
  and (_10978_, _10977_, _10973_);
  and (_10979_, _06458_, _05304_);
  nor (_10980_, _10979_, _10930_);
  nor (_10981_, _10980_, _04589_);
  nor (_10982_, _10981_, _10978_);
  nor (_10983_, _10982_, _03655_);
  nor (_10984_, _10930_, _05397_);
  not (_10985_, _10984_);
  nor (_10986_, _10936_, _04596_);
  and (_10987_, _10986_, _10985_);
  nor (_10988_, _10987_, _10983_);
  nor (_10989_, _10988_, _03773_);
  nor (_10990_, _10942_, _04594_);
  and (_10991_, _10990_, _10985_);
  or (_10992_, _10991_, _10989_);
  and (_10993_, _10992_, _04608_);
  nor (_10994_, _05959_, _10931_);
  nor (_10995_, _10994_, _10930_);
  nor (_10996_, _10995_, _04608_);
  or (_10997_, _10996_, _10993_);
  and (_10998_, _10997_, _04606_);
  nor (_10999_, _10998_, _10934_);
  nor (_11000_, _10999_, _03809_);
  nor (_11001_, _10948_, _04260_);
  or (_11002_, _11001_, _03816_);
  nor (_11003_, _11002_, _11000_);
  and (_11004_, _05895_, _05304_);
  or (_11005_, _10930_, _03820_);
  nor (_11006_, _11005_, _11004_);
  nor (_11007_, _11006_, _11003_);
  or (_11008_, _11007_, _43231_);
  or (_11009_, _43227_, \oc8051_golden_model_1.TH0 [7]);
  and (_11010_, _11009_, _41991_);
  and (_40764_, _11010_, _11008_);
  not (_11011_, \oc8051_golden_model_1.TH1 [7]);
  nor (_11012_, _05356_, _11011_);
  not (_11013_, _05356_);
  nor (_11014_, _06457_, _11013_);
  nor (_11015_, _11014_, _11012_);
  nor (_11016_, _11015_, _04606_);
  and (_11017_, _06247_, _05356_);
  nor (_11018_, _11017_, _11012_);
  and (_11019_, _11018_, _03650_);
  nor (_11020_, _11013_, _05289_);
  nor (_11021_, _11020_, _11012_);
  and (_11022_, _11021_, _07441_);
  and (_11023_, _05356_, \oc8051_golden_model_1.ACC [7]);
  nor (_11024_, _11023_, _11012_);
  nor (_11025_, _11024_, _04500_);
  nor (_11026_, _04499_, _11011_);
  or (_11027_, _11026_, _11025_);
  and (_11028_, _11027_, _04515_);
  and (_11029_, _06185_, _05356_);
  nor (_11030_, _11029_, _11012_);
  nor (_11031_, _11030_, _04515_);
  or (_11032_, _11031_, _11028_);
  and (_11033_, _11032_, _04524_);
  nor (_11034_, _11021_, _04524_);
  nor (_11035_, _11034_, _11033_);
  nor (_11036_, _11035_, _03603_);
  nor (_11037_, _11024_, _03611_);
  nor (_11038_, _11037_, _07441_);
  not (_11039_, _11038_);
  nor (_11040_, _11039_, _11036_);
  nor (_11041_, _11040_, _11022_);
  nor (_11042_, _11041_, _05969_);
  and (_11043_, _06171_, _05356_);
  nor (_11044_, _11012_, _05970_);
  not (_11045_, _11044_);
  nor (_11046_, _11045_, _11043_);
  or (_11047_, _11046_, _03644_);
  nor (_11048_, _11047_, _11042_);
  nor (_11049_, _06443_, _11013_);
  nor (_11050_, _11049_, _11012_);
  nor (_11051_, _11050_, _03275_);
  or (_11052_, _11051_, _03650_);
  nor (_11053_, _11052_, _11048_);
  nor (_11054_, _11053_, _11019_);
  or (_11055_, _11054_, _03649_);
  and (_11056_, _05961_, _05356_);
  or (_11057_, _11056_, _11012_);
  or (_11058_, _11057_, _04591_);
  and (_11059_, _11058_, _04589_);
  and (_11060_, _11059_, _11055_);
  and (_11061_, _06458_, _05356_);
  nor (_11062_, _11061_, _11012_);
  nor (_11063_, _11062_, _04589_);
  nor (_11064_, _11063_, _11060_);
  nor (_11065_, _11064_, _03655_);
  nor (_11066_, _11012_, _05397_);
  not (_11067_, _11066_);
  nor (_11068_, _11018_, _04596_);
  and (_11069_, _11068_, _11067_);
  nor (_11070_, _11069_, _11065_);
  nor (_11071_, _11070_, _03773_);
  nor (_11072_, _11024_, _04594_);
  and (_11073_, _11072_, _11067_);
  or (_11074_, _11073_, _11071_);
  and (_11075_, _11074_, _04608_);
  nor (_11076_, _05959_, _11013_);
  nor (_11077_, _11076_, _11012_);
  nor (_11078_, _11077_, _04608_);
  or (_11079_, _11078_, _11075_);
  and (_11080_, _11079_, _04606_);
  nor (_11081_, _11080_, _11016_);
  nor (_11082_, _11081_, _03809_);
  nor (_11083_, _11030_, _04260_);
  or (_11084_, _11083_, _03816_);
  nor (_11085_, _11084_, _11082_);
  and (_11086_, _05895_, _05356_);
  or (_11087_, _11012_, _03820_);
  nor (_11088_, _11087_, _11086_);
  nor (_11089_, _11088_, _11085_);
  or (_11090_, _11089_, _43231_);
  or (_11091_, _43227_, \oc8051_golden_model_1.TH1 [7]);
  and (_11092_, _11091_, _41991_);
  and (_40765_, _11092_, _11090_);
  not (_11093_, \oc8051_golden_model_1.TL0 [7]);
  nor (_11094_, _05350_, _11093_);
  not (_11095_, _05350_);
  nor (_11096_, _06457_, _11095_);
  nor (_11097_, _11096_, _11094_);
  nor (_11098_, _11097_, _04606_);
  and (_11099_, _06247_, _05350_);
  nor (_11100_, _11099_, _11094_);
  and (_11101_, _11100_, _03650_);
  nor (_11102_, _11095_, _05289_);
  nor (_11103_, _11102_, _11094_);
  and (_11104_, _11103_, _07441_);
  and (_11105_, _05350_, \oc8051_golden_model_1.ACC [7]);
  nor (_11106_, _11105_, _11094_);
  nor (_11107_, _11106_, _04500_);
  nor (_11108_, _04499_, _11093_);
  or (_11109_, _11108_, _11107_);
  and (_11110_, _11109_, _04515_);
  and (_11111_, _06185_, _05350_);
  nor (_11112_, _11111_, _11094_);
  nor (_11113_, _11112_, _04515_);
  or (_11114_, _11113_, _11110_);
  and (_11115_, _11114_, _04524_);
  nor (_11116_, _11103_, _04524_);
  nor (_11117_, _11116_, _11115_);
  nor (_11118_, _11117_, _03603_);
  nor (_11119_, _11106_, _03611_);
  nor (_11120_, _11119_, _07441_);
  not (_11121_, _11120_);
  nor (_11122_, _11121_, _11118_);
  nor (_11123_, _11122_, _11104_);
  nor (_11124_, _11123_, _05969_);
  and (_11125_, _06171_, _05350_);
  nor (_11126_, _11094_, _05970_);
  not (_11127_, _11126_);
  nor (_11128_, _11127_, _11125_);
  or (_11129_, _11128_, _03644_);
  nor (_11130_, _11129_, _11124_);
  nor (_11131_, _06443_, _11095_);
  nor (_11132_, _11131_, _11094_);
  nor (_11133_, _11132_, _03275_);
  or (_11134_, _11133_, _03650_);
  nor (_11135_, _11134_, _11130_);
  nor (_11136_, _11135_, _11101_);
  or (_11137_, _11136_, _03649_);
  and (_11138_, _05961_, _05350_);
  or (_11139_, _11138_, _11094_);
  or (_11140_, _11139_, _04591_);
  and (_11141_, _11140_, _04589_);
  and (_11142_, _11141_, _11137_);
  and (_11143_, _06458_, _05350_);
  nor (_11144_, _11143_, _11094_);
  nor (_11145_, _11144_, _04589_);
  nor (_11146_, _11145_, _11142_);
  nor (_11147_, _11146_, _03655_);
  nor (_11148_, _11094_, _05397_);
  not (_11149_, _11148_);
  nor (_11150_, _11100_, _04596_);
  and (_11151_, _11150_, _11149_);
  nor (_11152_, _11151_, _11147_);
  nor (_11153_, _11152_, _03773_);
  nor (_11154_, _11106_, _04594_);
  and (_11155_, _11154_, _11149_);
  nor (_11156_, _11155_, _03653_);
  not (_11157_, _11156_);
  nor (_11158_, _11157_, _11153_);
  nor (_11159_, _05959_, _11095_);
  or (_11160_, _11094_, _04608_);
  nor (_11161_, _11160_, _11159_);
  or (_11162_, _11161_, _03786_);
  nor (_11163_, _11162_, _11158_);
  nor (_11164_, _11163_, _11098_);
  nor (_11165_, _11164_, _03809_);
  nor (_11166_, _11112_, _04260_);
  or (_11167_, _11166_, _03816_);
  nor (_11168_, _11167_, _11165_);
  and (_11169_, _05895_, _05350_);
  nor (_11170_, _11169_, _11094_);
  and (_11171_, _11170_, _03816_);
  nor (_11172_, _11171_, _11168_);
  or (_11173_, _11172_, _43231_);
  or (_11174_, _43227_, \oc8051_golden_model_1.TL0 [7]);
  and (_11175_, _11174_, _41991_);
  and (_40766_, _11175_, _11173_);
  not (_11176_, \oc8051_golden_model_1.TL1 [7]);
  nor (_11177_, _05309_, _11176_);
  not (_11178_, _05309_);
  nor (_11179_, _06457_, _11178_);
  nor (_11180_, _11179_, _11177_);
  nor (_11181_, _11180_, _04606_);
  and (_11182_, _06247_, _05309_);
  nor (_11183_, _11182_, _11177_);
  and (_11184_, _11183_, _03650_);
  nor (_11185_, _11178_, _05289_);
  nor (_11186_, _11185_, _11177_);
  and (_11187_, _11186_, _07441_);
  and (_11188_, _05309_, \oc8051_golden_model_1.ACC [7]);
  nor (_11189_, _11188_, _11177_);
  nor (_11190_, _11189_, _04500_);
  nor (_11191_, _04499_, _11176_);
  or (_11192_, _11191_, _11190_);
  and (_11193_, _11192_, _04515_);
  and (_11194_, _06185_, _05309_);
  nor (_11195_, _11194_, _11177_);
  nor (_11196_, _11195_, _04515_);
  or (_11197_, _11196_, _11193_);
  and (_11198_, _11197_, _04524_);
  nor (_11199_, _11186_, _04524_);
  nor (_11200_, _11199_, _11198_);
  nor (_11201_, _11200_, _03603_);
  nor (_11202_, _11189_, _03611_);
  nor (_11203_, _11202_, _07441_);
  not (_11204_, _11203_);
  nor (_11205_, _11204_, _11201_);
  nor (_11206_, _11205_, _11187_);
  nor (_11207_, _11206_, _05969_);
  and (_11208_, _06171_, _05309_);
  nor (_11209_, _11177_, _05970_);
  not (_11210_, _11209_);
  nor (_11211_, _11210_, _11208_);
  or (_11212_, _11211_, _03644_);
  nor (_11213_, _11212_, _11207_);
  nor (_11214_, _06443_, _11178_);
  nor (_11215_, _11214_, _11177_);
  nor (_11216_, _11215_, _03275_);
  or (_11217_, _11216_, _03650_);
  nor (_11218_, _11217_, _11213_);
  nor (_11219_, _11218_, _11184_);
  or (_11220_, _11219_, _03649_);
  and (_11221_, _05961_, _05309_);
  or (_11222_, _11221_, _11177_);
  or (_11223_, _11222_, _04591_);
  and (_11224_, _11223_, _04589_);
  and (_11225_, _11224_, _11220_);
  and (_11226_, _06458_, _05309_);
  nor (_11227_, _11226_, _11177_);
  nor (_11228_, _11227_, _04589_);
  nor (_11229_, _11228_, _11225_);
  nor (_11230_, _11229_, _03655_);
  nor (_11231_, _11177_, _05397_);
  not (_11232_, _11231_);
  nor (_11233_, _11183_, _04596_);
  and (_11234_, _11233_, _11232_);
  nor (_11235_, _11234_, _11230_);
  nor (_11236_, _11235_, _03773_);
  nor (_11237_, _11189_, _04594_);
  and (_11238_, _11237_, _11232_);
  nor (_11239_, _11238_, _03653_);
  not (_11240_, _11239_);
  nor (_11241_, _11240_, _11236_);
  nor (_11242_, _05959_, _11178_);
  or (_11243_, _11177_, _04608_);
  nor (_11244_, _11243_, _11242_);
  or (_11245_, _11244_, _03786_);
  nor (_11246_, _11245_, _11241_);
  nor (_11247_, _11246_, _11181_);
  nor (_11248_, _11247_, _03809_);
  nor (_11249_, _11195_, _04260_);
  or (_11250_, _11249_, _03816_);
  nor (_11251_, _11250_, _11248_);
  and (_11252_, _05895_, _05309_);
  or (_11253_, _11177_, _03820_);
  nor (_11254_, _11253_, _11252_);
  nor (_11255_, _11254_, _11251_);
  or (_11256_, _11255_, _43231_);
  or (_11257_, _43227_, \oc8051_golden_model_1.TL1 [7]);
  and (_11258_, _11257_, _41991_);
  and (_40768_, _11258_, _11256_);
  not (_11259_, \oc8051_golden_model_1.TMOD [7]);
  nor (_11260_, _05343_, _11259_);
  not (_11261_, _05343_);
  nor (_11262_, _06457_, _11261_);
  nor (_11263_, _11262_, _11260_);
  nor (_11264_, _11263_, _04606_);
  and (_11265_, _06247_, _05343_);
  nor (_11266_, _11265_, _11260_);
  and (_11267_, _11266_, _03650_);
  nor (_11268_, _11261_, _05289_);
  nor (_11269_, _11268_, _11260_);
  and (_11270_, _11269_, _07441_);
  and (_11271_, _05343_, \oc8051_golden_model_1.ACC [7]);
  nor (_11272_, _11271_, _11260_);
  nor (_11273_, _11272_, _03611_);
  nor (_11274_, _11272_, _04500_);
  nor (_11275_, _04499_, _11259_);
  or (_11276_, _11275_, _11274_);
  and (_11277_, _11276_, _04515_);
  and (_11278_, _06185_, _05343_);
  nor (_11279_, _11278_, _11260_);
  nor (_11280_, _11279_, _04515_);
  or (_11281_, _11280_, _11277_);
  and (_11282_, _11281_, _04524_);
  nor (_11283_, _11269_, _04524_);
  nor (_11284_, _11283_, _11282_);
  nor (_11285_, _11284_, _03603_);
  or (_11286_, _11285_, _07441_);
  nor (_11287_, _11286_, _11273_);
  nor (_11288_, _11287_, _11270_);
  nor (_11289_, _11288_, _05969_);
  and (_11290_, _06171_, _05343_);
  nor (_11291_, _11260_, _05970_);
  not (_11292_, _11291_);
  nor (_11293_, _11292_, _11290_);
  or (_11294_, _11293_, _03644_);
  nor (_11295_, _11294_, _11289_);
  nor (_11296_, _06443_, _11261_);
  nor (_11297_, _11296_, _11260_);
  nor (_11298_, _11297_, _03275_);
  or (_11299_, _11298_, _03650_);
  nor (_11300_, _11299_, _11295_);
  nor (_11301_, _11300_, _11267_);
  or (_11302_, _11301_, _03649_);
  and (_11303_, _05961_, _05343_);
  or (_11304_, _11303_, _11260_);
  or (_11305_, _11304_, _04591_);
  and (_11306_, _11305_, _04589_);
  and (_11307_, _11306_, _11302_);
  and (_11308_, _06458_, _05343_);
  nor (_11309_, _11308_, _11260_);
  nor (_11310_, _11309_, _04589_);
  nor (_11311_, _11310_, _11307_);
  nor (_11312_, _11311_, _03655_);
  nor (_11313_, _11260_, _05397_);
  not (_11314_, _11313_);
  nor (_11315_, _11266_, _04596_);
  and (_11316_, _11315_, _11314_);
  nor (_11317_, _11316_, _11312_);
  nor (_11318_, _11317_, _03773_);
  nor (_11319_, _11272_, _04594_);
  and (_11320_, _11319_, _11314_);
  or (_11321_, _11320_, _11318_);
  and (_11322_, _11321_, _04608_);
  nor (_11323_, _05959_, _11261_);
  nor (_11324_, _11323_, _11260_);
  nor (_11325_, _11324_, _04608_);
  or (_11326_, _11325_, _11322_);
  and (_11327_, _11326_, _04606_);
  nor (_11328_, _11327_, _11264_);
  nor (_11329_, _11328_, _03809_);
  nor (_11330_, _11279_, _04260_);
  or (_11331_, _11330_, _03816_);
  nor (_11332_, _11331_, _11329_);
  and (_11333_, _05895_, _05343_);
  or (_11334_, _11260_, _03820_);
  nor (_11335_, _11334_, _11333_);
  nor (_11336_, _11335_, _11332_);
  or (_11337_, _11336_, _43231_);
  or (_11338_, _43227_, \oc8051_golden_model_1.TMOD [7]);
  and (_11339_, _11338_, _41991_);
  and (_40769_, _11339_, _11337_);
  not (_11340_, _02925_);
  and (_11341_, _05916_, _11340_);
  and (_11342_, _11341_, \oc8051_golden_model_1.PC [7]);
  and (_11343_, _11342_, \oc8051_golden_model_1.PC [8]);
  and (_11344_, _11343_, \oc8051_golden_model_1.PC [9]);
  and (_11345_, _11344_, \oc8051_golden_model_1.PC [10]);
  and (_11346_, _11345_, \oc8051_golden_model_1.PC [11]);
  and (_11347_, _11346_, \oc8051_golden_model_1.PC [12]);
  and (_11348_, _11347_, \oc8051_golden_model_1.PC [13]);
  and (_11349_, _11348_, \oc8051_golden_model_1.PC [14]);
  or (_11350_, _11349_, \oc8051_golden_model_1.PC [15]);
  nand (_11351_, _11349_, \oc8051_golden_model_1.PC [15]);
  and (_11352_, _11351_, _11350_);
  and (_11353_, _09696_, _10369_);
  or (_11354_, _11353_, _11352_);
  and (_11355_, _08541_, _07933_);
  or (_11356_, _11355_, _11352_);
  nor (_11357_, _08524_, _03784_);
  not (_11358_, _11357_);
  not (_11359_, _04208_);
  nor (_11360_, _04377_, _03954_);
  and (_11361_, _11360_, _11359_);
  or (_11362_, _11361_, _11352_);
  and (_11363_, _03237_, _03204_);
  not (_11364_, _11363_);
  or (_11365_, _10776_, _06874_);
  and (_11366_, _11365_, _11364_);
  nor (_11367_, _07942_, _03771_);
  not (_11368_, _11367_);
  nor (_11369_, _04814_, _04194_);
  nor (_11370_, _08490_, _11369_);
  or (_11371_, _11370_, _11352_);
  and (_11372_, _03219_, _03204_);
  not (_11373_, _11372_);
  nor (_11374_, _03562_, _03220_);
  or (_11375_, _11374_, _06874_);
  and (_11376_, _11375_, _11373_);
  not (_11377_, _06867_);
  nor (_11378_, _11377_, _03275_);
  nor (_11379_, _08160_, _03635_);
  not (_11380_, _11379_);
  and (_11381_, _08037_, _08128_);
  or (_11382_, _11381_, _11352_);
  nor (_11383_, _03274_, _03264_);
  not (_11384_, _11383_);
  nor (_11385_, _08880_, _06919_);
  and (_11386_, _11385_, _11384_);
  not (_11387_, _11386_);
  and (_11388_, _11387_, _11352_);
  not (_11389_, _10096_);
  and (_11390_, _06874_, _03603_);
  nor (_11391_, _09965_, _08063_);
  not (_11392_, _11391_);
  and (_11393_, _05744_, _05698_);
  and (_11394_, _06179_, _11393_);
  and (_11395_, _05490_, _05396_);
  and (_11396_, _11395_, _06176_);
  and (_11397_, _11396_, _11394_);
  and (_11398_, _05920_, \oc8051_golden_model_1.PC [8]);
  and (_11399_, _11398_, \oc8051_golden_model_1.PC [9]);
  and (_11400_, _11399_, \oc8051_golden_model_1.PC [10]);
  and (_11401_, _11400_, \oc8051_golden_model_1.PC [11]);
  and (_11402_, _11401_, \oc8051_golden_model_1.PC [12]);
  and (_11403_, _11402_, \oc8051_golden_model_1.PC [13]);
  and (_11404_, _11403_, \oc8051_golden_model_1.PC [14]);
  nor (_11405_, _11403_, \oc8051_golden_model_1.PC [14]);
  nor (_11406_, _11405_, _11404_);
  not (_11407_, _11406_);
  nor (_11408_, _11407_, _05958_);
  and (_11409_, _11407_, _05958_);
  nor (_11410_, _11409_, _11408_);
  not (_11411_, _11410_);
  nor (_11412_, _11402_, \oc8051_golden_model_1.PC [13]);
  nor (_11413_, _11412_, _11403_);
  not (_11414_, _11413_);
  nor (_11415_, _11414_, _05958_);
  and (_11416_, _11414_, _05958_);
  nor (_11417_, _11401_, \oc8051_golden_model_1.PC [12]);
  nor (_11418_, _11417_, _11402_);
  not (_11419_, _11418_);
  nor (_11420_, _11419_, _05958_);
  nor (_11421_, _11399_, \oc8051_golden_model_1.PC [10]);
  nor (_11422_, _11421_, _11400_);
  not (_11423_, _11422_);
  nor (_11424_, _11423_, _05958_);
  not (_11425_, _11424_);
  nor (_11426_, _11400_, \oc8051_golden_model_1.PC [11]);
  nor (_11427_, _11426_, _11401_);
  not (_11428_, _11427_);
  nor (_11429_, _11428_, _05958_);
  and (_11430_, _11428_, _05958_);
  nor (_11431_, _11430_, _11429_);
  and (_11432_, _11423_, _05958_);
  nor (_11433_, _11432_, _11424_);
  and (_11434_, _11433_, _11431_);
  nor (_11435_, _11398_, \oc8051_golden_model_1.PC [9]);
  nor (_11436_, _11435_, _11399_);
  not (_11437_, _11436_);
  nor (_11438_, _11437_, _05958_);
  and (_11439_, _11437_, _05958_);
  nor (_11440_, _11439_, _11438_);
  nor (_11441_, _05958_, _05923_);
  and (_11442_, _05958_, _05923_);
  and (_11443_, _05918_, _05915_);
  nor (_11444_, _11443_, \oc8051_golden_model_1.PC [6]);
  nor (_11445_, _11444_, _05919_);
  not (_11446_, _11445_);
  nor (_11447_, _11446_, _06281_);
  and (_11448_, _11446_, _06281_);
  nor (_11449_, _11448_, _11447_);
  not (_11450_, _11449_);
  and (_11451_, _05918_, \oc8051_golden_model_1.PC [4]);
  nor (_11452_, _11451_, \oc8051_golden_model_1.PC [5]);
  nor (_11453_, _11452_, _11443_);
  not (_11454_, _11453_);
  nor (_11455_, _11454_, _06313_);
  and (_11456_, _11454_, _06313_);
  nor (_11457_, _05918_, \oc8051_golden_model_1.PC [4]);
  nor (_11458_, _11457_, _11451_);
  not (_11459_, _11458_);
  nor (_11460_, _11459_, _06344_);
  nor (_11461_, _05917_, \oc8051_golden_model_1.PC [3]);
  nor (_11462_, _11461_, _05918_);
  not (_11463_, _11462_);
  nor (_11464_, _11463_, _03766_);
  and (_11465_, _11463_, _03766_);
  nor (_11466_, _02942_, \oc8051_golden_model_1.PC [2]);
  nor (_11467_, _11466_, _05917_);
  not (_11468_, _11467_);
  nor (_11469_, _11468_, _03943_);
  not (_11470_, _03321_);
  nor (_11471_, _04347_, _11470_);
  nor (_11472_, _04172_, \oc8051_golden_model_1.PC [0]);
  and (_11473_, _04347_, _11470_);
  nor (_11474_, _11473_, _11471_);
  and (_11475_, _11474_, _11472_);
  nor (_11476_, _11475_, _11471_);
  and (_11477_, _11468_, _03943_);
  nor (_11478_, _11477_, _11469_);
  not (_11479_, _11478_);
  nor (_11480_, _11479_, _11476_);
  nor (_11481_, _11480_, _11469_);
  nor (_11482_, _11481_, _11465_);
  nor (_11483_, _11482_, _11464_);
  and (_11484_, _11459_, _06344_);
  nor (_11485_, _11484_, _11460_);
  not (_11486_, _11485_);
  nor (_11487_, _11486_, _11483_);
  nor (_11488_, _11487_, _11460_);
  nor (_11489_, _11488_, _11456_);
  nor (_11490_, _11489_, _11455_);
  nor (_11491_, _11490_, _11450_);
  nor (_11492_, _11491_, _11447_);
  nor (_11493_, _11492_, _11442_);
  or (_11494_, _11493_, _11441_);
  nor (_11495_, _05920_, \oc8051_golden_model_1.PC [8]);
  nor (_11496_, _11495_, _11398_);
  not (_11497_, _11496_);
  nor (_11498_, _11497_, _05958_);
  and (_11499_, _11497_, _05958_);
  nor (_11500_, _11499_, _11498_);
  and (_11501_, _11500_, _11494_);
  and (_11502_, _11501_, _11440_);
  and (_11503_, _11502_, _11434_);
  nor (_11504_, _11498_, _11438_);
  not (_11505_, _11504_);
  and (_11506_, _11505_, _11434_);
  or (_11507_, _11506_, _11429_);
  nor (_11508_, _11507_, _11503_);
  and (_11509_, _11508_, _11425_);
  not (_11510_, _11509_);
  and (_11511_, _11419_, _05958_);
  nor (_11512_, _11511_, _11420_);
  and (_11513_, _11512_, _11510_);
  nor (_11514_, _11513_, _11420_);
  nor (_11515_, _11514_, _11416_);
  nor (_11516_, _11515_, _11415_);
  nor (_11517_, _11516_, _11411_);
  nor (_11518_, _11517_, _11408_);
  and (_11519_, _11377_, _05958_);
  nor (_11520_, _11377_, _05958_);
  nor (_11521_, _11520_, _11519_);
  and (_11522_, _11521_, _11518_);
  nor (_11523_, _11521_, _11518_);
  or (_11524_, _11523_, _11522_);
  or (_11525_, _11524_, _11397_);
  nand (_11526_, _11396_, _11394_);
  or (_11527_, _11526_, _06867_);
  and (_11528_, _11527_, _11525_);
  or (_11529_, _11528_, _04515_);
  or (_11530_, _06874_, _03948_);
  nor (_11531_, _04834_, _04821_);
  not (_11532_, _11531_);
  and (_11533_, _11532_, _11352_);
  and (_11534_, _11531_, \oc8051_golden_model_1.PC [15]);
  or (_11535_, _11534_, _04499_);
  and (_11536_, _03946_, _03170_);
  not (_11537_, _11536_);
  nor (_11538_, _04493_, _03261_);
  not (_11539_, _11538_);
  and (_11540_, _11539_, _08048_);
  and (_11541_, _11540_, _11537_);
  and (_11542_, _11541_, _11535_);
  or (_11543_, _11542_, _11533_);
  and (_11544_, _11543_, _11530_);
  not (_11545_, _11541_);
  and (_11546_, _11545_, _11352_);
  nand (_11547_, _06874_, _03947_);
  nand (_11548_, _11547_, _06054_);
  or (_11549_, _11548_, _11546_);
  or (_11550_, _11549_, _11544_);
  and (_11551_, _06046_, _06044_);
  and (_11552_, _04699_, _04491_);
  and (_11553_, _11552_, _05905_);
  and (_11554_, _11553_, _11551_);
  and (_11555_, _11554_, _06874_);
  nand (_11556_, _11553_, _11551_);
  and (_11557_, _06057_, \oc8051_golden_model_1.PC [8]);
  and (_11558_, _11557_, \oc8051_golden_model_1.PC [9]);
  and (_11559_, _11558_, \oc8051_golden_model_1.PC [10]);
  and (_11560_, _11559_, \oc8051_golden_model_1.PC [11]);
  and (_11561_, _11560_, \oc8051_golden_model_1.PC [12]);
  and (_11562_, _11561_, \oc8051_golden_model_1.PC [13]);
  and (_11563_, _11562_, \oc8051_golden_model_1.PC [14]);
  nor (_11564_, _11562_, \oc8051_golden_model_1.PC [14]);
  nor (_11565_, _11564_, _11563_);
  and (_11566_, _11565_, _03463_);
  nor (_11567_, _11565_, _03463_);
  nor (_11568_, _11567_, _11566_);
  not (_11569_, _11568_);
  nor (_11570_, _11561_, \oc8051_golden_model_1.PC [13]);
  nor (_11571_, _11570_, _11562_);
  and (_11572_, _11571_, _03463_);
  nor (_11573_, _11571_, _03463_);
  nor (_11574_, _11560_, \oc8051_golden_model_1.PC [12]);
  nor (_11575_, _11574_, _11561_);
  and (_11576_, _11575_, _03463_);
  nor (_11577_, _11558_, \oc8051_golden_model_1.PC [10]);
  nor (_11578_, _11577_, _11559_);
  and (_11579_, _11578_, _03463_);
  not (_11580_, _11579_);
  nor (_11581_, _11559_, \oc8051_golden_model_1.PC [11]);
  nor (_11582_, _11581_, _11560_);
  and (_11583_, _11582_, _03463_);
  nor (_11584_, _11582_, _03463_);
  nor (_11585_, _11584_, _11583_);
  nor (_11586_, _11578_, _03463_);
  nor (_11587_, _11586_, _11579_);
  and (_11588_, _11587_, _11585_);
  nor (_11589_, _11557_, \oc8051_golden_model_1.PC [9]);
  nor (_11590_, _11589_, _11558_);
  and (_11591_, _11590_, _03463_);
  nor (_11592_, _11590_, _03463_);
  nor (_11593_, _11592_, _11591_);
  and (_11594_, _06059_, _03463_);
  nor (_11595_, _06059_, _03463_);
  and (_11596_, _05915_, _03207_);
  nor (_11597_, _11596_, \oc8051_golden_model_1.PC [6]);
  nor (_11598_, _11597_, _06056_);
  not (_11599_, _11598_);
  nor (_11600_, _11599_, _03556_);
  and (_11601_, _11599_, _03556_);
  nor (_11602_, _11601_, _11600_);
  not (_11603_, _11602_);
  and (_11604_, _03207_, \oc8051_golden_model_1.PC [4]);
  nor (_11605_, _11604_, \oc8051_golden_model_1.PC [5]);
  nor (_11606_, _11605_, _11596_);
  not (_11607_, _11606_);
  nor (_11608_, _11607_, _03853_);
  and (_11609_, _11607_, _03853_);
  nor (_11610_, _03207_, \oc8051_golden_model_1.PC [4]);
  nor (_11611_, _11610_, _11604_);
  not (_11612_, _11611_);
  nor (_11613_, _11612_, _04308_);
  nor (_11614_, _03494_, _03211_);
  and (_11615_, _03494_, _03211_);
  nor (_11616_, _03898_, _03362_);
  nor (_11617_, _04434_, \oc8051_golden_model_1.PC [1]);
  nor (_11618_, _04042_, _02938_);
  and (_11619_, _04434_, \oc8051_golden_model_1.PC [1]);
  nor (_11620_, _11619_, _11617_);
  and (_11621_, _11620_, _11618_);
  nor (_11622_, _11621_, _11617_);
  and (_11623_, _03898_, _03362_);
  nor (_11624_, _11623_, _11616_);
  not (_11625_, _11624_);
  nor (_11626_, _11625_, _11622_);
  nor (_11627_, _11626_, _11616_);
  nor (_11628_, _11627_, _11615_);
  nor (_11629_, _11628_, _11614_);
  and (_11630_, _11612_, _04308_);
  nor (_11631_, _11630_, _11613_);
  not (_11632_, _11631_);
  nor (_11633_, _11632_, _11629_);
  nor (_11634_, _11633_, _11613_);
  nor (_11635_, _11634_, _11609_);
  nor (_11636_, _11635_, _11608_);
  nor (_11637_, _11636_, _11603_);
  nor (_11638_, _11637_, _11600_);
  nor (_11639_, _11638_, _11595_);
  or (_11640_, _11639_, _11594_);
  nor (_11641_, _06057_, \oc8051_golden_model_1.PC [8]);
  nor (_11642_, _11641_, _11557_);
  and (_11643_, _11642_, _03463_);
  nor (_11644_, _11642_, _03463_);
  nor (_11645_, _11644_, _11643_);
  and (_11646_, _11645_, _11640_);
  and (_11647_, _11646_, _11593_);
  and (_11648_, _11647_, _11588_);
  nor (_11649_, _11643_, _11591_);
  not (_11650_, _11649_);
  and (_11651_, _11650_, _11588_);
  or (_11652_, _11651_, _11583_);
  nor (_11653_, _11652_, _11648_);
  and (_11654_, _11653_, _11580_);
  not (_11655_, _11654_);
  nor (_11656_, _11575_, _03463_);
  nor (_11657_, _11656_, _11576_);
  and (_11658_, _11657_, _11655_);
  nor (_11659_, _11658_, _11576_);
  nor (_11660_, _11659_, _11573_);
  nor (_11661_, _11660_, _11572_);
  nor (_11662_, _11661_, _11569_);
  nor (_11663_, _11662_, _11566_);
  nor (_11664_, _06874_, _03463_);
  and (_11665_, _06874_, _03463_);
  nor (_11666_, _11665_, _11664_);
  and (_11667_, _11666_, _11663_);
  nor (_11668_, _11666_, _11663_);
  or (_11669_, _11668_, _11667_);
  and (_11670_, _11669_, _11556_);
  or (_11671_, _11670_, _11555_);
  or (_11672_, _11671_, _06054_);
  and (_11673_, _11672_, _11550_);
  nor (_11674_, _04509_, _03599_);
  not (_11675_, _11674_);
  or (_11676_, _11675_, _11673_);
  and (_11677_, _11676_, _11529_);
  or (_11678_, _11677_, _11392_);
  and (_11679_, _03604_, _03257_);
  and (_11680_, _11391_, _06068_);
  or (_11681_, _11680_, _11352_);
  and (_11682_, _11681_, _11679_);
  and (_11683_, _11682_, _11678_);
  and (_11684_, _08041_, _08102_);
  or (_11685_, _11679_, _06875_);
  nand (_11686_, _11685_, _11684_);
  or (_11687_, _11686_, _11683_);
  or (_11688_, _11684_, _11352_);
  and (_11689_, _11688_, _03611_);
  and (_11690_, _11689_, _11687_);
  or (_11691_, _11690_, _11390_);
  nor (_11692_, _09979_, _08106_);
  and (_11693_, _11692_, _11691_);
  not (_11694_, _11692_);
  and (_11695_, _11694_, _11352_);
  not (_11696_, _03260_);
  nor (_11697_, _03510_, _11696_);
  and (_11698_, _11697_, _03512_);
  not (_11699_, _11698_);
  or (_11700_, _11699_, _11695_);
  or (_11701_, _11700_, _11693_);
  or (_11702_, _11698_, _06874_);
  and (_11703_, _11702_, _09988_);
  and (_11704_, _11703_, _11701_);
  nand (_11705_, _10037_, _11377_);
  not (_11706_, _09988_);
  or (_11707_, _11524_, _10037_);
  and (_11708_, _11707_, _11706_);
  and (_11709_, _11708_, _11705_);
  or (_11710_, _11709_, _10041_);
  or (_11711_, _11710_, _11704_);
  and (_11712_, _11711_, _04046_);
  not (_11713_, _10089_);
  and (_11714_, _11524_, _11713_);
  and (_11715_, _10089_, _06867_);
  or (_11716_, _11715_, _10042_);
  or (_11717_, _11716_, _11714_);
  and (_11718_, _11717_, _11712_);
  not (_11719_, _09946_);
  and (_11720_, _11524_, _11719_);
  and (_11721_, _09946_, _06867_);
  or (_11722_, _11721_, _11720_);
  and (_11723_, _11722_, _03615_);
  or (_11724_, _11723_, _11718_);
  and (_11725_, _11724_, _09916_);
  or (_11726_, _11524_, _10133_);
  nand (_11727_, _10133_, _11377_);
  and (_11728_, _11727_, _03676_);
  and (_11729_, _11728_, _11726_);
  or (_11730_, _11729_, _11725_);
  and (_11731_, _11730_, _11389_);
  nand (_11732_, _11352_, _10096_);
  and (_11733_, _04999_, _03622_);
  and (_11734_, _11733_, _03593_);
  nand (_11735_, _11734_, _11732_);
  or (_11736_, _11735_, _11731_);
  or (_11737_, _11734_, _06874_);
  and (_11738_, _11737_, _11386_);
  and (_11739_, _11738_, _11736_);
  or (_11740_, _11739_, _11388_);
  and (_11741_, _03631_, _03265_);
  and (_11742_, _11741_, _11740_);
  or (_11743_, _11741_, _06875_);
  nand (_11744_, _11743_, _11381_);
  or (_11745_, _11744_, _11742_);
  and (_11746_, _11745_, _11382_);
  or (_11747_, _11746_, _11380_);
  or (_11748_, _11379_, _06874_);
  and (_11749_, _11748_, _03285_);
  and (_11750_, _11749_, _11747_);
  and (_11751_, _11352_, _03371_);
  nor (_11752_, _03500_, _03497_);
  not (_11753_, _11752_);
  or (_11754_, _11753_, _11751_);
  or (_11755_, _11754_, _11750_);
  or (_11756_, _11752_, _06874_);
  and (_11757_, _11756_, _08865_);
  and (_11758_, _11757_, _11755_);
  and (_11759_, _06889_, _05970_);
  nand (_11760_, _06867_, _03656_);
  nand (_11761_, _11760_, _11759_);
  or (_11762_, _11761_, _11758_);
  or (_11763_, _11759_, _06874_);
  and (_11764_, _11763_, _03275_);
  and (_11765_, _11764_, _11762_);
  or (_11766_, _11765_, _11378_);
  nor (_11767_, _07455_, _03313_);
  and (_11768_, _11767_, _11766_);
  not (_11769_, _11374_);
  not (_11770_, _11767_);
  and (_11771_, _11770_, _11352_);
  or (_11772_, _11771_, _11769_);
  or (_11773_, _11772_, _11768_);
  and (_11774_, _11773_, _11376_);
  and (_11775_, _11669_, _11372_);
  or (_11776_, _11775_, _06246_);
  or (_11777_, _11776_, _11774_);
  or (_11778_, _06874_, _05966_);
  and (_11779_, _11778_, _04582_);
  and (_11780_, _11779_, _11777_);
  and (_11781_, _06867_, _03650_);
  or (_11782_, _11781_, _08445_);
  or (_11783_, _11782_, _11780_);
  and (_11784_, _03648_, _03226_);
  not (_11785_, _11784_);
  nand (_11786_, _08445_, _06875_);
  and (_11787_, _11786_, _11785_);
  and (_11788_, _11787_, _11783_);
  and (_11789_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_11790_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_11791_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_11792_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_11793_, _11792_, _11791_);
  not (_11794_, _11793_);
  and (_11795_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_11796_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_11797_, _11796_, _11795_);
  not (_11798_, _11797_);
  and (_11799_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_11800_, _03302_, _03298_);
  nor (_11801_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_11802_, _11801_, _11799_);
  not (_11803_, _11802_);
  nor (_11804_, _11803_, _11800_);
  nor (_11805_, _11804_, _11799_);
  nor (_11806_, _11805_, _11798_);
  nor (_11807_, _11806_, _11795_);
  nor (_11808_, _11807_, _11794_);
  nor (_11809_, _11808_, _11791_);
  nor (_11810_, _11809_, _11790_);
  or (_11811_, _11810_, _11789_);
  and (_11812_, _11811_, _08984_);
  and (_11813_, _11812_, \oc8051_golden_model_1.DPH [2]);
  and (_11814_, _11813_, \oc8051_golden_model_1.DPH [3]);
  and (_11815_, _11814_, \oc8051_golden_model_1.DPH [4]);
  and (_11816_, _11815_, \oc8051_golden_model_1.DPH [5]);
  and (_11817_, _11816_, \oc8051_golden_model_1.DPH [6]);
  nand (_11818_, _11817_, \oc8051_golden_model_1.DPH [7]);
  or (_11819_, _11817_, \oc8051_golden_model_1.DPH [7]);
  and (_11820_, _11819_, _11784_);
  and (_11821_, _11820_, _11818_);
  nor (_11822_, _03561_, _03227_);
  not (_11823_, _11822_);
  or (_11824_, _11823_, _11821_);
  or (_11825_, _11824_, _11788_);
  and (_11826_, _03226_, _03204_);
  not (_11827_, _11826_);
  or (_11828_, _11822_, _06874_);
  and (_11829_, _11828_, _11827_);
  and (_11830_, _11829_, _11825_);
  or (_11831_, _11669_, _08820_);
  not (_11832_, _08820_);
  or (_11833_, _11832_, _06874_);
  and (_11834_, _11833_, _11826_);
  and (_11835_, _11834_, _11831_);
  or (_11836_, _11835_, _11830_);
  nor (_11837_, _04839_, _08453_);
  nor (_11838_, _11837_, _08451_);
  and (_11839_, _03666_, _03230_);
  nor (_11840_, _11839_, _07952_);
  and (_11841_, _11840_, _11838_);
  and (_11842_, _11841_, _11836_);
  nor (_11843_, _08472_, _03776_);
  not (_11844_, _11843_);
  not (_11845_, _11841_);
  and (_11846_, _11845_, _11352_);
  or (_11847_, _11846_, _11844_);
  or (_11848_, _11847_, _11842_);
  or (_11849_, _11843_, _06874_);
  and (_11850_, _11849_, _04591_);
  and (_11851_, _11850_, _11848_);
  nand (_11852_, _06867_, _03649_);
  nor (_11853_, _03778_, _03231_);
  nand (_11854_, _11853_, _11852_);
  or (_11855_, _11854_, _11851_);
  and (_11856_, _03230_, _03204_);
  not (_11857_, _11856_);
  or (_11858_, _11853_, _06874_);
  and (_11859_, _11858_, _11857_);
  and (_11860_, _11859_, _11855_);
  or (_11861_, _11669_, _11832_);
  or (_11862_, _08820_, _06874_);
  and (_11863_, _11862_, _11856_);
  and (_11864_, _11863_, _11861_);
  not (_11865_, _11370_);
  or (_11866_, _11865_, _11864_);
  or (_11867_, _11866_, _11860_);
  and (_11868_, _11867_, _11371_);
  or (_11869_, _11868_, _11368_);
  or (_11870_, _11367_, _06874_);
  and (_11871_, _11870_, _04596_);
  and (_11872_, _11871_, _11869_);
  nand (_11873_, _06867_, _03655_);
  nand (_11874_, _11873_, _10776_);
  or (_11875_, _11874_, _11872_);
  and (_11876_, _11875_, _11366_);
  not (_11877_, _11361_);
  or (_11878_, _11669_, \oc8051_golden_model_1.PSW [7]);
  or (_11879_, _06874_, _07911_);
  and (_11880_, _11879_, _11363_);
  and (_11881_, _11880_, _11878_);
  or (_11882_, _11881_, _11877_);
  or (_11883_, _11882_, _11876_);
  and (_11884_, _11883_, _11362_);
  or (_11885_, _11884_, _11358_);
  or (_11886_, _11357_, _06874_);
  and (_11887_, _11886_, _04608_);
  and (_11888_, _11887_, _11885_);
  nand (_11889_, _06867_, _03653_);
  nor (_11890_, _03786_, _03236_);
  nand (_11891_, _11890_, _11889_);
  or (_11892_, _11891_, _11888_);
  and (_11893_, _03235_, _03204_);
  not (_11894_, _11893_);
  or (_11895_, _11890_, _06874_);
  and (_11896_, _11895_, _11894_);
  and (_11897_, _11896_, _11892_);
  not (_11898_, _11355_);
  or (_11899_, _11669_, _07911_);
  or (_11900_, _06874_, \oc8051_golden_model_1.PSW [7]);
  and (_11901_, _11900_, _11893_);
  and (_11902_, _11901_, _11899_);
  or (_11903_, _11902_, _11898_);
  or (_11904_, _11903_, _11897_);
  and (_11905_, _11904_, _11356_);
  or (_11906_, _11905_, _08571_);
  or (_11907_, _08570_, _06874_);
  and (_11908_, _11907_, _08601_);
  and (_11909_, _11908_, _11906_);
  and (_11910_, _11352_, _08600_);
  or (_11911_, _11910_, _03792_);
  or (_11912_, _11911_, _11909_);
  nand (_11913_, _05289_, _03792_);
  and (_11914_, _11913_, _11912_);
  or (_11915_, _11914_, _03248_);
  nand (_11916_, _06875_, _03248_);
  and (_11917_, _11916_, _03796_);
  and (_11918_, _11917_, _11915_);
  not (_11919_, _11353_);
  not (_11920_, _09914_);
  or (_11921_, _11524_, _11920_);
  or (_11922_, _09914_, _06867_);
  and (_11923_, _11922_, _03652_);
  and (_11924_, _11923_, _11921_);
  or (_11925_, _11924_, _11919_);
  or (_11926_, _11925_, _11918_);
  and (_11927_, _11926_, _11354_);
  or (_11928_, _11927_, _08722_);
  or (_11929_, _08721_, _06874_);
  and (_11930_, _11929_, _08770_);
  and (_11931_, _11930_, _11928_);
  and (_11932_, _11352_, _08769_);
  or (_11933_, _11932_, _03521_);
  or (_11934_, _11933_, _11931_);
  nand (_11935_, _05289_, _03521_);
  and (_11936_, _11935_, _11934_);
  or (_11937_, _11936_, _03246_);
  nand (_11938_, _06875_, _03246_);
  and (_11939_, _11938_, _03520_);
  and (_11940_, _11939_, _11937_);
  or (_11941_, _11524_, _09914_);
  nand (_11942_, _09914_, _11377_);
  and (_11943_, _11942_, _11941_);
  and (_11944_, _11943_, _03519_);
  and (_11945_, _06814_, _06486_);
  not (_11946_, _11945_);
  or (_11947_, _11946_, _11944_);
  or (_11948_, _11947_, _11940_);
  or (_11949_, _11945_, _11352_);
  and (_11950_, _11949_, _04260_);
  and (_11951_, _11950_, _11948_);
  nor (_11952_, _08814_, _08809_);
  nand (_11953_, _06874_, _03809_);
  nand (_11954_, _11953_, _11952_);
  or (_11955_, _11954_, _11951_);
  not (_11956_, _03686_);
  or (_11957_, _11352_, _11952_);
  and (_11958_, _11957_, _11956_);
  and (_11959_, _11958_, _11955_);
  and (_11960_, _03686_, _03463_);
  or (_11961_, _11960_, _03243_);
  or (_11962_, _11961_, _11959_);
  nand (_11963_, _06875_, _03243_);
  and (_11964_, _11963_, _03206_);
  and (_11965_, _11964_, _11962_);
  and (_11966_, _11943_, _03205_);
  and (_11967_, _05913_, _06833_);
  not (_11968_, _11967_);
  or (_11969_, _11968_, _11966_);
  or (_11970_, _11969_, _11965_);
  or (_11971_, _11967_, _11352_);
  and (_11972_, _11971_, _03820_);
  and (_11973_, _11972_, _11970_);
  nor (_11974_, _08838_, _08831_);
  nand (_11975_, _06874_, _03816_);
  nand (_11976_, _11975_, _11974_);
  or (_11977_, _11976_, _11973_);
  not (_11978_, _03684_);
  or (_11979_, _11352_, _11974_);
  and (_11980_, _11979_, _11978_);
  and (_11981_, _11980_, _11977_);
  and (_11982_, _03241_, _03204_);
  nor (_11983_, _03684_, _03242_);
  not (_11984_, _11983_);
  or (_11985_, _03463_, _03242_);
  and (_11986_, _11985_, _11984_);
  or (_11987_, _11986_, _11982_);
  or (_11988_, _11987_, _11981_);
  nand (_11989_, _06875_, _03242_);
  not (_11990_, _11982_);
  or (_11991_, _11990_, _11352_);
  and (_11992_, _11991_, _11989_);
  and (_11993_, _11992_, _11988_);
  or (_11994_, _11993_, _43231_);
  or (_11995_, _43227_, \oc8051_golden_model_1.PC [15]);
  and (_11996_, _11995_, _41991_);
  and (_40770_, _11996_, _11994_);
  and (_11997_, _43231_, \oc8051_golden_model_1.P0INREG [7]);
  or (_11998_, _11997_, _01119_);
  and (_40771_, _11998_, _41991_);
  and (_11999_, _43231_, \oc8051_golden_model_1.P1INREG [7]);
  or (_12000_, _11999_, _00968_);
  and (_40772_, _12000_, _41991_);
  and (_12001_, _43231_, \oc8051_golden_model_1.P2INREG [7]);
  or (_12002_, _12001_, _01179_);
  and (_40774_, _12002_, _41991_);
  and (_12003_, _43231_, \oc8051_golden_model_1.P3INREG [7]);
  or (_12004_, _12003_, _01028_);
  and (_40775_, _12004_, _41991_);
  nor (_12005_, _04892_, _04638_);
  nor (_12006_, _12005_, _04893_);
  nor (_12007_, _05065_, _04892_);
  nor (_12008_, _12007_, _05206_);
  and (_12009_, _12008_, _04891_);
  and (_12010_, _12009_, _12006_);
  not (_12011_, _12010_);
  or (_12012_, _04510_, _04271_);
  and (_12013_, _12012_, _11968_);
  nand (_12014_, _03243_, _02938_);
  nor (_12015_, _05744_, \oc8051_golden_model_1.ACC [0]);
  nand (_12016_, _12015_, _04607_);
  nor (_12017_, _05744_, _06366_);
  and (_12018_, _05744_, _06366_);
  nor (_12019_, _12018_, _12017_);
  and (_12020_, _12019_, _04592_);
  or (_12021_, _04568_, _04491_);
  nand (_12022_, _08238_, _03594_);
  nor (_12023_, _10193_, _05332_);
  or (_12024_, _12023_, _06028_);
  nor (_12025_, _05744_, _06175_);
  or (_12026_, _06054_, _04510_);
  nand (_12027_, _03947_, _02938_);
  or (_12028_, _03947_, \oc8051_golden_model_1.ACC [0]);
  nand (_12029_, _12028_, _12027_);
  and (_12030_, _12029_, _06054_);
  nor (_12031_, _12030_, _04516_);
  and (_12032_, _12031_, _12026_);
  or (_12033_, _12032_, _12025_);
  and (_12034_, _12033_, _06040_);
  nand (_12035_, _10193_, _09809_);
  and (_12036_, _12035_, _04514_);
  or (_12037_, _12036_, _04857_);
  or (_12038_, _12037_, _12034_);
  nor (_12039_, _03257_, \oc8051_golden_model_1.PC [0]);
  nor (_12040_, _12039_, _04525_);
  and (_12041_, _12040_, _12038_);
  and (_12042_, _04525_, _04491_);
  or (_12043_, _12042_, _04533_);
  or (_12044_, _12043_, _12041_);
  and (_12045_, _12044_, _12024_);
  or (_12046_, _12045_, _03510_);
  nand (_12047_, _08238_, _03510_);
  and (_12048_, _12047_, _03508_);
  and (_12049_, _12048_, _12046_);
  nor (_12050_, _10194_, _03508_);
  and (_12051_, _12050_, _12035_);
  or (_12052_, _12051_, _12049_);
  and (_12053_, _12052_, _03253_);
  or (_12054_, _03253_, _02938_);
  nand (_12055_, _03593_, _12054_);
  or (_12056_, _12055_, _12053_);
  and (_12057_, _12056_, _12022_);
  or (_12058_, _12057_, _04551_);
  and (_12059_, _06836_, _04559_);
  nand (_12060_, _08237_, _04551_);
  or (_12061_, _12060_, _12059_);
  and (_12062_, _12061_, _12058_);
  or (_12063_, _12062_, _04550_);
  nor (_12064_, _09832_, _05332_);
  and (_12065_, _05332_, \oc8051_golden_model_1.PSW [7]);
  nor (_12066_, _12065_, _12064_);
  nand (_12067_, _12066_, _04550_);
  and (_12068_, _12067_, _03278_);
  and (_12069_, _12068_, _12063_);
  or (_12070_, _03278_, _02938_);
  nand (_12071_, _04568_, _12070_);
  or (_12072_, _12071_, _12069_);
  and (_12073_, _12072_, _12021_);
  or (_12074_, _12073_, _05971_);
  and (_12075_, _06836_, _06242_);
  or (_12076_, _12075_, _04571_);
  and (_12077_, _12076_, _12074_);
  and (_12078_, _05958_, _04491_);
  and (_12079_, _06427_, \oc8051_golden_model_1.PSW [0]);
  not (_12080_, _12079_);
  and (_12081_, _06388_, _06381_);
  and (_12082_, _12081_, \oc8051_golden_model_1.IP [0]);
  not (_12083_, _12082_);
  and (_12084_, _06432_, \oc8051_golden_model_1.ACC [0]);
  and (_12085_, _06380_, _06355_);
  and (_12086_, _06425_, _12085_);
  and (_12087_, _12086_, \oc8051_golden_model_1.B [0]);
  nor (_12088_, _12087_, _12084_);
  and (_12089_, _12088_, _12083_);
  and (_12090_, _12089_, _12080_);
  and (_12091_, _06368_, \oc8051_golden_model_1.SP [0]);
  not (_12092_, _12091_);
  and (_12093_, _06422_, \oc8051_golden_model_1.DPL [0]);
  and (_12094_, _06356_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_12095_, _12094_, _12093_);
  and (_12096_, _12095_, _12092_);
  and (_12097_, _12096_, _12090_);
  and (_12098_, _06389_, \oc8051_golden_model_1.IE [0]);
  not (_12099_, _12098_);
  and (_12100_, _06392_, \oc8051_golden_model_1.SCON [0]);
  and (_12101_, _06394_, \oc8051_golden_model_1.SBUF [0]);
  nor (_12102_, _12101_, _12100_);
  and (_12103_, _12102_, _12099_);
  and (_12104_, _06382_, \oc8051_golden_model_1.P3INREG [0]);
  and (_12105_, _06361_, \oc8051_golden_model_1.P2INREG [0]);
  and (_12106_, _06378_, \oc8051_golden_model_1.P1INREG [0]);
  or (_12107_, _12106_, _12105_);
  nor (_12108_, _12107_, _12104_);
  and (_12109_, _12108_, _12103_);
  and (_12110_, _06409_, \oc8051_golden_model_1.TH0 [0]);
  and (_12111_, _06411_, \oc8051_golden_model_1.TL1 [0]);
  nor (_12112_, _12111_, _12110_);
  and (_12113_, _06416_, \oc8051_golden_model_1.PCON [0]);
  and (_12114_, _06418_, \oc8051_golden_model_1.TCON [0]);
  nor (_12115_, _12114_, _12113_);
  and (_12116_, _12115_, _12112_);
  and (_12117_, _06400_, \oc8051_golden_model_1.DPH [0]);
  and (_12118_, _06367_, _06349_);
  and (_12119_, _12118_, \oc8051_golden_model_1.TMOD [0]);
  nor (_12120_, _12119_, _12117_);
  and (_12121_, _06404_, \oc8051_golden_model_1.TH1 [0]);
  and (_12122_, _06350_, \oc8051_golden_model_1.TL0 [0]);
  nor (_12123_, _12122_, _12121_);
  and (_12124_, _12123_, _12120_);
  and (_12125_, _12124_, _12116_);
  and (_12126_, _12125_, _12109_);
  and (_12127_, _12126_, _12097_);
  not (_12128_, _12127_);
  nor (_12129_, _12128_, _12078_);
  nor (_12130_, _12129_, _06242_);
  or (_12131_, _12130_, _06246_);
  or (_12132_, _12131_, _12077_);
  and (_12133_, _06246_, _04042_);
  nor (_12134_, _12133_, _04583_);
  and (_12135_, _12134_, _12132_);
  and (_12136_, _04583_, _06366_);
  or (_12137_, _12136_, _03227_);
  or (_12138_, _12137_, _12135_);
  and (_12139_, _03227_, _02938_);
  nor (_12140_, _12139_, _04592_);
  and (_12141_, _12140_, _12138_);
  or (_12142_, _12141_, _12020_);
  and (_12143_, _12142_, _05927_);
  and (_12144_, _05744_, \oc8051_golden_model_1.ACC [0]);
  nor (_12145_, _12144_, _12015_);
  and (_12146_, _12145_, _04590_);
  or (_12147_, _12146_, _12143_);
  and (_12148_, _12147_, _05926_);
  and (_12149_, _12018_, _04597_);
  or (_12150_, _12149_, _04595_);
  or (_12151_, _12150_, _12148_);
  or (_12152_, _12144_, _05925_);
  and (_12153_, _12152_, _12151_);
  or (_12154_, _12153_, _03238_);
  and (_12155_, _03238_, _02938_);
  nor (_12156_, _12155_, _04609_);
  and (_12157_, _12156_, _12154_);
  nor (_12158_, _12017_, _06471_);
  or (_12159_, _12158_, _04607_);
  or (_12160_, _12159_, _12157_);
  and (_12161_, _12160_, _12016_);
  or (_12162_, _12161_, _03248_);
  nand (_12163_, _03248_, _02938_);
  and (_12164_, _12163_, _06814_);
  and (_12165_, _12164_, _12162_);
  nor (_12166_, _06814_, _04491_);
  or (_12167_, _12166_, _12165_);
  and (_12168_, _12167_, _06486_);
  and (_12169_, _06622_, _04618_);
  or (_12170_, _12169_, _04617_);
  or (_12171_, _12170_, _12168_);
  nand (_12172_, _05744_, _04617_);
  and (_12173_, _12172_, _11956_);
  and (_12174_, _12173_, _12171_);
  and (_12175_, _03686_, _02938_);
  or (_12176_, _12175_, _03243_);
  or (_12177_, _12176_, _12174_);
  and (_12178_, _12177_, _12014_);
  or (_12179_, _12178_, _04624_);
  not (_12180_, _04624_);
  or (_12181_, _12064_, _12180_);
  and (_12182_, _12181_, _05913_);
  and (_12183_, _12182_, _12179_);
  or (_12184_, _12183_, _12013_);
  or (_12185_, _06622_, _06833_);
  and (_12186_, _12185_, _12184_);
  nor (_12187_, _12186_, _04633_);
  and (_12188_, _05744_, _04633_);
  or (_12189_, _12188_, _04892_);
  nor (_12190_, _12189_, _12187_);
  or (_12191_, _12190_, _12011_);
  nor (_12192_, _05228_, _04800_);
  nor (_12193_, _12192_, _05229_);
  nor (_12194_, _05228_, _05205_);
  nor (_12195_, _12194_, _05233_);
  and (_12196_, _12195_, _05227_);
  and (_12197_, _12196_, _12193_);
  or (_12198_, _12197_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_12199_, _05220_, _04801_);
  nor (_12200_, _05213_, _05216_);
  and (_12201_, _12200_, _12199_);
  and (_12202_, _12201_, _04645_);
  not (_12203_, _12202_);
  and (_12204_, _12203_, _12198_);
  and (_12205_, _12204_, _12191_);
  not (_12206_, _11642_);
  nor (_12207_, _12206_, _03686_);
  and (_12208_, _11496_, _03686_);
  or (_12209_, _12208_, _12207_);
  and (_12210_, _12209_, _12202_);
  or (_40790_, _12210_, _12205_);
  or (_12211_, _12197_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_12212_, _12211_, _12203_);
  not (_12213_, _12197_);
  nor (_12214_, _06045_, _05899_);
  and (_12215_, _12214_, _06827_);
  not (_12216_, _06481_);
  and (_12217_, _03248_, _02911_);
  and (_12218_, _05698_, _04347_);
  nor (_12219_, _05698_, _04347_);
  nor (_12220_, _12219_, _12218_);
  and (_12221_, _12220_, _04592_);
  or (_12222_, _05898_, _04568_);
  nand (_12223_, _08223_, _03594_);
  nor (_12224_, _10167_, _05314_);
  or (_12225_, _12224_, _06028_);
  not (_12226_, _06054_);
  nand (_12227_, _12214_, _12226_);
  nor (_12228_, _03947_, _03320_);
  and (_12229_, _03947_, _02911_);
  nor (_12230_, _12229_, _12228_);
  nand (_12231_, _12230_, _06054_);
  and (_12232_, _12231_, _12227_);
  and (_12233_, _12232_, _06175_);
  nor (_12234_, _06178_, _05745_);
  nor (_12235_, _12234_, _06175_);
  or (_12236_, _12235_, _12233_);
  or (_12237_, _12236_, _04514_);
  nand (_12238_, _10167_, _09755_);
  or (_12239_, _12238_, _06040_);
  and (_12240_, _12239_, _12237_);
  or (_12241_, _12240_, _04857_);
  nor (_12242_, _03257_, _02911_);
  nor (_12243_, _12242_, _04525_);
  and (_12244_, _12243_, _12241_);
  and (_12245_, _05898_, _04525_);
  or (_12246_, _12245_, _04533_);
  or (_12247_, _12246_, _12244_);
  and (_12248_, _12247_, _12225_);
  or (_12249_, _12248_, _03510_);
  nand (_12250_, _08223_, _03510_);
  and (_12251_, _12250_, _03508_);
  and (_12252_, _12251_, _12249_);
  not (_12253_, _10168_);
  and (_12254_, _12238_, _12253_);
  and (_12255_, _12254_, _03507_);
  or (_12256_, _12255_, _12252_);
  and (_12257_, _12256_, _03253_);
  or (_12258_, _03253_, \oc8051_golden_model_1.PC [1]);
  nand (_12259_, _03593_, _12258_);
  or (_12260_, _12259_, _12257_);
  and (_12261_, _12260_, _12223_);
  or (_12262_, _12261_, _04551_);
  and (_12263_, _06835_, _04559_);
  nand (_12264_, _08222_, _04551_);
  or (_12265_, _12264_, _12263_);
  and (_12266_, _12265_, _12262_);
  or (_12267_, _12266_, _04550_);
  nor (_12268_, _09778_, _05314_);
  and (_12269_, _05314_, \oc8051_golden_model_1.PSW [7]);
  nor (_12270_, _12269_, _12268_);
  nand (_12271_, _12270_, _04550_);
  and (_12272_, _12271_, _03278_);
  and (_12273_, _12272_, _12267_);
  or (_12274_, _03278_, \oc8051_golden_model_1.PC [1]);
  nand (_12275_, _04568_, _12274_);
  or (_12276_, _12275_, _12273_);
  and (_12277_, _12276_, _12222_);
  or (_12278_, _12277_, _05971_);
  and (_12279_, _06835_, _06242_);
  or (_12280_, _12279_, _04571_);
  and (_12281_, _12280_, _12278_);
  and (_12282_, _05958_, _05898_);
  and (_12283_, _06350_, \oc8051_golden_model_1.TL0 [1]);
  not (_12284_, _12283_);
  and (_12285_, _06356_, \oc8051_golden_model_1.P0INREG [1]);
  and (_12286_, _06361_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_12287_, _12286_, _12285_);
  and (_12288_, _12287_, _12284_);
  and (_12289_, _06368_, \oc8051_golden_model_1.SP [1]);
  not (_12290_, _12289_);
  and (_12291_, _06372_, \oc8051_golden_model_1.TMOD [1]);
  not (_12292_, _12291_);
  and (_12293_, _06378_, \oc8051_golden_model_1.P1INREG [1]);
  and (_12294_, _06382_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_12295_, _12294_, _12293_);
  and (_12296_, _12295_, _12292_);
  and (_12297_, _12296_, _12290_);
  and (_12298_, _12297_, _12288_);
  and (_12299_, _06389_, \oc8051_golden_model_1.IE [1]);
  not (_12300_, _12299_);
  and (_12301_, _06392_, \oc8051_golden_model_1.SCON [1]);
  and (_12302_, _06394_, \oc8051_golden_model_1.SBUF [1]);
  nor (_12303_, _12302_, _12301_);
  and (_12304_, _12303_, _12300_);
  and (_12305_, _06400_, \oc8051_golden_model_1.DPH [1]);
  and (_12306_, _06404_, \oc8051_golden_model_1.TH1 [1]);
  nor (_12307_, _12306_, _12305_);
  and (_12308_, _12307_, _12304_);
  and (_12309_, _12308_, _12298_);
  and (_12310_, _06409_, \oc8051_golden_model_1.TH0 [1]);
  and (_12311_, _06411_, \oc8051_golden_model_1.TL1 [1]);
  nor (_12312_, _12311_, _12310_);
  and (_12313_, _06416_, \oc8051_golden_model_1.PCON [1]);
  and (_12314_, _06418_, \oc8051_golden_model_1.TCON [1]);
  nor (_12315_, _12314_, _12313_);
  and (_12316_, _12315_, _12312_);
  and (_12317_, _06422_, \oc8051_golden_model_1.DPL [1]);
  not (_12318_, _12317_);
  and (_12319_, _06429_, \oc8051_golden_model_1.B [1]);
  and (_12320_, _06435_, \oc8051_golden_model_1.IP [1]);
  nor (_12321_, _12320_, _12319_);
  and (_12322_, _06427_, \oc8051_golden_model_1.PSW [1]);
  and (_12323_, _06432_, \oc8051_golden_model_1.ACC [1]);
  nor (_12324_, _12323_, _12322_);
  and (_12325_, _12324_, _12321_);
  and (_12326_, _12325_, _12318_);
  and (_12327_, _12326_, _12316_);
  and (_12328_, _12327_, _12309_);
  not (_12329_, _12328_);
  nor (_12330_, _12329_, _12282_);
  nor (_12331_, _12330_, _06242_);
  or (_12332_, _12331_, _06246_);
  or (_12333_, _12332_, _12281_);
  and (_12334_, _06246_, _04434_);
  nor (_12335_, _12334_, _04583_);
  and (_12336_, _12335_, _12333_);
  and (_12337_, _04583_, _06249_);
  or (_12338_, _12337_, _03227_);
  or (_12339_, _12338_, _12336_);
  and (_12340_, _03227_, \oc8051_golden_model_1.PC [1]);
  nor (_12341_, _12340_, _04592_);
  and (_12342_, _12341_, _12339_);
  or (_12343_, _12342_, _12221_);
  and (_12344_, _12343_, _05927_);
  nor (_12345_, _05698_, _03320_);
  and (_12346_, _05698_, _03320_);
  nor (_12347_, _12346_, _12345_);
  and (_12348_, _12347_, _04590_);
  or (_12349_, _12348_, _12344_);
  and (_12350_, _12349_, _05926_);
  and (_12351_, _12219_, _04597_);
  or (_12352_, _12351_, _04595_);
  or (_12353_, _12352_, _12350_);
  or (_12354_, _12345_, _05925_);
  and (_12355_, _12354_, _12353_);
  or (_12356_, _12355_, _03238_);
  and (_12357_, _03238_, \oc8051_golden_model_1.PC [1]);
  nor (_12358_, _12357_, _04609_);
  and (_12359_, _12358_, _12356_);
  nor (_12360_, _12218_, _06471_);
  or (_12361_, _12360_, _04607_);
  or (_12362_, _12361_, _12359_);
  nand (_12363_, _12346_, _04607_);
  and (_12364_, _12363_, _06475_);
  and (_12365_, _12364_, _12362_);
  or (_12366_, _12365_, _12217_);
  and (_12367_, _12366_, _12216_);
  nor (_12368_, _12214_, _12216_);
  or (_12369_, _12368_, _04781_);
  or (_12370_, _12369_, _12367_);
  nand (_12371_, _12214_, _04781_);
  and (_12372_, _12371_, _06486_);
  and (_12373_, _12372_, _12370_);
  or (_12374_, _06837_, _06623_);
  and (_12375_, _12374_, _04618_);
  or (_12376_, _12375_, _04617_);
  or (_12377_, _12376_, _12373_);
  nand (_12378_, _12234_, _04617_);
  and (_12379_, _12378_, _12377_);
  or (_12380_, _12379_, _03686_);
  not (_12381_, _03243_);
  nand (_12382_, _03686_, _11470_);
  and (_12383_, _12382_, _12381_);
  and (_12384_, _12383_, _12380_);
  and (_12385_, _03243_, _02911_);
  or (_12386_, _04624_, _12385_);
  or (_12387_, _12386_, _12384_);
  or (_12388_, _12268_, _12180_);
  and (_12389_, _12388_, _05913_);
  and (_12390_, _12389_, _12387_);
  or (_12391_, _12390_, _12215_);
  and (_12392_, _12391_, _06833_);
  nor (_12393_, _06837_, _06623_);
  and (_12394_, _12393_, _04271_);
  or (_12395_, _12394_, _04633_);
  or (_12396_, _12395_, _12392_);
  or (_12397_, _12234_, _04805_);
  and (_12398_, _12397_, _05227_);
  and (_12399_, _12398_, _12396_);
  or (_12400_, _12399_, _12213_);
  and (_12401_, _12400_, _12212_);
  not (_12402_, _11590_);
  nor (_12403_, _12402_, _03686_);
  and (_12404_, _11436_, _03686_);
  or (_12405_, _12404_, _12403_);
  and (_12406_, _12405_, _12202_);
  or (_40792_, _12406_, _12401_);
  or (_12407_, _12197_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_12408_, _12407_, _12203_);
  nor (_12409_, _05899_, _07889_);
  nor (_12410_, _12409_, _07890_);
  and (_12411_, _12410_, _06827_);
  nor (_12412_, _05792_, _03943_);
  and (_12413_, _12412_, _04597_);
  nor (_12414_, _10156_, _05318_);
  or (_12415_, _12414_, _06028_);
  nand (_12416_, _10156_, _09730_);
  or (_12417_, _12416_, _06040_);
  and (_12418_, _03947_, _03356_);
  nor (_12419_, _03947_, _07634_);
  or (_12420_, _12419_, _12418_);
  and (_12421_, _12420_, _06054_);
  and (_12422_, _06045_, _05130_);
  nor (_12423_, _06045_, _05130_);
  or (_12424_, _12423_, _12422_);
  and (_12425_, _12424_, _12226_);
  or (_12426_, _12425_, _12421_);
  and (_12427_, _12426_, _06175_);
  and (_12428_, _06178_, _05792_);
  nor (_12429_, _06178_, _05792_);
  nor (_12430_, _12429_, _12428_);
  nor (_12431_, _12430_, _06175_);
  or (_12432_, _12431_, _12427_);
  or (_12433_, _12432_, _04514_);
  and (_12434_, _12433_, _12417_);
  or (_12435_, _12434_, _04857_);
  nor (_12436_, _03356_, _03257_);
  nor (_12437_, _12436_, _04525_);
  and (_12438_, _12437_, _12435_);
  and (_12439_, _07889_, _04525_);
  or (_12440_, _12439_, _04533_);
  or (_12441_, _12440_, _12438_);
  and (_12442_, _12441_, _12415_);
  or (_12443_, _12442_, _03510_);
  nand (_12444_, _08208_, _03510_);
  and (_12445_, _12444_, _03508_);
  and (_12446_, _12445_, _12443_);
  not (_12447_, _10157_);
  and (_12448_, _12416_, _12447_);
  and (_12449_, _12448_, _03507_);
  or (_12450_, _12449_, _12446_);
  and (_12451_, _12450_, _03253_);
  or (_12452_, _03362_, _03253_);
  nand (_12453_, _03593_, _12452_);
  or (_12454_, _12453_, _12451_);
  nand (_12455_, _08208_, _03594_);
  and (_12456_, _12455_, _12454_);
  or (_12457_, _12456_, _04551_);
  and (_12458_, _06839_, _04559_);
  nand (_12459_, _08207_, _04551_);
  or (_12460_, _12459_, _12458_);
  and (_12461_, _12460_, _12457_);
  or (_12462_, _12461_, _04550_);
  nor (_12463_, _09753_, _05318_);
  and (_12464_, _05318_, \oc8051_golden_model_1.PSW [7]);
  nor (_12465_, _12464_, _12463_);
  nand (_12466_, _12465_, _04550_);
  and (_12467_, _12466_, _03278_);
  and (_12468_, _12467_, _12462_);
  or (_12469_, _03362_, _03278_);
  nand (_12470_, _04568_, _12469_);
  or (_12471_, _12470_, _12468_);
  nand (_12472_, _05130_, _06238_);
  and (_12473_, _12472_, _12471_);
  or (_12474_, _12473_, _05971_);
  and (_12475_, _06839_, _06242_);
  or (_12476_, _12475_, _04571_);
  and (_12477_, _12476_, _12474_);
  nor (_12478_, _06247_, _05130_);
  and (_12479_, _06368_, \oc8051_golden_model_1.SP [2]);
  not (_12480_, _12479_);
  and (_12481_, _06350_, \oc8051_golden_model_1.TL0 [2]);
  not (_12482_, _12481_);
  and (_12483_, _06378_, \oc8051_golden_model_1.P1INREG [2]);
  and (_12484_, _06382_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_12485_, _12484_, _12483_);
  and (_12486_, _12485_, _12482_);
  and (_12487_, _06356_, \oc8051_golden_model_1.P0INREG [2]);
  and (_12488_, _06361_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_12489_, _12488_, _12487_);
  and (_12490_, _12489_, _12486_);
  and (_12491_, _12490_, _12480_);
  and (_12492_, _06389_, \oc8051_golden_model_1.IE [2]);
  not (_12493_, _12492_);
  and (_12494_, _06392_, \oc8051_golden_model_1.SCON [2]);
  and (_12495_, _06394_, \oc8051_golden_model_1.SBUF [2]);
  nor (_12496_, _12495_, _12494_);
  and (_12497_, _12496_, _12493_);
  and (_12498_, _06427_, \oc8051_golden_model_1.PSW [2]);
  and (_12499_, _06432_, \oc8051_golden_model_1.ACC [2]);
  nor (_12500_, _12499_, _12498_);
  and (_12501_, _06429_, \oc8051_golden_model_1.B [2]);
  and (_12502_, _06435_, \oc8051_golden_model_1.IP [2]);
  nor (_12503_, _12502_, _12501_);
  and (_12504_, _12503_, _12500_);
  and (_12505_, _12504_, _12497_);
  and (_12506_, _12505_, _12491_);
  and (_12507_, _06409_, \oc8051_golden_model_1.TH0 [2]);
  and (_12508_, _06411_, \oc8051_golden_model_1.TL1 [2]);
  nor (_12509_, _12508_, _12507_);
  and (_12510_, _06416_, \oc8051_golden_model_1.PCON [2]);
  and (_12511_, _06418_, \oc8051_golden_model_1.TCON [2]);
  nor (_12512_, _12511_, _12510_);
  and (_12513_, _12512_, _12509_);
  and (_12514_, _06372_, \oc8051_golden_model_1.TMOD [2]);
  and (_12515_, _06404_, \oc8051_golden_model_1.TH1 [2]);
  nor (_12516_, _12515_, _12514_);
  and (_12517_, _06422_, \oc8051_golden_model_1.DPL [2]);
  and (_12518_, _06400_, \oc8051_golden_model_1.DPH [2]);
  nor (_12519_, _12518_, _12517_);
  and (_12520_, _12519_, _12516_);
  and (_12521_, _12520_, _12513_);
  and (_12522_, _12521_, _12506_);
  not (_12523_, _12522_);
  nor (_12524_, _12523_, _12478_);
  nor (_12525_, _12524_, _06242_);
  or (_12526_, _12525_, _06246_);
  or (_12527_, _12526_, _12477_);
  and (_12528_, _06246_, _03898_);
  nor (_12529_, _12528_, _04583_);
  and (_12530_, _12529_, _12527_);
  and (_12531_, _04583_, _06414_);
  or (_12532_, _12531_, _03227_);
  or (_12533_, _12532_, _12530_);
  and (_12534_, _03362_, _03227_);
  nor (_12535_, _12534_, _04592_);
  and (_12536_, _12535_, _12533_);
  and (_12537_, _05792_, _03943_);
  nor (_12538_, _12537_, _12412_);
  and (_12539_, _12538_, _04592_);
  or (_12540_, _12539_, _04590_);
  or (_12541_, _12540_, _12536_);
  nor (_12542_, _05792_, _07634_);
  and (_12543_, _05792_, _07634_);
  nor (_12544_, _12543_, _12542_);
  or (_12545_, _12544_, _05927_);
  and (_12546_, _12545_, _05926_);
  and (_12547_, _12546_, _12541_);
  or (_12548_, _12547_, _12413_);
  and (_12549_, _12548_, _05925_);
  and (_12550_, _12542_, _04595_);
  or (_12551_, _12550_, _03238_);
  or (_12552_, _12551_, _12549_);
  and (_12553_, _03362_, _03238_);
  nor (_12554_, _12553_, _04609_);
  and (_12555_, _12554_, _12552_);
  nor (_12556_, _12537_, _06471_);
  or (_12557_, _12556_, _04607_);
  or (_12558_, _12557_, _12555_);
  nand (_12559_, _12543_, _04607_);
  and (_12560_, _12559_, _06475_);
  and (_12561_, _12560_, _12558_);
  and (_12562_, _03356_, _03248_);
  or (_12563_, _06479_, _12562_);
  or (_12564_, _12563_, _12561_);
  nor (_12565_, _06480_, _04781_);
  not (_12566_, _06479_);
  or (_12567_, _12424_, _12566_);
  and (_12568_, _12567_, _12565_);
  and (_12569_, _12568_, _12564_);
  not (_12570_, _12565_);
  and (_12571_, _12424_, _12570_);
  or (_12572_, _12571_, _04618_);
  or (_12573_, _12572_, _12569_);
  nor (_12574_, _06623_, _06714_);
  and (_12575_, _06623_, _06714_);
  or (_12576_, _12575_, _06486_);
  or (_12577_, _12576_, _12574_);
  and (_12578_, _12577_, _04811_);
  and (_12579_, _12578_, _12573_);
  nor (_12580_, _12430_, _04811_);
  or (_12581_, _12580_, _03686_);
  or (_12582_, _12581_, _12579_);
  nand (_12583_, _11468_, _03686_);
  and (_12584_, _12583_, _12381_);
  and (_12585_, _12584_, _12582_);
  and (_12586_, _03356_, _03243_);
  or (_12587_, _04624_, _12586_);
  or (_12588_, _12587_, _12585_);
  or (_12589_, _12463_, _12180_);
  and (_12590_, _12589_, _05913_);
  and (_12591_, _12590_, _12588_);
  or (_12592_, _12591_, _12411_);
  and (_12593_, _12592_, _06833_);
  or (_12594_, _06837_, _06839_);
  nor (_12595_, _07991_, _06833_);
  and (_12596_, _12595_, _12594_);
  or (_12597_, _12596_, _04633_);
  or (_12598_, _12597_, _12593_);
  nor (_12599_, _05793_, _05745_);
  nor (_12600_, _12599_, _05794_);
  or (_12601_, _12600_, _04805_);
  and (_12602_, _12601_, _05227_);
  and (_12603_, _12602_, _12598_);
  or (_12604_, _12603_, _12213_);
  and (_12605_, _12604_, _12408_);
  and (_12606_, _11422_, _03686_);
  not (_12607_, _11578_);
  nor (_12608_, _12607_, _03686_);
  or (_12609_, _12608_, _12606_);
  and (_12610_, _12609_, _12202_);
  or (_40793_, _12610_, _12605_);
  or (_12611_, _12197_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_12612_, _12611_, _12203_);
  nor (_12613_, _12575_, _06668_);
  or (_12614_, _12613_, _06716_);
  and (_12615_, _12614_, _04618_);
  and (_12616_, _03248_, _03210_);
  nor (_12617_, _05649_, _07628_);
  and (_12618_, _05649_, _07628_);
  nor (_12619_, _12618_, _12617_);
  or (_12620_, _12619_, _05927_);
  nor (_12621_, _03278_, _03211_);
  nor (_12622_, _10216_, _05296_);
  or (_12623_, _12622_, _06028_);
  nor (_12624_, _12428_, _05649_);
  nor (_12625_, _12624_, _06180_);
  nand (_12626_, _12625_, _04516_);
  nor (_12627_, _12422_, _04944_);
  or (_12628_, _12627_, _06047_);
  and (_12629_, _12628_, _12226_);
  nor (_12630_, _03947_, _07628_);
  and (_12631_, _03947_, _03210_);
  or (_12632_, _12631_, _12630_);
  and (_12633_, _12632_, _06054_);
  or (_12634_, _12633_, _04516_);
  or (_12635_, _12634_, _12629_);
  and (_12636_, _12635_, _06040_);
  and (_12637_, _12636_, _12626_);
  nand (_12638_, _10216_, _09861_);
  and (_12639_, _12638_, _04514_);
  or (_12640_, _12639_, _04857_);
  or (_12641_, _12640_, _12637_);
  nor (_12642_, _03257_, _03210_);
  nor (_12643_, _12642_, _04525_);
  and (_12644_, _12643_, _12641_);
  and (_12645_, _07888_, _04525_);
  or (_12646_, _12645_, _04533_);
  or (_12647_, _12646_, _12644_);
  and (_12648_, _12647_, _12623_);
  or (_12649_, _12648_, _03510_);
  nand (_12650_, _08191_, _03510_);
  and (_12651_, _12650_, _03508_);
  and (_12652_, _12651_, _12649_);
  not (_12653_, _10217_);
  and (_12654_, _12638_, _12653_);
  and (_12655_, _12654_, _03507_);
  or (_12656_, _12655_, _12652_);
  and (_12657_, _12656_, _03253_);
  or (_12658_, _03253_, _03211_);
  nand (_12659_, _03593_, _12658_);
  or (_12660_, _12659_, _12657_);
  nand (_12661_, _08191_, _03594_);
  and (_12662_, _12661_, _12660_);
  or (_12663_, _12662_, _04551_);
  and (_12664_, _06838_, _04559_);
  nand (_12665_, _08190_, _04551_);
  or (_12666_, _12665_, _12664_);
  and (_12667_, _12666_, _12663_);
  or (_12668_, _12667_, _04550_);
  and (_12669_, _05296_, \oc8051_golden_model_1.PSW [7]);
  nor (_12670_, _09884_, _05296_);
  nor (_12671_, _12670_, _12669_);
  nand (_12672_, _12671_, _04550_);
  and (_12673_, _12672_, _03278_);
  and (_12674_, _12673_, _12668_);
  or (_12675_, _12674_, _12621_);
  and (_12676_, _12675_, _04568_);
  nor (_12677_, _04944_, _04568_);
  or (_12678_, _12677_, _04570_);
  or (_12679_, _12678_, _12676_);
  nand (_12680_, _06668_, _05971_);
  and (_12681_, _12680_, _06242_);
  and (_12682_, _12681_, _12679_);
  nor (_12683_, _06247_, _04944_);
  and (_12684_, _06422_, \oc8051_golden_model_1.DPL [3]);
  and (_12685_, _06350_, \oc8051_golden_model_1.TL0 [3]);
  nor (_12686_, _12685_, _12684_);
  and (_12687_, _06400_, \oc8051_golden_model_1.DPH [3]);
  and (_12688_, _06404_, \oc8051_golden_model_1.TH1 [3]);
  nor (_12689_, _12688_, _12687_);
  and (_12691_, _12689_, _12686_);
  and (_12692_, _06389_, \oc8051_golden_model_1.IE [3]);
  not (_12693_, _12692_);
  and (_12694_, _06392_, \oc8051_golden_model_1.SCON [3]);
  and (_12695_, _06394_, \oc8051_golden_model_1.SBUF [3]);
  nor (_12696_, _12695_, _12694_);
  and (_12697_, _12696_, _12693_);
  and (_12698_, _06432_, \oc8051_golden_model_1.ACC [3]);
  and (_12699_, _06435_, \oc8051_golden_model_1.IP [3]);
  nor (_12700_, _12699_, _12698_);
  and (_12701_, _06427_, \oc8051_golden_model_1.PSW [3]);
  and (_12702_, _06429_, \oc8051_golden_model_1.B [3]);
  nor (_12703_, _12702_, _12701_);
  and (_12704_, _12703_, _12700_);
  and (_12705_, _12704_, _12697_);
  and (_12706_, _12705_, _12691_);
  and (_12707_, _06409_, \oc8051_golden_model_1.TH0 [3]);
  and (_12708_, _06411_, \oc8051_golden_model_1.TL1 [3]);
  nor (_12709_, _12708_, _12707_);
  and (_12710_, _06416_, \oc8051_golden_model_1.PCON [3]);
  and (_12712_, _06418_, \oc8051_golden_model_1.TCON [3]);
  nor (_12713_, _12712_, _12710_);
  and (_12714_, _12713_, _12709_);
  and (_12715_, _06368_, \oc8051_golden_model_1.SP [3]);
  not (_12716_, _12715_);
  and (_12717_, _06356_, \oc8051_golden_model_1.P0INREG [3]);
  not (_12718_, _12717_);
  and (_12719_, _06378_, \oc8051_golden_model_1.P1INREG [3]);
  and (_12720_, _06382_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_12721_, _12720_, _12719_);
  and (_12722_, _12721_, _12718_);
  and (_12723_, _06372_, \oc8051_golden_model_1.TMOD [3]);
  and (_12724_, _06361_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_12725_, _12724_, _12723_);
  and (_12726_, _12725_, _12722_);
  and (_12727_, _12726_, _12716_);
  and (_12728_, _12727_, _12714_);
  and (_12729_, _12728_, _12706_);
  not (_12730_, _12729_);
  nor (_12731_, _12730_, _12683_);
  nor (_12732_, _12731_, _06242_);
  or (_12733_, _12732_, _06246_);
  or (_12734_, _12733_, _12682_);
  and (_12735_, _06246_, _03494_);
  nor (_12736_, _12735_, _04583_);
  and (_12737_, _12736_, _12734_);
  and (_12738_, _04583_, _06347_);
  or (_12739_, _12738_, _03227_);
  or (_12740_, _12739_, _12737_);
  and (_12741_, _03227_, _03211_);
  nor (_12742_, _12741_, _04592_);
  and (_12743_, _12742_, _12740_);
  nor (_12744_, _05649_, _03766_);
  and (_12745_, _05649_, _03766_);
  nor (_12746_, _12745_, _12744_);
  and (_12747_, _12746_, _04592_);
  or (_12748_, _12747_, _04590_);
  or (_12749_, _12748_, _12743_);
  and (_12750_, _12749_, _12620_);
  or (_12751_, _12750_, _04597_);
  or (_12752_, _12744_, _05926_);
  and (_12753_, _12752_, _05925_);
  and (_12754_, _12753_, _12751_);
  and (_12755_, _12617_, _04595_);
  or (_12756_, _12755_, _03238_);
  or (_12757_, _12756_, _12754_);
  and (_12758_, _03238_, _03211_);
  nor (_12759_, _12758_, _04609_);
  and (_12760_, _12759_, _12757_);
  nor (_12761_, _12745_, _06471_);
  or (_12762_, _12761_, _04607_);
  or (_12763_, _12762_, _12760_);
  nand (_12764_, _12618_, _04607_);
  and (_12765_, _12764_, _06475_);
  and (_12766_, _12765_, _12763_);
  or (_12767_, _12766_, _12616_);
  and (_12768_, _12767_, _12216_);
  and (_12769_, _12628_, _06481_);
  or (_12770_, _12769_, _04781_);
  or (_12771_, _12770_, _12768_);
  not (_12772_, _04781_);
  or (_12773_, _12628_, _12772_);
  and (_12774_, _12773_, _06486_);
  and (_12775_, _12774_, _12771_);
  or (_12776_, _12775_, _12615_);
  and (_12777_, _12776_, _04811_);
  nor (_12778_, _12625_, _04811_);
  or (_12779_, _12778_, _03686_);
  or (_12780_, _12779_, _12777_);
  nand (_12781_, _11463_, _03686_);
  and (_12782_, _12781_, _12381_);
  and (_12783_, _12782_, _12780_);
  and (_12784_, _03243_, _03210_);
  or (_12785_, _04624_, _12784_);
  or (_12786_, _12785_, _12783_);
  not (_12787_, _05912_);
  or (_12788_, _12670_, _12180_);
  and (_12789_, _12788_, _12787_);
  and (_12790_, _12789_, _12786_);
  nor (_12791_, _07890_, _07888_);
  nor (_12792_, _12791_, _05901_);
  and (_12793_, _12792_, _05912_);
  or (_12794_, _12793_, _04642_);
  or (_12795_, _12794_, _12790_);
  not (_12796_, _04642_);
  or (_12797_, _12792_, _12796_);
  and (_12798_, _12797_, _06833_);
  and (_12799_, _12798_, _12795_);
  or (_12800_, _07991_, _06838_);
  nor (_12801_, _06841_, _06833_);
  and (_12802_, _12801_, _12800_);
  or (_12803_, _12802_, _04633_);
  or (_12804_, _12803_, _12799_);
  nor (_12805_, _05794_, _05650_);
  nor (_12806_, _12805_, _05795_);
  or (_12807_, _12806_, _04805_);
  and (_12808_, _12807_, _05227_);
  and (_12809_, _12808_, _12804_);
  or (_12810_, _12809_, _12213_);
  and (_12811_, _12810_, _12612_);
  and (_12812_, _11427_, _03686_);
  and (_12813_, _11582_, _11956_);
  or (_12814_, _12813_, _12812_);
  and (_12815_, _12814_, _12202_);
  or (_40795_, _12815_, _12811_);
  or (_12816_, _12197_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_12817_, _12816_, _12203_);
  and (_12818_, _06180_, _05888_);
  nor (_12819_, _06180_, _05888_);
  nor (_12820_, _12819_, _12818_);
  nand (_12821_, _12820_, _04617_);
  nor (_12822_, _06047_, _05840_);
  and (_12823_, _06047_, _05840_);
  or (_12824_, _12823_, _12822_);
  or (_12825_, _12824_, _12216_);
  nor (_12826_, _09804_, _09781_);
  and (_12827_, _09781_, \oc8051_golden_model_1.PSW [7]);
  nor (_12828_, _12827_, _12826_);
  nor (_12829_, _12828_, _05007_);
  nand (_12830_, _09782_, _10180_);
  or (_12831_, _12830_, _06040_);
  or (_12832_, _12824_, _06054_);
  and (_12833_, _11611_, _03947_);
  nor (_12834_, _03947_, _07536_);
  nor (_12835_, _12834_, _12833_);
  nand (_12836_, _12835_, _06054_);
  and (_12837_, _12836_, _12832_);
  or (_12838_, _12837_, _04509_);
  or (_12839_, _06843_, _06068_);
  and (_12840_, _12839_, _12838_);
  or (_12841_, _12840_, _04516_);
  nand (_12842_, _12820_, _04516_);
  and (_12843_, _12842_, _12841_);
  or (_12844_, _12843_, _04514_);
  and (_12845_, _12844_, _12831_);
  or (_12846_, _12845_, _04857_);
  nor (_12847_, _11611_, _03257_);
  nor (_12848_, _12847_, _04525_);
  and (_12849_, _12848_, _12846_);
  and (_12850_, _07872_, _04525_);
  or (_12851_, _12850_, _04533_);
  or (_12852_, _12851_, _12849_);
  nor (_12853_, _09781_, _10180_);
  or (_12854_, _12853_, _06028_);
  and (_12855_, _12854_, _12852_);
  or (_12856_, _12855_, _03510_);
  nand (_12857_, _08269_, _03510_);
  and (_12858_, _12857_, _03508_);
  and (_12859_, _12858_, _12856_);
  not (_12860_, _10181_);
  and (_12861_, _12830_, _12860_);
  and (_12862_, _12861_, _03507_);
  or (_12863_, _12862_, _12859_);
  and (_12864_, _12863_, _03253_);
  or (_12865_, _11612_, _03253_);
  nand (_12866_, _12865_, _03593_);
  or (_12867_, _12866_, _12864_);
  nand (_12868_, _08269_, _03594_);
  and (_12869_, _12868_, _12867_);
  or (_12870_, _12869_, _04551_);
  and (_12871_, _06843_, _04559_);
  nand (_12872_, _08268_, _04551_);
  or (_12873_, _12872_, _12871_);
  and (_12874_, _12873_, _05007_);
  and (_12875_, _12874_, _12870_);
  or (_12876_, _12875_, _12829_);
  and (_12877_, _12876_, _03278_);
  or (_12878_, _11612_, _03278_);
  nand (_12879_, _12878_, _04568_);
  or (_12880_, _12879_, _12877_);
  nand (_12881_, _05840_, _06238_);
  and (_12882_, _12881_, _12880_);
  or (_12883_, _12882_, _05971_);
  and (_12884_, _06843_, _06242_);
  or (_12885_, _12884_, _04571_);
  and (_12886_, _12885_, _12883_);
  nor (_12887_, _06247_, _05840_);
  and (_12888_, _06350_, \oc8051_golden_model_1.TL0 [4]);
  not (_12889_, _12888_);
  and (_12890_, _06356_, \oc8051_golden_model_1.P0INREG [4]);
  and (_12891_, _06361_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_12892_, _12891_, _12890_);
  and (_12893_, _12892_, _12889_);
  and (_12894_, _06368_, \oc8051_golden_model_1.SP [4]);
  not (_12895_, _12894_);
  and (_12896_, _06372_, \oc8051_golden_model_1.TMOD [4]);
  not (_12897_, _12896_);
  and (_12898_, _06378_, \oc8051_golden_model_1.P1INREG [4]);
  and (_12899_, _06382_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_12900_, _12899_, _12898_);
  and (_12901_, _12900_, _12897_);
  and (_12902_, _12901_, _12895_);
  and (_12903_, _12902_, _12893_);
  and (_12904_, _06389_, \oc8051_golden_model_1.IE [4]);
  not (_12905_, _12904_);
  and (_12906_, _06392_, \oc8051_golden_model_1.SCON [4]);
  and (_12907_, _06394_, \oc8051_golden_model_1.SBUF [4]);
  nor (_12908_, _12907_, _12906_);
  and (_12909_, _12908_, _12905_);
  and (_12910_, _06400_, \oc8051_golden_model_1.DPH [4]);
  and (_12911_, _06404_, \oc8051_golden_model_1.TH1 [4]);
  nor (_12912_, _12911_, _12910_);
  and (_12913_, _12912_, _12909_);
  and (_12914_, _12913_, _12903_);
  and (_12915_, _06422_, \oc8051_golden_model_1.DPL [4]);
  not (_12916_, _12915_);
  and (_12917_, _06427_, \oc8051_golden_model_1.PSW [4]);
  and (_12918_, _06429_, \oc8051_golden_model_1.B [4]);
  nor (_12919_, _12918_, _12917_);
  and (_12920_, _06432_, \oc8051_golden_model_1.ACC [4]);
  and (_12921_, _06435_, \oc8051_golden_model_1.IP [4]);
  nor (_12922_, _12921_, _12920_);
  and (_12923_, _12922_, _12919_);
  and (_12924_, _12923_, _12916_);
  and (_12925_, _06388_, _06346_);
  and (_12926_, _12925_, \oc8051_golden_model_1.TCON [4]);
  and (_12927_, _06409_, \oc8051_golden_model_1.TH0 [4]);
  nor (_12928_, _12927_, _12926_);
  and (_12929_, _06416_, \oc8051_golden_model_1.PCON [4]);
  and (_12930_, _06411_, \oc8051_golden_model_1.TL1 [4]);
  nor (_12931_, _12930_, _12929_);
  and (_12932_, _12931_, _12928_);
  and (_12933_, _12932_, _12924_);
  and (_12934_, _12933_, _12914_);
  not (_12935_, _12934_);
  nor (_12936_, _12935_, _12887_);
  nor (_12937_, _12936_, _06242_);
  or (_12938_, _12937_, _06246_);
  or (_12939_, _12938_, _12886_);
  and (_12940_, _06246_, _04308_);
  nor (_12941_, _12940_, _04583_);
  and (_12942_, _12941_, _12939_);
  and (_12943_, _06375_, _04583_);
  or (_12944_, _12943_, _03227_);
  or (_12945_, _12944_, _12942_);
  and (_12946_, _11612_, _03227_);
  nor (_12947_, _12946_, _04592_);
  and (_12948_, _12947_, _12945_);
  and (_12949_, _06344_, _05888_);
  nor (_12950_, _06344_, _05888_);
  nor (_12951_, _12950_, _12949_);
  and (_12952_, _12951_, _04592_);
  or (_12953_, _12952_, _04590_);
  or (_12954_, _12953_, _12948_);
  nor (_12955_, _05888_, _07536_);
  and (_12956_, _05888_, _07536_);
  nor (_12957_, _12956_, _12955_);
  or (_12958_, _12957_, _05927_);
  and (_12959_, _12958_, _05926_);
  and (_12960_, _12959_, _12954_);
  and (_12961_, _12950_, _04597_);
  or (_12962_, _12961_, _04595_);
  or (_12963_, _12962_, _12960_);
  or (_12964_, _12955_, _05925_);
  and (_12965_, _12964_, _12963_);
  or (_12966_, _12965_, _03238_);
  and (_12967_, _11612_, _03238_);
  nor (_12968_, _12967_, _04609_);
  and (_12969_, _12968_, _12966_);
  nor (_12970_, _12949_, _06471_);
  or (_12971_, _12970_, _04607_);
  or (_12972_, _12971_, _12969_);
  nand (_12973_, _12956_, _04607_);
  and (_12974_, _12973_, _06475_);
  and (_12975_, _12974_, _12972_);
  and (_12976_, _11611_, _03248_);
  or (_12977_, _12976_, _06481_);
  or (_12978_, _12977_, _12975_);
  and (_12979_, _12978_, _12825_);
  or (_12980_, _12979_, _04781_);
  or (_12981_, _12824_, _12772_);
  and (_12982_, _12981_, _06486_);
  and (_12983_, _12982_, _12980_);
  and (_12984_, _06716_, _06806_);
  nor (_12985_, _06716_, _06806_);
  or (_12986_, _12985_, _12984_);
  and (_12987_, _12986_, _04618_);
  or (_12988_, _12987_, _04617_);
  or (_12989_, _12988_, _12983_);
  and (_12990_, _12989_, _12821_);
  or (_12991_, _12990_, _03686_);
  nand (_12992_, _11459_, _03686_);
  and (_12993_, _12992_, _12381_);
  and (_12994_, _12993_, _12991_);
  and (_12995_, _11611_, _03243_);
  or (_12996_, _12995_, _04624_);
  or (_12997_, _12996_, _12994_);
  or (_12998_, _12826_, _12180_);
  and (_12999_, _12998_, _05913_);
  and (_13000_, _12999_, _12997_);
  or (_13001_, _05901_, _07872_);
  and (_13002_, _05901_, _07872_);
  nor (_13003_, _05913_, _13002_);
  and (_13004_, _13003_, _13001_);
  or (_13005_, _13004_, _13000_);
  and (_13006_, _13005_, _06833_);
  or (_13007_, _06841_, _06843_);
  nor (_13008_, _07968_, _06833_);
  and (_13009_, _13008_, _13007_);
  or (_13010_, _13009_, _04633_);
  or (_13011_, _13010_, _13006_);
  nor (_13012_, _05889_, _05795_);
  nor (_13013_, _13012_, _05890_);
  or (_13014_, _13013_, _04805_);
  and (_13015_, _13014_, _05227_);
  and (_13016_, _13015_, _13011_);
  or (_13017_, _13016_, _12213_);
  and (_13018_, _13017_, _12817_);
  and (_13019_, _11418_, _03686_);
  not (_13020_, _11575_);
  nor (_13021_, _13020_, _03686_);
  or (_13022_, _13021_, _13019_);
  and (_13023_, _13022_, _12202_);
  or (_40796_, _13023_, _13018_);
  nor (_13024_, _12010_, _05492_);
  nor (_13025_, _07968_, _06842_);
  nor (_13026_, _13025_, _06845_);
  or (_13027_, _13026_, _06833_);
  nor (_13028_, _09910_, _09886_);
  and (_13029_, _09886_, \oc8051_golden_model_1.PSW [7]);
  nor (_13030_, _13029_, _13028_);
  nor (_13031_, _13030_, _05007_);
  nor (_13032_, _09886_, _10228_);
  or (_13033_, _13032_, _06028_);
  nor (_13034_, _12818_, _05600_);
  nor (_13035_, _13034_, _06181_);
  nor (_13036_, _13035_, _06175_);
  or (_13037_, _06842_, _06068_);
  nor (_13038_, _12823_, _05552_);
  or (_13039_, _13038_, _06048_);
  and (_13040_, _13039_, _12226_);
  nand (_13041_, _11607_, _03947_);
  or (_13042_, _03947_, \oc8051_golden_model_1.ACC [5]);
  and (_13043_, _13042_, _13041_);
  and (_13044_, _13043_, _06054_);
  or (_13045_, _13044_, _04509_);
  or (_13046_, _13045_, _13040_);
  and (_13047_, _13046_, _06175_);
  and (_13048_, _13047_, _13037_);
  or (_13049_, _13048_, _13036_);
  and (_13050_, _13049_, _06040_);
  nand (_13051_, _09887_, _10228_);
  and (_13052_, _13051_, _04514_);
  or (_13053_, _13052_, _04857_);
  or (_13054_, _13053_, _13050_);
  nor (_13055_, _11606_, _03257_);
  nor (_13056_, _13055_, _04525_);
  and (_13057_, _13056_, _13054_);
  and (_13058_, _07871_, _04525_);
  or (_13059_, _13058_, _04533_);
  or (_13060_, _13059_, _13057_);
  and (_13061_, _13060_, _13033_);
  or (_13062_, _13061_, _03510_);
  nand (_13063_, _08255_, _03510_);
  and (_13064_, _13063_, _03508_);
  and (_13065_, _13064_, _13062_);
  not (_13066_, _10229_);
  and (_13067_, _13051_, _13066_);
  and (_13068_, _13067_, _03507_);
  or (_13069_, _13068_, _13065_);
  and (_13070_, _13069_, _03253_);
  or (_13071_, _11607_, _03253_);
  nand (_13072_, _13071_, _03593_);
  or (_13073_, _13072_, _13070_);
  nand (_13074_, _08255_, _03594_);
  and (_13075_, _13074_, _13073_);
  or (_13076_, _13075_, _04551_);
  and (_13077_, _06842_, _04559_);
  nand (_13078_, _08254_, _04551_);
  or (_13079_, _13078_, _13077_);
  and (_13080_, _13079_, _05007_);
  and (_13081_, _13080_, _13076_);
  or (_13082_, _13081_, _13031_);
  and (_13083_, _13082_, _03278_);
  or (_13084_, _11607_, _03278_);
  nand (_13085_, _13084_, _04568_);
  or (_13086_, _13085_, _13083_);
  nand (_13087_, _05552_, _06238_);
  and (_13088_, _13087_, _13086_);
  or (_13089_, _13088_, _05971_);
  and (_13090_, _06842_, _06242_);
  or (_13091_, _13090_, _04571_);
  and (_13092_, _13091_, _13089_);
  nor (_13093_, _06247_, _05552_);
  and (_13094_, _06368_, \oc8051_golden_model_1.SP [5]);
  not (_13095_, _13094_);
  and (_13096_, _06350_, \oc8051_golden_model_1.TL0 [5]);
  not (_13097_, _13096_);
  and (_13098_, _06378_, \oc8051_golden_model_1.P1INREG [5]);
  and (_13099_, _06382_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_13100_, _13099_, _13098_);
  and (_13101_, _13100_, _13097_);
  and (_13102_, _06356_, \oc8051_golden_model_1.P0INREG [5]);
  and (_13103_, _06361_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_13104_, _13103_, _13102_);
  and (_13105_, _13104_, _13101_);
  and (_13106_, _13105_, _13095_);
  and (_13107_, _06389_, \oc8051_golden_model_1.IE [5]);
  not (_13108_, _13107_);
  and (_13109_, _06392_, \oc8051_golden_model_1.SCON [5]);
  and (_13110_, _06394_, \oc8051_golden_model_1.SBUF [5]);
  nor (_13111_, _13110_, _13109_);
  and (_13112_, _13111_, _13108_);
  and (_13113_, _06427_, \oc8051_golden_model_1.PSW [5]);
  and (_13114_, _06429_, \oc8051_golden_model_1.B [5]);
  nor (_13115_, _13114_, _13113_);
  and (_13116_, _06432_, \oc8051_golden_model_1.ACC [5]);
  and (_13117_, _06435_, \oc8051_golden_model_1.IP [5]);
  nor (_13118_, _13117_, _13116_);
  and (_13119_, _13118_, _13115_);
  and (_13120_, _13119_, _13112_);
  and (_13121_, _13120_, _13106_);
  and (_13122_, _06409_, \oc8051_golden_model_1.TH0 [5]);
  and (_13123_, _06411_, \oc8051_golden_model_1.TL1 [5]);
  nor (_13124_, _13123_, _13122_);
  and (_13125_, _06416_, \oc8051_golden_model_1.PCON [5]);
  and (_13126_, _06418_, \oc8051_golden_model_1.TCON [5]);
  nor (_13127_, _13126_, _13125_);
  and (_13128_, _13127_, _13124_);
  and (_13129_, _06372_, \oc8051_golden_model_1.TMOD [5]);
  and (_13130_, _06404_, \oc8051_golden_model_1.TH1 [5]);
  nor (_13131_, _13130_, _13129_);
  and (_13132_, _06422_, \oc8051_golden_model_1.DPL [5]);
  and (_13133_, _06400_, \oc8051_golden_model_1.DPH [5]);
  nor (_13134_, _13133_, _13132_);
  and (_13135_, _13134_, _13131_);
  and (_13136_, _13135_, _13128_);
  and (_13137_, _13136_, _13121_);
  not (_13138_, _13137_);
  nor (_13139_, _13138_, _13093_);
  nor (_13140_, _13139_, _06242_);
  or (_13141_, _13140_, _06246_);
  or (_13142_, _13141_, _13092_);
  and (_13143_, _06246_, _03853_);
  nor (_13144_, _13143_, _04583_);
  and (_13145_, _13144_, _13142_);
  and (_13146_, _06358_, _04583_);
  or (_13147_, _13146_, _03227_);
  or (_13148_, _13147_, _13145_);
  and (_13149_, _11607_, _03227_);
  nor (_13150_, _13149_, _04592_);
  and (_13151_, _13150_, _13148_);
  and (_13152_, _06313_, _05600_);
  nor (_13153_, _06313_, _05600_);
  nor (_13154_, _13153_, _13152_);
  and (_13155_, _13154_, _04592_);
  or (_13156_, _13155_, _04590_);
  or (_13157_, _13156_, _13151_);
  nor (_13158_, _05600_, _07530_);
  and (_13159_, _05600_, _07530_);
  nor (_13160_, _13159_, _13158_);
  or (_13161_, _13160_, _05927_);
  and (_13162_, _13161_, _05926_);
  and (_13163_, _13162_, _13157_);
  and (_13164_, _13153_, _04597_);
  or (_13165_, _13164_, _13163_);
  and (_13166_, _13165_, _05925_);
  and (_13167_, _13158_, _04595_);
  or (_13168_, _13167_, _03238_);
  or (_13169_, _13168_, _13166_);
  and (_13170_, _11607_, _03238_);
  nor (_13171_, _13170_, _04609_);
  and (_13172_, _13171_, _13169_);
  nor (_13173_, _13152_, _06471_);
  or (_13174_, _13173_, _04607_);
  or (_13175_, _13174_, _13172_);
  nand (_13176_, _13159_, _04607_);
  and (_13177_, _13176_, _06475_);
  and (_13178_, _13177_, _13175_);
  and (_13179_, _11606_, _03248_);
  and (_13180_, _03589_, _03066_);
  or (_13181_, _06479_, _13180_);
  or (_13182_, _13181_, _13179_);
  or (_13183_, _13182_, _06480_);
  or (_13184_, _13183_, _13178_);
  not (_13185_, _04250_);
  and (_13186_, _13039_, _13185_);
  or (_13187_, _13186_, _06814_);
  and (_13188_, _13187_, _13184_);
  and (_13189_, _13039_, _04250_);
  or (_13190_, _13189_, _04618_);
  or (_13191_, _13190_, _13188_);
  nor (_13192_, _12984_, _06761_);
  or (_13193_, _06808_, _06486_);
  or (_13194_, _13193_, _13192_);
  and (_13195_, _13194_, _04811_);
  and (_13196_, _13195_, _13191_);
  nor (_13197_, _13035_, _04811_);
  or (_13198_, _13197_, _03686_);
  or (_13199_, _13198_, _13196_);
  nand (_13200_, _11454_, _03686_);
  and (_13201_, _13200_, _12381_);
  and (_13202_, _13201_, _13199_);
  and (_13203_, _11606_, _03243_);
  or (_13204_, _13203_, _04624_);
  or (_13205_, _13204_, _13202_);
  or (_13206_, _13028_, _12180_);
  and (_13207_, _13206_, _05913_);
  and (_13208_, _13207_, _13205_);
  or (_13209_, _13002_, _07871_);
  nor (_13210_, _05913_, _05903_);
  and (_13211_, _13210_, _13209_);
  or (_13212_, _13211_, _04271_);
  or (_13213_, _13212_, _13208_);
  and (_13214_, _13213_, _13027_);
  or (_13215_, _13214_, _04633_);
  nor (_13216_, _05890_, _05601_);
  nor (_13217_, _13216_, _05891_);
  or (_13218_, _13217_, _04805_);
  and (_13219_, _13218_, _04891_);
  and (_13220_, _13219_, _13215_);
  and (_13221_, _13220_, _12010_);
  or (_13222_, _13221_, _13024_);
  and (_13223_, _13222_, _12203_);
  and (_13224_, _11413_, _03686_);
  and (_13225_, _11571_, _11956_);
  or (_13226_, _13225_, _13224_);
  and (_13227_, _13226_, _12202_);
  or (_40797_, _13227_, _13223_);
  or (_13228_, _12197_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_13229_, _13228_, _12203_);
  and (_13230_, _05903_, _05442_);
  nor (_13231_, _05903_, _05442_);
  or (_13232_, _13231_, _13230_);
  or (_13233_, _13232_, _12787_);
  nor (_13234_, _06181_, _05490_);
  nor (_13235_, _13234_, _06182_);
  nor (_13236_, _13235_, _04811_);
  nor (_13237_, _06808_, _06532_);
  or (_13238_, _13237_, _06809_);
  and (_13239_, _13238_, _04618_);
  nor (_13240_, _06048_, _05442_);
  or (_13241_, _13240_, _06049_);
  or (_13242_, _13241_, _12216_);
  and (_13243_, _06281_, _05490_);
  nor (_13244_, _06281_, _05490_);
  nor (_13245_, _13244_, _13243_);
  and (_13246_, _13245_, _04592_);
  nor (_13247_, _09858_, _09834_);
  and (_13248_, _09834_, \oc8051_golden_model_1.PSW [7]);
  nor (_13249_, _13248_, _13247_);
  nor (_13250_, _13249_, _05007_);
  nor (_13251_, _09834_, _10204_);
  or (_13252_, _13251_, _06028_);
  or (_13253_, _13241_, _06054_);
  nor (_13254_, _03947_, _07484_);
  and (_13255_, _11598_, _03947_);
  nor (_13256_, _13255_, _13254_);
  nand (_13257_, _13256_, _06054_);
  and (_13258_, _13257_, _13253_);
  or (_13259_, _13258_, _04509_);
  or (_13260_, _06531_, _06068_);
  and (_13261_, _13260_, _13259_);
  and (_13262_, _13261_, _06175_);
  nor (_13263_, _13235_, _06175_);
  or (_13264_, _13263_, _13262_);
  and (_13265_, _13264_, _06040_);
  nand (_13266_, _09835_, _10204_);
  and (_13267_, _13266_, _04514_);
  or (_13268_, _13267_, _04857_);
  or (_13269_, _13268_, _13265_);
  nor (_13270_, _11598_, _03257_);
  nor (_13271_, _13270_, _04525_);
  and (_13272_, _13271_, _13269_);
  and (_13273_, _07856_, _04525_);
  or (_13274_, _13273_, _04533_);
  or (_13275_, _13274_, _13272_);
  and (_13276_, _13275_, _13252_);
  or (_13277_, _13276_, _03510_);
  nand (_13278_, _08173_, _03510_);
  and (_13279_, _13278_, _03508_);
  and (_13280_, _13279_, _13277_);
  not (_13281_, _10205_);
  and (_13282_, _13266_, _13281_);
  and (_13283_, _13282_, _03507_);
  or (_13284_, _13283_, _13280_);
  and (_13285_, _13284_, _03253_);
  or (_13286_, _11599_, _03253_);
  nand (_13287_, _13286_, _03593_);
  or (_13288_, _13287_, _13285_);
  nand (_13289_, _08173_, _03594_);
  and (_13290_, _13289_, _13288_);
  or (_13291_, _13290_, _04551_);
  and (_13292_, _06531_, _04559_);
  nand (_13293_, _08172_, _04551_);
  or (_13294_, _13293_, _13292_);
  and (_13295_, _13294_, _05007_);
  and (_13296_, _13295_, _13291_);
  or (_13297_, _13296_, _13250_);
  and (_13298_, _13297_, _03278_);
  or (_13299_, _11599_, _03278_);
  nand (_13300_, _13299_, _04568_);
  or (_13301_, _13300_, _13298_);
  nand (_13302_, _05442_, _06238_);
  and (_13303_, _13302_, _13301_);
  or (_13304_, _13303_, _05971_);
  and (_13305_, _06531_, _06242_);
  or (_13306_, _13305_, _04571_);
  and (_13307_, _13306_, _13304_);
  nor (_13308_, _06247_, _05442_);
  and (_13309_, _06350_, \oc8051_golden_model_1.TL0 [6]);
  not (_13310_, _13309_);
  and (_13311_, _06356_, \oc8051_golden_model_1.P0INREG [6]);
  and (_13312_, _06361_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_13313_, _13312_, _13311_);
  and (_13314_, _13313_, _13310_);
  and (_13315_, _06368_, \oc8051_golden_model_1.SP [6]);
  not (_13316_, _13315_);
  and (_13317_, _06372_, \oc8051_golden_model_1.TMOD [6]);
  not (_13318_, _13317_);
  and (_13319_, _06378_, \oc8051_golden_model_1.P1INREG [6]);
  and (_13320_, _06382_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_13321_, _13320_, _13319_);
  and (_13322_, _13321_, _13318_);
  and (_13323_, _13322_, _13316_);
  and (_13324_, _13323_, _13314_);
  and (_13325_, _06389_, \oc8051_golden_model_1.IE [6]);
  not (_13326_, _13325_);
  and (_13327_, _06392_, \oc8051_golden_model_1.SCON [6]);
  and (_13328_, _06394_, \oc8051_golden_model_1.SBUF [6]);
  nor (_13329_, _13328_, _13327_);
  and (_13330_, _13329_, _13326_);
  and (_13331_, _06400_, \oc8051_golden_model_1.DPH [6]);
  and (_13332_, _06404_, \oc8051_golden_model_1.TH1 [6]);
  nor (_13333_, _13332_, _13331_);
  and (_13334_, _13333_, _13330_);
  and (_13335_, _13334_, _13324_);
  and (_13336_, _06409_, \oc8051_golden_model_1.TH0 [6]);
  and (_13337_, _06411_, \oc8051_golden_model_1.TL1 [6]);
  nor (_13338_, _13337_, _13336_);
  and (_13339_, _06416_, \oc8051_golden_model_1.PCON [6]);
  and (_13340_, _06418_, \oc8051_golden_model_1.TCON [6]);
  nor (_13341_, _13340_, _13339_);
  and (_13342_, _13341_, _13338_);
  and (_13343_, _06422_, \oc8051_golden_model_1.DPL [6]);
  not (_13344_, _13343_);
  and (_13345_, _06429_, \oc8051_golden_model_1.B [6]);
  and (_13346_, _06435_, \oc8051_golden_model_1.IP [6]);
  nor (_13347_, _13346_, _13345_);
  and (_13348_, _06427_, \oc8051_golden_model_1.PSW [6]);
  and (_13349_, _06432_, \oc8051_golden_model_1.ACC [6]);
  nor (_13350_, _13349_, _13348_);
  and (_13351_, _13350_, _13347_);
  and (_13352_, _13351_, _13344_);
  and (_13353_, _13352_, _13342_);
  and (_13354_, _13353_, _13335_);
  not (_13355_, _13354_);
  nor (_13356_, _13355_, _13308_);
  nor (_13357_, _13356_, _06242_);
  or (_13358_, _13357_, _06246_);
  or (_13359_, _13358_, _13307_);
  and (_13360_, _06246_, _03556_);
  nor (_13361_, _13360_, _04583_);
  and (_13362_, _13361_, _13359_);
  not (_13363_, _06281_);
  and (_13364_, _13363_, _04583_);
  or (_13365_, _13364_, _03227_);
  or (_13366_, _13365_, _13362_);
  and (_13367_, _11599_, _03227_);
  nor (_13368_, _13367_, _04592_);
  and (_13369_, _13368_, _13366_);
  or (_13370_, _13369_, _13246_);
  and (_13371_, _13370_, _05927_);
  nor (_13372_, _05490_, _07484_);
  and (_13373_, _05490_, _07484_);
  nor (_13374_, _13373_, _13372_);
  and (_13375_, _13374_, _04590_);
  or (_13376_, _13375_, _13371_);
  and (_13377_, _13376_, _05926_);
  and (_13378_, _13244_, _04597_);
  or (_13379_, _13378_, _04595_);
  or (_13380_, _13379_, _13377_);
  or (_13381_, _13372_, _05925_);
  and (_13382_, _13381_, _13380_);
  or (_13383_, _13382_, _03238_);
  and (_13384_, _11599_, _03238_);
  nor (_13385_, _13384_, _04609_);
  and (_13386_, _13385_, _13383_);
  nor (_13387_, _13243_, _06471_);
  or (_13388_, _13387_, _04607_);
  or (_13389_, _13388_, _13386_);
  nand (_13390_, _13373_, _04607_);
  and (_13391_, _13390_, _06475_);
  and (_13392_, _13391_, _13389_);
  and (_13393_, _11598_, _03248_);
  or (_13394_, _13393_, _06481_);
  or (_13395_, _13394_, _13392_);
  and (_13396_, _13395_, _13242_);
  or (_13397_, _13396_, _04781_);
  or (_13398_, _13241_, _12772_);
  and (_13399_, _13398_, _06486_);
  and (_13400_, _13399_, _13397_);
  or (_13401_, _13400_, _13239_);
  and (_13402_, _13401_, _04811_);
  or (_13403_, _13402_, _13236_);
  and (_13404_, _13403_, _11956_);
  and (_13405_, _11445_, _03686_);
  or (_13406_, _13405_, _03243_);
  or (_13407_, _13406_, _13404_);
  and (_13408_, _11599_, _03243_);
  nor (_13409_, _13408_, _04624_);
  and (_13410_, _13409_, _13407_);
  and (_13411_, _13247_, _04624_);
  or (_13412_, _13411_, _05912_);
  or (_13413_, _13412_, _13410_);
  and (_13414_, _13413_, _13233_);
  or (_13415_, _13414_, _04642_);
  or (_13416_, _13232_, _12796_);
  and (_13417_, _13416_, _06833_);
  and (_13418_, _13417_, _13415_);
  or (_13419_, _06845_, _06531_);
  nor (_13420_, _06846_, _06833_);
  and (_13421_, _13420_, _13419_);
  or (_13422_, _13421_, _04633_);
  or (_13423_, _13422_, _13418_);
  nor (_13424_, _05891_, _05491_);
  nor (_13425_, _13424_, _05892_);
  or (_13426_, _13425_, _04805_);
  and (_13427_, _13426_, _04891_);
  and (_13428_, _13427_, _13423_);
  or (_13429_, _13428_, _12213_);
  and (_13430_, _13429_, _13229_);
  and (_13431_, _11406_, _03686_);
  and (_13432_, _11565_, _11956_);
  or (_13433_, _13432_, _13431_);
  and (_13434_, _13433_, _12202_);
  or (_40799_, _13434_, _13430_);
  or (_13435_, _12011_, _06853_);
  or (_13436_, _12197_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_13437_, _13436_, _12203_);
  and (_13438_, _13437_, _13435_);
  and (_13439_, _12202_, _06877_);
  or (_40800_, _13439_, _13438_);
  and (_13440_, _05229_, _04800_);
  and (_13441_, _13440_, _12195_);
  or (_13442_, _13441_, \oc8051_golden_model_1.IRAM[1] [0]);
  nor (_13443_, _12188_, _05228_);
  not (_13444_, _13443_);
  nor (_13445_, _13444_, _12187_);
  not (_13446_, _13441_);
  or (_13447_, _13446_, _13445_);
  nand (_13448_, _13447_, _13442_);
  not (_13449_, _05213_);
  or (_13450_, _05220_, _13449_);
  or (_13451_, _13450_, _43231_);
  nor (_13452_, _13451_, rst);
  not (_13453_, _05216_);
  nor (_13454_, _05220_, _13453_);
  and (_13455_, _13454_, _43227_);
  and (_13456_, _13455_, _41991_);
  nor (_13457_, _13456_, _13452_);
  nor (_13458_, _05220_, _04079_);
  and (_13459_, _13458_, _43227_);
  and (_13460_, _13459_, _41991_);
  not (_13461_, _13460_);
  nor (_13462_, _05220_, \oc8051_golden_model_1.SP [1]);
  and (_13463_, _13462_, _43227_);
  and (_13464_, _13463_, _41991_);
  nor (_13465_, _13464_, _13461_);
  and (_13466_, _13465_, _13457_);
  nor (_13467_, _13466_, _13448_);
  and (_13468_, _12201_, _04948_);
  and (_13469_, _13468_, _12209_);
  or (_40804_, _13469_, _13467_);
  not (_13470_, _13468_);
  or (_13471_, _13441_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_13472_, _13471_, _13470_);
  or (_13473_, _13446_, _12399_);
  and (_13474_, _13473_, _13472_);
  and (_13475_, _13468_, _12405_);
  or (_40806_, _13475_, _13474_);
  or (_13476_, _13441_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_13477_, _13476_, _13470_);
  or (_13478_, _13446_, _12603_);
  and (_13479_, _13478_, _13477_);
  and (_13480_, _13468_, _12609_);
  or (_40807_, _13480_, _13479_);
  or (_13481_, _13441_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_13482_, _13481_, _13470_);
  or (_13483_, _13446_, _12809_);
  and (_13484_, _13483_, _13482_);
  and (_13485_, _13468_, _12814_);
  or (_40808_, _13485_, _13484_);
  or (_13486_, _13441_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_13487_, _13486_, _13470_);
  or (_13488_, _13446_, _13016_);
  and (_13489_, _13488_, _13487_);
  and (_13490_, _13468_, _13022_);
  or (_40809_, _13490_, _13489_);
  and (_13491_, _12005_, _04800_);
  and (_13492_, _13491_, _12008_);
  nor (_13493_, _13492_, _05494_);
  and (_13494_, _13492_, _13220_);
  or (_13495_, _13494_, _13493_);
  and (_13496_, _13495_, _13470_);
  and (_13497_, _13468_, _13226_);
  or (_40810_, _13497_, _13496_);
  or (_13498_, _13441_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_13499_, _13498_, _13470_);
  or (_13500_, _13446_, _13428_);
  and (_13501_, _13500_, _13499_);
  not (_13502_, _05220_);
  and (_13503_, _13433_, _13502_);
  and (_13504_, _13503_, _43227_);
  and (_13505_, _13504_, _41991_);
  and (_13506_, _13466_, _13505_);
  or (_40812_, _13506_, _13501_);
  or (_13507_, _13441_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_13508_, _13507_, _13470_);
  or (_13509_, _13446_, _06854_);
  and (_13510_, _13509_, _13508_);
  and (_13511_, _13468_, _06877_);
  or (_40813_, _13511_, _13510_);
  and (_13512_, _04893_, _04638_);
  and (_13513_, _13512_, _12008_);
  not (_13514_, _13513_);
  or (_13515_, _13514_, _12190_);
  nor (_13516_, _13513_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_13517_, _12201_, _06070_);
  nor (_13518_, _13517_, _13516_);
  and (_13519_, _13518_, _13515_);
  and (_13520_, _12209_, _12199_);
  and (_13521_, _13520_, _13517_);
  or (_40817_, _13521_, _13519_);
  not (_13522_, _13517_);
  or (_13523_, _13513_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_13524_, _13523_, _13522_);
  and (_13525_, _12192_, _04638_);
  and (_13526_, _13525_, _12195_);
  not (_13527_, _13526_);
  or (_13528_, _13527_, _12399_);
  and (_13529_, _13528_, _13524_);
  and (_13530_, _13517_, _12405_);
  or (_40818_, _13530_, _13529_);
  or (_13531_, _13513_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_13532_, _13531_, _13522_);
  and (_13533_, _12601_, _04891_);
  and (_13534_, _13533_, _12598_);
  or (_13535_, _13514_, _13534_);
  and (_13536_, _13535_, _13532_);
  and (_13537_, _13517_, _12609_);
  or (_40819_, _13537_, _13536_);
  and (_13538_, _12814_, _12199_);
  or (_13539_, _13538_, _13522_);
  and (_13540_, _12807_, _04891_);
  and (_13541_, _13540_, _12804_);
  and (_13542_, _13513_, _13541_);
  nor (_13543_, _13513_, _04901_);
  or (_13544_, _13543_, _13517_);
  or (_13545_, _13544_, _13542_);
  and (_40821_, _13545_, _13539_);
  or (_13546_, _13513_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_13547_, _13546_, _13522_);
  and (_13548_, _13014_, _04891_);
  and (_13549_, _13548_, _13011_);
  or (_13550_, _13514_, _13549_);
  and (_13551_, _13550_, _13547_);
  and (_13552_, _13022_, _12199_);
  and (_13553_, _13552_, _13517_);
  or (_40822_, _13553_, _13551_);
  nor (_13554_, _13513_, _05500_);
  and (_13555_, _13513_, _13220_);
  or (_13556_, _13555_, _13554_);
  and (_13557_, _13556_, _13522_);
  and (_13558_, _13226_, _12199_);
  and (_13559_, _13558_, _13517_);
  or (_40823_, _13559_, _13557_);
  or (_13560_, _13513_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_13561_, _13560_, _13522_);
  or (_13562_, _13514_, _13428_);
  and (_13563_, _13562_, _13561_);
  and (_13564_, _13517_, _13433_);
  or (_40824_, _13564_, _13563_);
  or (_13565_, _13513_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_13566_, _13565_, _13522_);
  or (_13567_, _13527_, _06854_);
  and (_13568_, _13567_, _13566_);
  and (_13569_, _06877_, _12199_);
  and (_13570_, _13517_, _13569_);
  or (_40825_, _13570_, _13568_);
  and (_13571_, _12195_, _05231_);
  or (_13572_, _13571_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_13573_, _12201_, _04644_);
  not (_13574_, _13573_);
  and (_13575_, _13574_, _13572_);
  not (_13576_, _13571_);
  or (_13577_, _13576_, _13445_);
  and (_13578_, _13577_, _13575_);
  and (_13579_, _13573_, _13520_);
  or (_40829_, _13579_, _13578_);
  or (_13580_, _13571_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_13581_, _13580_, _13574_);
  or (_13582_, _13576_, _12399_);
  and (_13583_, _13582_, _13581_);
  and (_13584_, _13573_, _12405_);
  or (_40831_, _13584_, _13583_);
  or (_13585_, _13571_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_13586_, _13585_, _13574_);
  or (_13587_, _13576_, _12603_);
  and (_13588_, _13587_, _13586_);
  and (_13589_, _13573_, _12609_);
  or (_40832_, _13589_, _13588_);
  or (_13590_, _13571_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_13591_, _13590_, _13574_);
  or (_13592_, _13576_, _12809_);
  and (_13593_, _13592_, _13591_);
  and (_13594_, _13573_, _13538_);
  or (_40833_, _13594_, _13593_);
  or (_13595_, _13571_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_13596_, _13595_, _13574_);
  or (_13597_, _13576_, _13016_);
  and (_13598_, _13597_, _13596_);
  and (_13599_, _13573_, _13552_);
  or (_40834_, _13599_, _13598_);
  and (_13600_, _12008_, _04894_);
  nor (_13601_, _13600_, _05498_);
  and (_13602_, _13600_, _13220_);
  or (_13603_, _13602_, _13601_);
  and (_13604_, _13603_, _13574_);
  and (_13605_, _13573_, _13558_);
  or (_40835_, _13605_, _13604_);
  or (_13607_, _13571_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_13608_, _13607_, _13574_);
  or (_13609_, _13576_, _13428_);
  and (_13610_, _13609_, _13608_);
  and (_13611_, _13573_, _13433_);
  or (_40837_, _13611_, _13610_);
  or (_13612_, _13571_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_13613_, _13612_, _13574_);
  or (_13614_, _13576_, _06854_);
  and (_13616_, _13614_, _13613_);
  and (_13617_, _13573_, _13569_);
  or (_40838_, _13617_, _13616_);
  and (_13618_, _12194_, _05065_);
  and (_13619_, _13618_, _12193_);
  not (_13620_, _13619_);
  or (_13621_, _13620_, _13445_);
  and (_13622_, _05221_, _05213_);
  and (_13623_, _13622_, _13453_);
  and (_13624_, _13623_, _04645_);
  not (_13626_, _13624_);
  or (_13627_, _13619_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_13628_, _13627_, _13626_);
  and (_13629_, _13628_, _13621_);
  and (_13630_, _12209_, _05221_);
  and (_13631_, _13624_, _13630_);
  or (_40842_, _13631_, _13629_);
  or (_13632_, _13620_, _12399_);
  or (_13633_, _13619_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_13634_, _13633_, _13626_);
  and (_13636_, _13634_, _13632_);
  and (_13637_, _12405_, _05221_);
  and (_13638_, _13637_, _13624_);
  or (_40843_, _13638_, _13636_);
  and (_13639_, _12199_, _05213_);
  and (_13640_, _13639_, _13453_);
  and (_13641_, _13640_, _04645_);
  not (_13642_, _13641_);
  and (_13643_, _05206_, _05065_);
  and (_13644_, _13643_, _12006_);
  or (_13646_, _13644_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_13647_, _13646_, _13642_);
  not (_13648_, _13644_);
  or (_13649_, _13648_, _13534_);
  and (_13650_, _13649_, _13647_);
  and (_13651_, _12609_, _05221_);
  and (_13652_, _13651_, _13624_);
  or (_40844_, _13652_, _13650_);
  or (_13653_, _13620_, _12809_);
  or (_13654_, _13619_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_13656_, _13654_, _13626_);
  and (_13657_, _13656_, _13653_);
  and (_13658_, _12814_, _05221_);
  and (_13659_, _13624_, _13658_);
  or (_40846_, _13659_, _13657_);
  or (_13660_, _13644_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_13661_, _13660_, _13642_);
  or (_13662_, _13648_, _13549_);
  and (_13663_, _13662_, _13661_);
  and (_13664_, _13641_, _13552_);
  or (_40847_, _13664_, _13663_);
  nor (_13666_, _13644_, _05512_);
  and (_13667_, _13644_, _13220_);
  or (_13668_, _13667_, _13666_);
  and (_13669_, _13668_, _13642_);
  and (_13670_, _13641_, _13558_);
  or (_40848_, _13670_, _13669_);
  or (_13671_, _13644_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_13672_, _13671_, _13642_);
  or (_13673_, _13648_, _13428_);
  and (_13675_, _13673_, _13672_);
  and (_13676_, _13433_, _12199_);
  and (_13677_, _13676_, _13641_);
  or (_40849_, _13677_, _13675_);
  or (_13678_, _13644_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_13679_, _13678_, _13642_);
  or (_13680_, _13620_, _06854_);
  and (_13681_, _13680_, _13679_);
  and (_13682_, _13641_, _13569_);
  or (_40850_, _13682_, _13681_);
  and (_13684_, _13643_, _13491_);
  or (_13685_, _13684_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_13686_, _13640_, _04948_);
  not (_13687_, _13686_);
  and (_13688_, _13687_, _13685_);
  not (_13689_, _13684_);
  or (_13690_, _13689_, _12190_);
  and (_13691_, _13690_, _13688_);
  and (_13692_, _13686_, _13520_);
  or (_40854_, _13692_, _13691_);
  and (_13694_, _13618_, _13440_);
  not (_13695_, _13694_);
  or (_13696_, _13695_, _12399_);
  and (_13697_, _13623_, _04948_);
  not (_13698_, _13697_);
  or (_13699_, _13694_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_13700_, _13699_, _13698_);
  and (_13701_, _13700_, _13696_);
  and (_13702_, _13697_, _13637_);
  or (_40855_, _13702_, _13701_);
  or (_13704_, _13684_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_13705_, _13704_, _13687_);
  or (_13706_, _13689_, _13534_);
  and (_13707_, _13706_, _13705_);
  and (_13708_, _13697_, _13651_);
  or (_40857_, _13708_, _13707_);
  or (_13709_, _13695_, _12809_);
  or (_13710_, _13694_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_13711_, _13710_, _13698_);
  and (_13712_, _13711_, _13709_);
  and (_13714_, _13697_, _13658_);
  or (_40858_, _13714_, _13712_);
  or (_13715_, _13684_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_13716_, _13715_, _13687_);
  or (_13717_, _13689_, _13549_);
  and (_13718_, _13717_, _13716_);
  and (_13719_, _13686_, _13552_);
  or (_40859_, _13719_, _13718_);
  nor (_13720_, _13684_, _05514_);
  and (_13721_, _13684_, _13220_);
  or (_13723_, _13721_, _13720_);
  and (_13724_, _13723_, _13687_);
  and (_13725_, _13686_, _13558_);
  or (_40860_, _13725_, _13724_);
  or (_13726_, _13684_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_13727_, _13726_, _13687_);
  or (_13728_, _13689_, _13428_);
  and (_13729_, _13728_, _13727_);
  and (_13730_, _13686_, _13676_);
  or (_40861_, _13730_, _13729_);
  or (_13732_, _13684_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_13733_, _13732_, _13687_);
  or (_13734_, _13695_, _06854_);
  and (_13735_, _13734_, _13733_);
  and (_13736_, _13686_, _13569_);
  or (_40863_, _13736_, _13735_);
  and (_13737_, _13643_, _13512_);
  or (_13738_, _13737_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_13739_, _13640_, _06070_);
  not (_13740_, _13739_);
  and (_13741_, _13740_, _13738_);
  not (_13742_, _13737_);
  or (_13743_, _13742_, _12190_);
  and (_13744_, _13743_, _13741_);
  and (_13745_, _13739_, _13520_);
  or (_40866_, _13745_, _13744_);
  and (_13746_, _13618_, _13525_);
  not (_13747_, _13746_);
  or (_13748_, _13747_, _12399_);
  and (_13749_, _13623_, _06070_);
  not (_13750_, _13749_);
  or (_13751_, _13746_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_13752_, _13751_, _13750_);
  and (_13753_, _13752_, _13748_);
  and (_13754_, _13749_, _13637_);
  or (_40867_, _13754_, _13753_);
  or (_13755_, _13737_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_13756_, _13755_, _13740_);
  or (_13757_, _13742_, _13534_);
  and (_13758_, _13757_, _13756_);
  and (_13759_, _13749_, _13651_);
  or (_40869_, _13759_, _13758_);
  or (_13760_, _13747_, _12809_);
  or (_13761_, _13746_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_13762_, _13761_, _13750_);
  and (_13763_, _13762_, _13760_);
  and (_13764_, _13749_, _13658_);
  or (_40870_, _13764_, _13763_);
  or (_13765_, _13737_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_13766_, _13765_, _13740_);
  or (_13767_, _13742_, _13549_);
  and (_13768_, _13767_, _13766_);
  and (_13769_, _13739_, _13552_);
  or (_40871_, _13769_, _13768_);
  nor (_13770_, _13737_, _05508_);
  and (_13771_, _13737_, _13220_);
  or (_13772_, _13771_, _13770_);
  and (_13773_, _13772_, _13740_);
  and (_13774_, _13739_, _13558_);
  or (_40872_, _13774_, _13773_);
  or (_13775_, _13737_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_13776_, _13775_, _13740_);
  or (_13777_, _13742_, _13428_);
  and (_13778_, _13777_, _13776_);
  and (_13779_, _13739_, _13676_);
  or (_40873_, _13779_, _13778_);
  or (_13780_, _13737_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_13781_, _13780_, _13740_);
  or (_13782_, _13747_, _06854_);
  and (_13783_, _13782_, _13781_);
  and (_13784_, _13739_, _13569_);
  or (_40875_, _13784_, _13783_);
  and (_13785_, _13643_, _04894_);
  not (_13786_, _13785_);
  or (_13787_, _13786_, _12190_);
  or (_13788_, _13785_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_13789_, _13640_, _04644_);
  not (_13790_, _13789_);
  and (_13791_, _13790_, _13788_);
  and (_13792_, _13791_, _13787_);
  and (_13793_, _13789_, _13520_);
  or (_40878_, _13793_, _13792_);
  and (_13794_, _13618_, _05231_);
  not (_13795_, _13794_);
  or (_13796_, _13795_, _12399_);
  and (_13797_, _13623_, _04644_);
  not (_13798_, _13797_);
  or (_13799_, _13794_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_13800_, _13799_, _13798_);
  and (_13801_, _13800_, _13796_);
  and (_13802_, _13797_, _13637_);
  or (_40880_, _13802_, _13801_);
  or (_13803_, _13785_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_13804_, _13803_, _13790_);
  or (_13805_, _13786_, _13534_);
  and (_13806_, _13805_, _13804_);
  and (_13807_, _13797_, _13651_);
  or (_40881_, _13807_, _13806_);
  or (_13808_, _13795_, _12809_);
  or (_13809_, _13794_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_13810_, _13809_, _13798_);
  and (_13811_, _13810_, _13808_);
  and (_13812_, _13797_, _13658_);
  or (_40882_, _13812_, _13811_);
  or (_13813_, _13785_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_13814_, _13813_, _13790_);
  or (_13815_, _13786_, _13549_);
  and (_13816_, _13815_, _13814_);
  and (_13817_, _13789_, _13552_);
  or (_40883_, _13817_, _13816_);
  nor (_13818_, _13785_, _05506_);
  and (_13819_, _13785_, _13220_);
  or (_13820_, _13819_, _13818_);
  and (_13821_, _13820_, _13790_);
  and (_13822_, _13789_, _13558_);
  or (_40884_, _13822_, _13821_);
  or (_13823_, _13785_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_13824_, _13823_, _13790_);
  or (_13825_, _13786_, _13428_);
  and (_13826_, _13825_, _13824_);
  and (_13827_, _13789_, _13676_);
  or (_40886_, _13827_, _13826_);
  or (_13828_, _13785_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_13829_, _13828_, _13790_);
  or (_13830_, _13795_, _06854_);
  and (_13831_, _13830_, _13829_);
  and (_13832_, _13789_, _13569_);
  or (_40887_, _13832_, _13831_);
  and (_13833_, _05233_, _05205_);
  and (_13834_, _13833_, _12193_);
  not (_13835_, _13834_);
  or (_13836_, _13835_, _13445_);
  and (_13837_, _05222_, _13449_);
  and (_13838_, _13837_, _04645_);
  not (_13839_, _13838_);
  or (_13840_, _13834_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_13841_, _13840_, _13839_);
  and (_13842_, _13841_, _13836_);
  and (_13843_, _13838_, _13630_);
  or (_40891_, _13843_, _13842_);
  or (_13844_, _13835_, _12399_);
  or (_13845_, _13834_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_13846_, _13845_, _13839_);
  and (_13847_, _13846_, _13844_);
  and (_13848_, _13838_, _13637_);
  or (_40892_, _13848_, _13847_);
  or (_13849_, _13834_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_13850_, _13849_, _13839_);
  or (_13851_, _13835_, _12603_);
  and (_13852_, _13851_, _13850_);
  and (_13853_, _13838_, _13651_);
  or (_40893_, _13853_, _13852_);
  or (_13854_, _13835_, _12809_);
  or (_13855_, _13834_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_13856_, _13855_, _13839_);
  and (_13857_, _13856_, _13854_);
  and (_13858_, _13838_, _13658_);
  or (_40895_, _13858_, _13857_);
  or (_13859_, _13834_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_13860_, _13859_, _13839_);
  or (_13861_, _13835_, _13016_);
  and (_13862_, _13861_, _13860_);
  and (_13863_, _13022_, _05221_);
  and (_13864_, _13838_, _13863_);
  or (_40896_, _13864_, _13862_);
  and (_13865_, _13218_, _05227_);
  nand (_13866_, _13865_, _13215_);
  nand (_13867_, _13834_, _13866_);
  or (_13868_, _13834_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_13869_, _13868_, _13839_);
  and (_13870_, _13869_, _13867_);
  and (_13871_, _13226_, _05221_);
  and (_13872_, _13838_, _13871_);
  or (_40897_, _13872_, _13870_);
  or (_13873_, _13834_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_13874_, _13873_, _13839_);
  or (_13875_, _13835_, _13428_);
  and (_13876_, _13875_, _13874_);
  and (_13877_, _13433_, _05221_);
  and (_13878_, _13838_, _13877_);
  or (_40898_, _13878_, _13876_);
  or (_13879_, _13834_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_13880_, _13879_, _13839_);
  or (_13881_, _13835_, _06854_);
  and (_13882_, _13881_, _13880_);
  and (_13883_, _13838_, _06878_);
  or (_40899_, _13883_, _13882_);
  and (_13884_, _13833_, _13440_);
  not (_13885_, _13884_);
  or (_13886_, _13885_, _13445_);
  and (_13887_, _13837_, _04948_);
  not (_13888_, _13887_);
  or (_13889_, _13884_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_13890_, _13889_, _13888_);
  and (_13891_, _13890_, _13886_);
  and (_13892_, _13887_, _13630_);
  or (_40903_, _13892_, _13891_);
  or (_13893_, _13885_, _12399_);
  or (_13894_, _13884_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_13895_, _13894_, _13888_);
  and (_13896_, _13895_, _13893_);
  and (_13897_, _13887_, _13637_);
  or (_40904_, _13897_, _13896_);
  or (_13898_, _13884_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_13899_, _13898_, _13888_);
  or (_13900_, _13885_, _12603_);
  and (_13901_, _13900_, _13899_);
  and (_13902_, _13887_, _13651_);
  or (_40906_, _13902_, _13901_);
  or (_13903_, _13885_, _12809_);
  or (_13904_, _13884_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_13905_, _13904_, _13888_);
  and (_13906_, _13905_, _13903_);
  and (_13907_, _13887_, _13658_);
  or (_40907_, _13907_, _13906_);
  or (_13908_, _13884_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_13909_, _13908_, _13888_);
  or (_13910_, _13885_, _13016_);
  and (_13911_, _13910_, _13909_);
  and (_13912_, _13887_, _13863_);
  or (_40908_, _13912_, _13911_);
  nand (_13913_, _13884_, _13866_);
  or (_13914_, _13884_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_13915_, _13914_, _13888_);
  and (_13916_, _13915_, _13913_);
  and (_13917_, _13887_, _13871_);
  or (_40909_, _13917_, _13916_);
  or (_13918_, _13884_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_13919_, _13918_, _13888_);
  or (_13920_, _13885_, _13428_);
  and (_13921_, _13920_, _13919_);
  and (_13922_, _13887_, _13877_);
  or (_40910_, _13922_, _13921_);
  or (_13923_, _13884_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_13924_, _13923_, _13888_);
  or (_13925_, _13885_, _06854_);
  and (_13926_, _13925_, _13924_);
  and (_13927_, _13887_, _06878_);
  or (_40912_, _13927_, _13926_);
  and (_13928_, _13833_, _13525_);
  not (_13929_, _13928_);
  or (_13930_, _13929_, _13445_);
  and (_13931_, _13837_, _06070_);
  not (_13932_, _13931_);
  or (_13933_, _13928_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_13934_, _13933_, _13932_);
  and (_13935_, _13934_, _13930_);
  and (_13936_, _13931_, _13630_);
  or (_40915_, _13936_, _13935_);
  or (_13937_, _13929_, _12399_);
  or (_13938_, _13928_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_13939_, _13938_, _13932_);
  and (_13940_, _13939_, _13937_);
  and (_13941_, _13931_, _13637_);
  or (_40916_, _13941_, _13940_);
  or (_13942_, _13928_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_13943_, _13942_, _13932_);
  or (_13944_, _13929_, _12603_);
  and (_13945_, _13944_, _13943_);
  and (_13946_, _13931_, _13651_);
  or (_40918_, _13946_, _13945_);
  or (_13947_, _13929_, _12809_);
  or (_13948_, _13928_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_13949_, _13948_, _13932_);
  and (_13950_, _13949_, _13947_);
  and (_13951_, _13931_, _13658_);
  or (_40919_, _13951_, _13950_);
  or (_13952_, _13929_, _13016_);
  or (_13953_, _13928_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_13954_, _13953_, _13932_);
  and (_13955_, _13954_, _13952_);
  and (_13956_, _13931_, _13863_);
  or (_40920_, _13956_, _13955_);
  nand (_13957_, _13928_, _13866_);
  or (_13958_, _13928_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_13959_, _13958_, _13932_);
  and (_13960_, _13959_, _13957_);
  and (_13961_, _13931_, _13871_);
  or (_40921_, _13961_, _13960_);
  or (_13962_, _13928_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_13963_, _13962_, _13932_);
  or (_13964_, _13929_, _13428_);
  and (_13965_, _13964_, _13963_);
  and (_13966_, _13931_, _13877_);
  or (_40922_, _13966_, _13965_);
  or (_13967_, _13928_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_13968_, _13967_, _13932_);
  or (_13969_, _13929_, _06854_);
  and (_13970_, _13969_, _13968_);
  and (_13971_, _13931_, _06878_);
  or (_40924_, _13971_, _13970_);
  and (_13972_, _13833_, _05231_);
  or (_13973_, _13972_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_13974_, _13837_, _04644_);
  not (_13975_, _13974_);
  and (_13976_, _13975_, _13973_);
  not (_13977_, _13972_);
  or (_13978_, _13977_, _13445_);
  and (_13979_, _13978_, _13976_);
  and (_13980_, _13974_, _13630_);
  or (_40927_, _13980_, _13979_);
  or (_13981_, _13977_, _12399_);
  or (_13982_, _13972_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_13983_, _13982_, _13975_);
  and (_13984_, _13983_, _13981_);
  and (_13985_, _13974_, _13637_);
  or (_40929_, _13985_, _13984_);
  or (_13986_, _13972_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_13987_, _13986_, _13975_);
  or (_13988_, _13977_, _12603_);
  and (_13989_, _13988_, _13987_);
  and (_13990_, _13974_, _13651_);
  or (_40930_, _13990_, _13989_);
  or (_13991_, _13977_, _12809_);
  or (_13992_, _13972_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_13993_, _13992_, _13975_);
  and (_13994_, _13993_, _13991_);
  and (_13995_, _13974_, _13658_);
  or (_40931_, _13995_, _13994_);
  or (_13996_, _13972_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_13997_, _13996_, _13975_);
  or (_13998_, _13977_, _13016_);
  and (_13999_, _13998_, _13997_);
  and (_14000_, _13974_, _13863_);
  or (_40932_, _14000_, _13999_);
  nand (_14001_, _13972_, _13866_);
  or (_14002_, _13972_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_14003_, _14002_, _13975_);
  and (_14004_, _14003_, _14001_);
  and (_14005_, _13974_, _13871_);
  or (_40933_, _14005_, _14004_);
  or (_14006_, _13972_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_14007_, _14006_, _13975_);
  or (_14008_, _13977_, _13428_);
  and (_14009_, _14008_, _14007_);
  and (_14010_, _13974_, _13877_);
  or (_40935_, _14010_, _14009_);
  or (_14011_, _13972_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_14012_, _14011_, _13975_);
  or (_14013_, _13977_, _06854_);
  and (_14014_, _14013_, _14012_);
  and (_14015_, _13974_, _06878_);
  or (_40936_, _14015_, _14014_);
  and (_14016_, _12006_, _05208_);
  and (_14017_, _14016_, _12190_);
  or (_14018_, _14016_, _04482_);
  not (_14019_, _04645_);
  nand (_14020_, _13639_, _05216_);
  or (_14021_, _14020_, _14019_);
  nand (_14022_, _14021_, _14018_);
  or (_14023_, _14022_, _14017_);
  and (_14024_, _05223_, _04645_);
  not (_14025_, _14024_);
  or (_14026_, _14025_, _13630_);
  and (_40940_, _14026_, _14023_);
  or (_14027_, _14016_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_14028_, _14027_, _14025_);
  and (_14029_, _12193_, _05234_);
  not (_14030_, _14029_);
  or (_14031_, _14030_, _12399_);
  and (_14032_, _14031_, _14028_);
  and (_14033_, _14024_, _13637_);
  or (_40941_, _14033_, _14032_);
  or (_14034_, _14016_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_14035_, _14034_, _14025_);
  not (_14036_, _14016_);
  or (_14037_, _14036_, _13534_);
  and (_14038_, _14037_, _14035_);
  and (_14039_, _14024_, _13651_);
  or (_40942_, _14039_, _14038_);
  or (_14040_, _14016_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_14041_, _14040_, _14025_);
  or (_14042_, _14036_, _13541_);
  and (_14043_, _14042_, _14041_);
  and (_14044_, _14024_, _13658_);
  or (_40943_, _14044_, _14043_);
  or (_14045_, _14016_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_14046_, _14045_, _14025_);
  or (_14047_, _14036_, _13549_);
  and (_14048_, _14047_, _14046_);
  and (_14049_, _14024_, _13863_);
  or (_40944_, _14049_, _14048_);
  nand (_14050_, _14029_, _13866_);
  or (_14051_, _14029_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_14052_, _14051_, _14025_);
  and (_14053_, _14052_, _14050_);
  and (_14054_, _14024_, _13871_);
  or (_40946_, _14054_, _14053_);
  or (_14055_, _14016_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_14056_, _14055_, _14025_);
  or (_14057_, _14036_, _13428_);
  and (_14058_, _14057_, _14056_);
  and (_14059_, _14024_, _13877_);
  or (_40947_, _14059_, _14058_);
  or (_14060_, _14016_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_14061_, _14060_, _14025_);
  or (_14062_, _14030_, _06854_);
  and (_14063_, _14062_, _14061_);
  and (_14064_, _14024_, _06878_);
  or (_40948_, _14064_, _14063_);
  and (_14065_, _13491_, _05208_);
  or (_14066_, _14065_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_14067_, _05223_, _04948_);
  not (_14068_, _14067_);
  and (_14069_, _14068_, _14066_);
  and (_14070_, _13440_, _05234_);
  not (_14071_, _14070_);
  or (_14072_, _14071_, _13445_);
  and (_14073_, _14072_, _14069_);
  and (_14074_, _14067_, _13630_);
  or (_40952_, _14074_, _14073_);
  or (_14075_, _14071_, _12399_);
  or (_14076_, _14070_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_14077_, _14076_, _14068_);
  and (_14078_, _14077_, _14075_);
  and (_14079_, _14067_, _13637_);
  or (_40953_, _14079_, _14078_);
  or (_14080_, _14065_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_14081_, _14080_, _14068_);
  not (_14082_, _14065_);
  or (_14083_, _14082_, _13534_);
  and (_14084_, _14083_, _14081_);
  and (_14085_, _14067_, _13651_);
  or (_40954_, _14085_, _14084_);
  not (_14086_, _04948_);
  or (_14087_, _14020_, _14086_);
  or (_14088_, _14087_, _13538_);
  and (_14089_, _14065_, _13541_);
  or (_14090_, _14065_, _04936_);
  nand (_14091_, _14090_, _14087_);
  or (_14092_, _14091_, _14089_);
  and (_40955_, _14092_, _14088_);
  or (_14093_, _14065_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_14094_, _14093_, _14068_);
  or (_14095_, _14082_, _13549_);
  and (_14096_, _14095_, _14094_);
  and (_14097_, _14067_, _13863_);
  or (_40957_, _14097_, _14096_);
  nand (_14098_, _14070_, _13866_);
  or (_14099_, _14070_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_14100_, _14099_, _14068_);
  and (_14101_, _14100_, _14098_);
  and (_14102_, _14067_, _13871_);
  or (_40958_, _14102_, _14101_);
  or (_14103_, _14065_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_14104_, _14103_, _14068_);
  or (_14105_, _14082_, _13428_);
  and (_14106_, _14105_, _14104_);
  and (_14107_, _14067_, _13877_);
  or (_40959_, _14107_, _14106_);
  or (_14108_, _14065_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_14109_, _14108_, _14068_);
  or (_14110_, _14071_, _06854_);
  and (_14111_, _14110_, _14109_);
  and (_14112_, _14067_, _06878_);
  or (_40960_, _14112_, _14111_);
  and (_14113_, _13512_, _05208_);
  or (_14114_, _14113_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_14115_, _06070_, _05223_);
  not (_14116_, _14115_);
  and (_14117_, _14116_, _14114_);
  and (_14118_, _13525_, _05234_);
  not (_14119_, _14118_);
  or (_14120_, _14119_, _13445_);
  and (_14121_, _14120_, _14117_);
  and (_14122_, _14115_, _13630_);
  or (_40964_, _14122_, _14121_);
  or (_14123_, _14119_, _12399_);
  or (_14124_, _14118_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_14125_, _14124_, _14116_);
  and (_14126_, _14125_, _14123_);
  and (_14127_, _14115_, _13637_);
  or (_40965_, _14127_, _14126_);
  or (_14128_, _14113_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_14129_, _14128_, _14116_);
  not (_14130_, _14113_);
  or (_14131_, _14130_, _13534_);
  and (_14132_, _14131_, _14129_);
  and (_14133_, _14115_, _13651_);
  or (_40966_, _14133_, _14132_);
  not (_14134_, _06070_);
  or (_14135_, _14134_, _14020_);
  or (_14136_, _14135_, _13538_);
  and (_14137_, _14113_, _13541_);
  or (_14138_, _14113_, _04931_);
  nand (_14139_, _14138_, _14135_);
  or (_14140_, _14139_, _14137_);
  and (_40967_, _14140_, _14136_);
  or (_14141_, _14113_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_14142_, _14141_, _14116_);
  or (_14143_, _14130_, _13549_);
  and (_14144_, _14143_, _14142_);
  and (_14145_, _14115_, _13863_);
  or (_40969_, _14145_, _14144_);
  nand (_14146_, _14118_, _13866_);
  or (_14147_, _14118_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_14148_, _14147_, _14116_);
  and (_14149_, _14148_, _14146_);
  and (_14150_, _14115_, _13871_);
  or (_40970_, _14150_, _14149_);
  or (_14151_, _14113_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_14152_, _14151_, _14116_);
  or (_14153_, _14130_, _13428_);
  and (_14154_, _14153_, _14152_);
  and (_14155_, _14115_, _13877_);
  or (_40971_, _14155_, _14154_);
  or (_14156_, _14113_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_14157_, _14156_, _14116_);
  or (_14158_, _14119_, _06854_);
  and (_14159_, _14158_, _14157_);
  and (_14160_, _14115_, _06878_);
  or (_40972_, _14160_, _14159_);
  not (_14161_, _04644_);
  or (_14162_, _14020_, _14161_);
  or (_14163_, _13520_, _14162_);
  and (_14164_, _12190_, _05209_);
  or (_14165_, _05209_, _04477_);
  nand (_14166_, _14165_, _14162_);
  or (_14167_, _14166_, _14164_);
  and (_40976_, _14167_, _14163_);
  or (_14168_, _12399_, _05236_);
  or (_14169_, _05235_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_14170_, _14169_, _05225_);
  and (_14171_, _14170_, _14168_);
  and (_14172_, _13637_, _05224_);
  or (_40977_, _14172_, _14171_);
  not (_14173_, _05209_);
  or (_14174_, _13534_, _14173_);
  or (_14175_, _05209_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_14176_, _14175_, _05225_);
  and (_14177_, _14176_, _14174_);
  and (_14178_, _13651_, _05224_);
  or (_40978_, _14178_, _14177_);
  or (_14179_, _13538_, _14162_);
  and (_14180_, _13541_, _05209_);
  or (_14181_, _05209_, _04929_);
  nand (_14182_, _14181_, _14162_);
  or (_14183_, _14182_, _14180_);
  and (_40979_, _14183_, _14179_);
  or (_14184_, _05209_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_14185_, _14184_, _05225_);
  or (_14186_, _13549_, _14173_);
  and (_14187_, _14186_, _14185_);
  and (_14188_, _13863_, _05224_);
  or (_40981_, _14188_, _14187_);
  nand (_14189_, _13866_, _05235_);
  or (_14190_, _05235_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_14191_, _14190_, _05225_);
  and (_14192_, _14191_, _14189_);
  and (_14193_, _13871_, _05224_);
  or (_40982_, _14193_, _14192_);
  or (_14194_, _05209_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_14195_, _14194_, _05225_);
  or (_14196_, _13428_, _14173_);
  and (_14197_, _14196_, _14195_);
  and (_14198_, _13877_, _05224_);
  or (_40983_, _14198_, _14197_);
  nor (_14199_, _43227_, _07467_);
  nor (_14200_, _05379_, _07467_);
  and (_14201_, _12145_, _05379_);
  or (_14202_, _14201_, _14200_);
  and (_14203_, _14202_, _03778_);
  nor (_14204_, _05744_, _06883_);
  or (_14205_, _14204_, _14200_);
  or (_14206_, _14205_, _04515_);
  and (_14207_, _05379_, \oc8051_golden_model_1.ACC [0]);
  or (_14208_, _14207_, _14200_);
  and (_14209_, _14208_, _04499_);
  nor (_14210_, _04499_, _07467_);
  or (_14211_, _14210_, _03599_);
  or (_14212_, _14211_, _14209_);
  and (_14213_, _14212_, _03516_);
  and (_14214_, _14213_, _14206_);
  and (_14215_, _12035_, _05992_);
  nor (_14216_, _05992_, _07467_);
  or (_14217_, _14216_, _14215_);
  and (_14218_, _14217_, _03515_);
  or (_14219_, _14218_, _14214_);
  and (_14220_, _14219_, _04524_);
  and (_14221_, _05379_, _04491_);
  or (_14222_, _14221_, _14200_);
  and (_14223_, _14222_, _03597_);
  or (_14224_, _14223_, _03603_);
  or (_14225_, _14224_, _14220_);
  or (_14226_, _14208_, _03611_);
  and (_14227_, _14226_, _03512_);
  and (_14228_, _14227_, _14225_);
  and (_14229_, _14200_, _03511_);
  or (_14230_, _14229_, _03504_);
  or (_14231_, _14230_, _14228_);
  or (_14232_, _14205_, _03505_);
  and (_14233_, _14232_, _14231_);
  or (_14234_, _14233_, _06919_);
  nor (_14235_, _07400_, _07398_);
  nor (_14236_, _14235_, _07401_);
  or (_14237_, _14236_, _06925_);
  and (_14238_, _14237_, _03501_);
  and (_14239_, _14238_, _14234_);
  nor (_14240_, _12066_, _07442_);
  or (_14241_, _14240_, _14216_);
  and (_14242_, _14241_, _03500_);
  or (_14243_, _14242_, _07441_);
  or (_14244_, _14243_, _14239_);
  or (_14245_, _14222_, _06889_);
  and (_14246_, _14245_, _05970_);
  and (_14247_, _14246_, _14244_);
  and (_14248_, _06836_, _05379_);
  or (_14249_, _14248_, _14200_);
  and (_14250_, _14249_, _05969_);
  or (_14251_, _14250_, _03644_);
  or (_14252_, _14251_, _14247_);
  nor (_14253_, _12129_, _06883_);
  or (_14254_, _14200_, _03275_);
  or (_14255_, _14254_, _14253_);
  and (_14256_, _14255_, _07805_);
  and (_14257_, _14256_, _14252_);
  nand (_14258_, _07803_, _03397_);
  or (_14259_, _07797_, _07772_);
  or (_14260_, _07803_, _14259_);
  and (_14261_, _14260_, _07455_);
  and (_14262_, _14261_, _14258_);
  or (_14263_, _14262_, _08861_);
  or (_14264_, _14263_, _14257_);
  and (_14265_, _12019_, _05379_);
  or (_14266_, _14200_, _04591_);
  or (_14267_, _14266_, _14265_);
  and (_14268_, _05379_, _06366_);
  or (_14269_, _14268_, _14200_);
  or (_14270_, _14269_, _04582_);
  and (_14271_, _14270_, _04589_);
  and (_14272_, _14271_, _14267_);
  and (_14273_, _14272_, _14264_);
  or (_14274_, _14273_, _14203_);
  and (_14275_, _14274_, _04596_);
  nand (_14276_, _14269_, _03655_);
  nor (_14277_, _14276_, _14204_);
  or (_14278_, _14277_, _14275_);
  and (_14279_, _14278_, _04594_);
  or (_14280_, _14200_, _05744_);
  and (_14281_, _14208_, _03773_);
  and (_14282_, _14281_, _14280_);
  or (_14283_, _14282_, _03653_);
  or (_14284_, _14283_, _14279_);
  nor (_14285_, _12017_, _06883_);
  or (_14286_, _14200_, _04608_);
  or (_14287_, _14286_, _14285_);
  and (_14288_, _14287_, _04606_);
  and (_14289_, _14288_, _14284_);
  nor (_14290_, _12015_, _06883_);
  or (_14291_, _14290_, _14200_);
  and (_14292_, _14291_, _03786_);
  or (_14293_, _14292_, _03809_);
  or (_14294_, _14293_, _14289_);
  or (_14295_, _14205_, _04260_);
  and (_14296_, _14295_, _03206_);
  and (_14297_, _14296_, _14294_);
  and (_14298_, _14200_, _03205_);
  or (_14299_, _14298_, _03816_);
  or (_14300_, _14299_, _14297_);
  or (_14301_, _14205_, _03820_);
  and (_14302_, _14301_, _43227_);
  and (_14303_, _14302_, _14300_);
  or (_14304_, _14303_, _14199_);
  and (_43424_, _14304_, _41991_);
  nor (_14305_, _43227_, _07461_);
  nor (_14306_, _05992_, _07461_);
  and (_14307_, _12224_, _05992_);
  or (_14308_, _14307_, _14306_);
  and (_14309_, _14308_, _03511_);
  nor (_14310_, _05379_, _07461_);
  and (_14311_, _05379_, _05898_);
  or (_14312_, _14311_, _14310_);
  or (_14313_, _14312_, _04524_);
  or (_14314_, _05379_, \oc8051_golden_model_1.B [1]);
  and (_14315_, _12234_, _05379_);
  not (_14316_, _14315_);
  and (_14317_, _14316_, _14314_);
  or (_14318_, _14317_, _04515_);
  nand (_14319_, _05379_, _03320_);
  and (_14320_, _14319_, _14314_);
  and (_14321_, _14320_, _04499_);
  nor (_14322_, _04499_, _07461_);
  or (_14323_, _14322_, _03599_);
  or (_14324_, _14323_, _14321_);
  and (_14325_, _14324_, _03516_);
  and (_14326_, _14325_, _14318_);
  and (_14327_, _12238_, _05992_);
  or (_14328_, _14327_, _14306_);
  and (_14329_, _14328_, _03515_);
  or (_14330_, _14329_, _03597_);
  or (_14331_, _14330_, _14326_);
  and (_14332_, _14331_, _14313_);
  or (_14333_, _14332_, _03603_);
  or (_14334_, _14320_, _03611_);
  and (_14335_, _14334_, _03512_);
  and (_14336_, _14335_, _14333_);
  or (_14337_, _14336_, _14309_);
  and (_14338_, _14337_, _03505_);
  and (_14339_, _14327_, _12253_);
  or (_14340_, _14339_, _14306_);
  and (_14341_, _14340_, _03504_);
  or (_14342_, _14341_, _06919_);
  or (_14343_, _14342_, _14338_);
  nor (_14344_, _07403_, _07346_);
  nor (_14345_, _14344_, _07404_);
  or (_14346_, _14345_, _06925_);
  and (_14347_, _14346_, _03501_);
  and (_14348_, _14347_, _14343_);
  nor (_14349_, _12270_, _07442_);
  or (_14350_, _14349_, _14306_);
  and (_14351_, _14350_, _03500_);
  or (_14352_, _14351_, _07441_);
  or (_14353_, _14352_, _14348_);
  or (_14354_, _14312_, _06889_);
  and (_14355_, _14354_, _14353_);
  or (_14356_, _14355_, _05969_);
  and (_14357_, _06835_, _05379_);
  or (_14358_, _14310_, _05970_);
  or (_14359_, _14358_, _14357_);
  and (_14360_, _14359_, _03275_);
  and (_14361_, _14360_, _14356_);
  nand (_14362_, _12330_, _05379_);
  and (_14363_, _14314_, _03644_);
  and (_14364_, _14363_, _14362_);
  or (_14365_, _14364_, _07455_);
  or (_14366_, _14365_, _14361_);
  nor (_14367_, _07798_, _07796_);
  or (_14368_, _14367_, _07799_);
  nor (_14369_, _14368_, _07803_);
  and (_14370_, _07803_, _07769_);
  or (_14371_, _14370_, _14369_);
  or (_14372_, _14371_, _07805_);
  and (_14373_, _14372_, _04582_);
  and (_14374_, _14373_, _14366_);
  nand (_14375_, _05379_, _04347_);
  and (_14376_, _14375_, _03650_);
  and (_14377_, _14376_, _14314_);
  or (_14378_, _14377_, _14374_);
  and (_14379_, _14378_, _04591_);
  or (_14380_, _12220_, _06883_);
  and (_14381_, _14314_, _03649_);
  and (_14382_, _14381_, _14380_);
  or (_14383_, _14382_, _14379_);
  and (_14384_, _14383_, _04589_);
  or (_14385_, _12347_, _06883_);
  and (_14386_, _14314_, _03778_);
  and (_14387_, _14386_, _14385_);
  or (_14388_, _14387_, _14384_);
  and (_14389_, _14388_, _04596_);
  or (_14390_, _12219_, _06883_);
  and (_14391_, _14314_, _03655_);
  and (_14392_, _14391_, _14390_);
  or (_14393_, _14392_, _14389_);
  and (_14394_, _14393_, _04594_);
  or (_14395_, _14310_, _05699_);
  and (_14396_, _14320_, _03773_);
  and (_14397_, _14396_, _14395_);
  or (_14398_, _14397_, _14394_);
  and (_14399_, _14398_, _03787_);
  or (_14400_, _14375_, _05699_);
  and (_14401_, _14314_, _03653_);
  and (_14402_, _14401_, _14400_);
  or (_14403_, _14319_, _05699_);
  and (_14404_, _14314_, _03786_);
  and (_14405_, _14404_, _14403_);
  or (_14406_, _14405_, _03809_);
  or (_14407_, _14406_, _14402_);
  or (_14408_, _14407_, _14399_);
  or (_14409_, _14317_, _04260_);
  and (_14410_, _14409_, _03206_);
  and (_14411_, _14410_, _14408_);
  and (_14412_, _14308_, _03205_);
  or (_14413_, _14412_, _03816_);
  or (_14414_, _14413_, _14411_);
  or (_14415_, _14310_, _03820_);
  or (_14416_, _14415_, _14315_);
  and (_14417_, _14416_, _43227_);
  and (_14418_, _14417_, _14414_);
  or (_14419_, _14418_, _14305_);
  and (_43425_, _14419_, _41991_);
  nor (_14420_, _43227_, _07475_);
  nor (_14421_, _05379_, _07475_);
  nor (_14422_, _06883_, _05130_);
  or (_14423_, _14422_, _14421_);
  or (_14424_, _14423_, _06889_);
  and (_14425_, _12416_, _05992_);
  and (_14426_, _14425_, _12447_);
  nor (_14427_, _05992_, _07475_);
  or (_14428_, _14427_, _03505_);
  or (_14429_, _14428_, _14426_);
  or (_14430_, _14423_, _04524_);
  nor (_14431_, _12430_, _06883_);
  or (_14432_, _14431_, _14421_);
  or (_14433_, _14432_, _04515_);
  and (_14434_, _05379_, \oc8051_golden_model_1.ACC [2]);
  or (_14435_, _14434_, _14421_);
  and (_14436_, _14435_, _04499_);
  nor (_14437_, _04499_, _07475_);
  or (_14438_, _14437_, _03599_);
  or (_14439_, _14438_, _14436_);
  and (_14440_, _14439_, _03516_);
  and (_14441_, _14440_, _14433_);
  or (_14442_, _14427_, _14425_);
  and (_14443_, _14442_, _03515_);
  or (_14444_, _14443_, _03597_);
  or (_14445_, _14444_, _14441_);
  and (_14446_, _14445_, _14430_);
  or (_14447_, _14446_, _03603_);
  or (_14448_, _14435_, _03611_);
  and (_14449_, _14448_, _03512_);
  and (_14450_, _14449_, _14447_);
  and (_14451_, _12414_, _05992_);
  or (_14452_, _14451_, _14427_);
  and (_14453_, _14452_, _03511_);
  or (_14454_, _14453_, _03504_);
  or (_14455_, _14454_, _14450_);
  and (_14456_, _14455_, _14429_);
  or (_14457_, _14456_, _06919_);
  nor (_14458_, _07406_, _07301_);
  nor (_14459_, _14458_, _07407_);
  or (_14460_, _14459_, _06925_);
  and (_14461_, _14460_, _03501_);
  and (_14462_, _14461_, _14457_);
  nor (_14463_, _12465_, _07442_);
  or (_14464_, _14463_, _14427_);
  and (_14465_, _14464_, _03500_);
  or (_14466_, _14465_, _07441_);
  or (_14467_, _14466_, _14462_);
  and (_14468_, _14467_, _14424_);
  or (_14469_, _14468_, _05969_);
  and (_14470_, _06839_, _05379_);
  or (_14471_, _14421_, _05970_);
  or (_14472_, _14471_, _14470_);
  and (_14473_, _14472_, _14469_);
  or (_14474_, _14473_, _03644_);
  nor (_14475_, _12524_, _06883_);
  or (_14476_, _14421_, _03275_);
  or (_14477_, _14476_, _14475_);
  and (_14478_, _14477_, _07805_);
  and (_14479_, _14478_, _14474_);
  not (_14480_, _07803_);
  or (_14481_, _14480_, _07759_);
  nor (_14482_, _07799_, _07770_);
  not (_14483_, _14482_);
  and (_14484_, _14483_, _07762_);
  nor (_14485_, _14483_, _07762_);
  nor (_14486_, _14485_, _14484_);
  or (_14487_, _14486_, _07803_);
  and (_14488_, _14487_, _07455_);
  and (_14489_, _14488_, _14481_);
  or (_14490_, _14489_, _08861_);
  or (_14491_, _14490_, _14479_);
  and (_14492_, _12538_, _05379_);
  or (_14493_, _14421_, _04591_);
  or (_14494_, _14493_, _14492_);
  and (_14495_, _05379_, _06414_);
  or (_14496_, _14495_, _14421_);
  or (_14497_, _14496_, _04582_);
  and (_14498_, _14497_, _04589_);
  and (_14499_, _14498_, _14494_);
  and (_14500_, _14499_, _14491_);
  and (_14501_, _12544_, _05379_);
  or (_14502_, _14501_, _14421_);
  and (_14503_, _14502_, _03778_);
  or (_14504_, _14503_, _14500_);
  and (_14505_, _14504_, _04596_);
  or (_14506_, _14421_, _05793_);
  and (_14507_, _14496_, _03655_);
  and (_14508_, _14507_, _14506_);
  or (_14509_, _14508_, _14505_);
  and (_14510_, _14509_, _04594_);
  and (_14511_, _14435_, _03773_);
  and (_14512_, _14511_, _14506_);
  or (_14513_, _14512_, _03653_);
  or (_14514_, _14513_, _14510_);
  nor (_14515_, _12537_, _06883_);
  or (_14516_, _14421_, _04608_);
  or (_14517_, _14516_, _14515_);
  and (_14518_, _14517_, _04606_);
  and (_14519_, _14518_, _14514_);
  nor (_14520_, _12543_, _06883_);
  or (_14521_, _14520_, _14421_);
  and (_14522_, _14521_, _03786_);
  or (_14523_, _14522_, _03809_);
  or (_14524_, _14523_, _14519_);
  or (_14525_, _14432_, _04260_);
  and (_14526_, _14525_, _03206_);
  and (_14527_, _14526_, _14524_);
  and (_14528_, _14452_, _03205_);
  or (_14529_, _14528_, _03816_);
  or (_14530_, _14529_, _14527_);
  and (_14531_, _12600_, _05379_);
  or (_14532_, _14421_, _03820_);
  or (_14533_, _14532_, _14531_);
  and (_14534_, _14533_, _43227_);
  and (_14535_, _14534_, _14530_);
  or (_14536_, _14535_, _14420_);
  and (_43426_, _14536_, _41991_);
  nor (_14537_, _43227_, _07476_);
  nor (_14538_, _05379_, _07476_);
  nor (_14539_, _12731_, _06883_);
  or (_14540_, _14539_, _14538_);
  and (_14541_, _14540_, _03644_);
  nor (_14542_, _05992_, _07476_);
  and (_14543_, _12638_, _05992_);
  or (_14544_, _14543_, _14542_);
  or (_14545_, _14542_, _12653_);
  and (_14546_, _14545_, _14544_);
  or (_14547_, _14546_, _03505_);
  nor (_14548_, _12625_, _06883_);
  or (_14549_, _14548_, _14538_);
  or (_14550_, _14549_, _04515_);
  and (_14551_, _05379_, \oc8051_golden_model_1.ACC [3]);
  or (_14552_, _14551_, _14538_);
  and (_14553_, _14552_, _04499_);
  nor (_14554_, _04499_, _07476_);
  or (_14555_, _14554_, _03599_);
  or (_14556_, _14555_, _14553_);
  and (_14557_, _14556_, _03516_);
  and (_14558_, _14557_, _14550_);
  and (_14559_, _14544_, _03515_);
  or (_14560_, _14559_, _03597_);
  or (_14561_, _14560_, _14558_);
  nor (_14562_, _06883_, _04944_);
  or (_14563_, _14562_, _14538_);
  or (_14564_, _14563_, _04524_);
  and (_14565_, _14564_, _14561_);
  or (_14566_, _14565_, _03603_);
  or (_14567_, _14552_, _03611_);
  and (_14568_, _14567_, _03512_);
  and (_14569_, _14568_, _14566_);
  and (_14570_, _12622_, _05992_);
  or (_14571_, _14570_, _14542_);
  and (_14572_, _14571_, _03511_);
  or (_14573_, _14572_, _03504_);
  or (_14574_, _14573_, _14569_);
  and (_14575_, _14574_, _14547_);
  or (_14576_, _14575_, _06919_);
  nor (_14577_, _07409_, _07243_);
  nor (_14578_, _14577_, _07410_);
  or (_14579_, _14578_, _06925_);
  and (_14580_, _14579_, _03501_);
  and (_14581_, _14580_, _14576_);
  nor (_14582_, _12671_, _07442_);
  or (_14583_, _14582_, _14542_);
  and (_14584_, _14583_, _03500_);
  or (_14585_, _14584_, _07441_);
  or (_14586_, _14585_, _14581_);
  or (_14587_, _14563_, _06889_);
  and (_14588_, _14587_, _14586_);
  or (_14589_, _14588_, _05969_);
  and (_14590_, _06838_, _05379_);
  or (_14591_, _14538_, _05970_);
  or (_14592_, _14591_, _14590_);
  and (_14593_, _14592_, _03275_);
  and (_14594_, _14593_, _14589_);
  or (_14595_, _14594_, _14541_);
  and (_14596_, _14595_, _07805_);
  nor (_14597_, _14484_, _07761_);
  nor (_14598_, _14597_, _07754_);
  and (_14599_, _14597_, _07754_);
  or (_14600_, _14599_, _14598_);
  or (_14601_, _14600_, _07803_);
  or (_14602_, _14480_, _07751_);
  and (_14603_, _14602_, _07455_);
  and (_14604_, _14603_, _14601_);
  or (_14605_, _14604_, _08861_);
  or (_14606_, _14605_, _14596_);
  and (_14607_, _12746_, _05379_);
  or (_14608_, _14538_, _04591_);
  or (_14609_, _14608_, _14607_);
  and (_14610_, _05379_, _06347_);
  or (_14611_, _14610_, _14538_);
  or (_14612_, _14611_, _04582_);
  and (_14613_, _14612_, _04589_);
  and (_14614_, _14613_, _14609_);
  and (_14615_, _14614_, _14606_);
  and (_14616_, _12619_, _05379_);
  or (_14617_, _14616_, _14538_);
  and (_14618_, _14617_, _03778_);
  or (_14619_, _14618_, _14615_);
  and (_14620_, _14619_, _04596_);
  or (_14621_, _14538_, _05650_);
  and (_14622_, _14611_, _03655_);
  and (_14623_, _14622_, _14621_);
  or (_14624_, _14623_, _14620_);
  and (_14625_, _14624_, _04594_);
  and (_14626_, _14552_, _03773_);
  and (_14627_, _14626_, _14621_);
  or (_14628_, _14627_, _03653_);
  or (_14629_, _14628_, _14625_);
  nor (_14630_, _12745_, _06883_);
  or (_14631_, _14538_, _04608_);
  or (_14632_, _14631_, _14630_);
  and (_14633_, _14632_, _04606_);
  and (_14634_, _14633_, _14629_);
  nor (_14635_, _12618_, _06883_);
  or (_14636_, _14635_, _14538_);
  and (_14637_, _14636_, _03786_);
  or (_14638_, _14637_, _03809_);
  or (_14639_, _14638_, _14634_);
  or (_14640_, _14549_, _04260_);
  and (_14641_, _14640_, _03206_);
  and (_14642_, _14641_, _14639_);
  and (_14643_, _14571_, _03205_);
  or (_14644_, _14643_, _03816_);
  or (_14645_, _14644_, _14642_);
  and (_14646_, _12806_, _05379_);
  or (_14647_, _14538_, _03820_);
  or (_14648_, _14647_, _14646_);
  and (_14649_, _14648_, _43227_);
  and (_14650_, _14649_, _14645_);
  or (_14651_, _14650_, _14537_);
  and (_43428_, _14651_, _41991_);
  nor (_14652_, _43227_, _07477_);
  nor (_14653_, _05379_, _07477_);
  nor (_14654_, _12936_, _06883_);
  or (_14655_, _14654_, _14653_);
  and (_14656_, _14655_, _03644_);
  nor (_14657_, _05840_, _06883_);
  or (_14658_, _14657_, _14653_);
  or (_14659_, _14658_, _06889_);
  nor (_14660_, _05992_, _07477_);
  and (_14661_, _12853_, _05992_);
  or (_14662_, _14661_, _14660_);
  and (_14663_, _14662_, _03511_);
  nor (_14664_, _12820_, _06883_);
  or (_14665_, _14664_, _14653_);
  or (_14666_, _14665_, _04515_);
  and (_14667_, _05379_, \oc8051_golden_model_1.ACC [4]);
  or (_14668_, _14667_, _14653_);
  and (_14669_, _14668_, _04499_);
  nor (_14670_, _04499_, _07477_);
  or (_14671_, _14670_, _03599_);
  or (_14672_, _14671_, _14669_);
  and (_14673_, _14672_, _03516_);
  and (_14674_, _14673_, _14666_);
  and (_14675_, _12830_, _05992_);
  or (_14676_, _14675_, _14660_);
  and (_14677_, _14676_, _03515_);
  or (_14678_, _14677_, _03597_);
  or (_14679_, _14678_, _14674_);
  or (_14680_, _14658_, _04524_);
  and (_14681_, _14680_, _14679_);
  or (_14682_, _14681_, _03603_);
  or (_14683_, _14668_, _03611_);
  and (_14684_, _14683_, _03512_);
  and (_14685_, _14684_, _14682_);
  or (_14686_, _14685_, _14663_);
  and (_14687_, _14686_, _03505_);
  or (_14688_, _14660_, _12860_);
  and (_14689_, _14688_, _03504_);
  and (_14690_, _14689_, _14676_);
  or (_14691_, _14690_, _06919_);
  or (_14692_, _14691_, _14687_);
  nor (_14693_, _07414_, _07412_);
  nor (_14694_, _14693_, _07415_);
  or (_14695_, _14694_, _06925_);
  and (_14696_, _14695_, _03501_);
  and (_14697_, _14696_, _14692_);
  nor (_14698_, _12828_, _07442_);
  or (_14699_, _14698_, _14660_);
  and (_14700_, _14699_, _03500_);
  or (_14701_, _14700_, _07441_);
  or (_14702_, _14701_, _14697_);
  and (_14703_, _14702_, _14659_);
  or (_14704_, _14703_, _05969_);
  and (_14705_, _06843_, _05379_);
  or (_14706_, _14653_, _05970_);
  or (_14707_, _14706_, _14705_);
  and (_14708_, _14707_, _03275_);
  and (_14709_, _14708_, _14704_);
  or (_14710_, _14709_, _14656_);
  and (_14711_, _14710_, _07805_);
  or (_14712_, _14480_, _07743_);
  nor (_14713_, _14597_, _07753_);
  or (_14714_, _14713_, _07752_);
  nand (_14715_, _14714_, _07791_);
  or (_14716_, _14714_, _07791_);
  and (_14717_, _14716_, _14715_);
  or (_14718_, _14717_, _07803_);
  and (_14719_, _14718_, _07455_);
  and (_14720_, _14719_, _14712_);
  or (_14721_, _14720_, _08861_);
  or (_14722_, _14721_, _14711_);
  and (_14723_, _12951_, _05379_);
  or (_14724_, _14653_, _04591_);
  or (_14725_, _14724_, _14723_);
  and (_14726_, _06375_, _05379_);
  or (_14727_, _14726_, _14653_);
  or (_14728_, _14727_, _04582_);
  and (_14729_, _14728_, _04589_);
  and (_14730_, _14729_, _14725_);
  and (_14731_, _14730_, _14722_);
  and (_14732_, _12957_, _05379_);
  or (_14733_, _14732_, _14653_);
  and (_14734_, _14733_, _03778_);
  or (_14735_, _14734_, _14731_);
  and (_14736_, _14735_, _04596_);
  or (_14737_, _14653_, _05889_);
  and (_14738_, _14727_, _03655_);
  and (_14739_, _14738_, _14737_);
  or (_14740_, _14739_, _14736_);
  and (_14741_, _14740_, _04594_);
  and (_14742_, _14668_, _03773_);
  and (_14743_, _14742_, _14737_);
  or (_14744_, _14743_, _03653_);
  or (_14745_, _14744_, _14741_);
  nor (_14746_, _12949_, _06883_);
  or (_14747_, _14653_, _04608_);
  or (_14748_, _14747_, _14746_);
  and (_14749_, _14748_, _04606_);
  and (_14750_, _14749_, _14745_);
  nor (_14751_, _12956_, _06883_);
  or (_14752_, _14751_, _14653_);
  and (_14753_, _14752_, _03786_);
  or (_14754_, _14753_, _03809_);
  or (_14755_, _14754_, _14750_);
  or (_14756_, _14665_, _04260_);
  and (_14757_, _14756_, _03206_);
  and (_14758_, _14757_, _14755_);
  and (_14759_, _14662_, _03205_);
  or (_14760_, _14759_, _03816_);
  or (_14761_, _14760_, _14758_);
  and (_14762_, _13013_, _05379_);
  or (_14763_, _14653_, _03820_);
  or (_14764_, _14763_, _14762_);
  and (_14765_, _14764_, _43227_);
  and (_14766_, _14765_, _14761_);
  or (_14767_, _14766_, _14652_);
  and (_43429_, _14767_, _41991_);
  nor (_14768_, _43227_, _07478_);
  nor (_14769_, _05379_, _07478_);
  nor (_14770_, _13139_, _06883_);
  or (_14771_, _14770_, _14769_);
  and (_14772_, _14771_, _03644_);
  nor (_14773_, _05552_, _06883_);
  or (_14774_, _14773_, _14769_);
  or (_14775_, _14774_, _06889_);
  nor (_14776_, _05992_, _07478_);
  and (_14777_, _13032_, _05992_);
  or (_14778_, _14777_, _14776_);
  and (_14779_, _14778_, _03511_);
  nor (_14780_, _13035_, _06883_);
  or (_14781_, _14780_, _14769_);
  or (_14782_, _14781_, _04515_);
  and (_14783_, _05379_, \oc8051_golden_model_1.ACC [5]);
  or (_14784_, _14783_, _14769_);
  and (_14785_, _14784_, _04499_);
  nor (_14786_, _04499_, _07478_);
  or (_14787_, _14786_, _03599_);
  or (_14788_, _14787_, _14785_);
  and (_14789_, _14788_, _03516_);
  and (_14790_, _14789_, _14782_);
  and (_14791_, _13051_, _05992_);
  or (_14792_, _14791_, _14776_);
  and (_14793_, _14792_, _03515_);
  or (_14794_, _14793_, _03597_);
  or (_14795_, _14794_, _14790_);
  or (_14796_, _14774_, _04524_);
  and (_14797_, _14796_, _14795_);
  or (_14798_, _14797_, _03603_);
  or (_14799_, _14784_, _03611_);
  and (_14800_, _14799_, _03512_);
  and (_14801_, _14800_, _14798_);
  or (_14802_, _14801_, _14779_);
  and (_14803_, _14802_, _03505_);
  or (_14804_, _14776_, _13066_);
  and (_14805_, _14804_, _03504_);
  and (_14806_, _14805_, _14792_);
  or (_14807_, _14806_, _06919_);
  or (_14808_, _14807_, _14803_);
  or (_14809_, _07116_, _07117_);
  and (_14810_, _14809_, _07416_);
  nor (_14811_, _14810_, _07417_);
  or (_14812_, _14811_, _06925_);
  and (_14813_, _14812_, _03501_);
  and (_14814_, _14813_, _14808_);
  nor (_14815_, _13030_, _07442_);
  or (_14816_, _14815_, _14776_);
  and (_14817_, _14816_, _03500_);
  or (_14818_, _14817_, _07441_);
  or (_14819_, _14818_, _14814_);
  and (_14820_, _14819_, _14775_);
  or (_14821_, _14820_, _05969_);
  and (_14822_, _06842_, _05379_);
  or (_14823_, _14769_, _05970_);
  or (_14824_, _14823_, _14822_);
  and (_14825_, _14824_, _03275_);
  and (_14826_, _14825_, _14821_);
  or (_14827_, _14826_, _14772_);
  and (_14828_, _14827_, _07805_);
  not (_14829_, _07781_);
  and (_14830_, _14715_, _14829_);
  nor (_14831_, _14830_, _07790_);
  and (_14832_, _14830_, _07790_);
  or (_14833_, _14832_, _14831_);
  nor (_14834_, _07803_, _07805_);
  and (_14835_, _14834_, _14833_);
  and (_14836_, _07735_, _07455_);
  and (_14837_, _14836_, _07803_);
  or (_14838_, _14837_, _08861_);
  or (_14839_, _14838_, _14835_);
  or (_14840_, _14839_, _14828_);
  and (_14841_, _13154_, _05379_);
  or (_14842_, _14769_, _04591_);
  or (_14843_, _14842_, _14841_);
  and (_14844_, _06358_, _05379_);
  or (_14845_, _14844_, _14769_);
  or (_14846_, _14845_, _04582_);
  and (_14847_, _14846_, _04589_);
  and (_14848_, _14847_, _14843_);
  and (_14849_, _14848_, _14840_);
  and (_14850_, _13160_, _05379_);
  or (_14851_, _14850_, _14769_);
  and (_14852_, _14851_, _03778_);
  or (_14853_, _14852_, _14849_);
  and (_14854_, _14853_, _04596_);
  or (_14855_, _14769_, _05601_);
  and (_14856_, _14845_, _03655_);
  and (_14857_, _14856_, _14855_);
  or (_14858_, _14857_, _14854_);
  and (_14859_, _14858_, _04594_);
  and (_14860_, _14784_, _03773_);
  and (_14861_, _14860_, _14855_);
  or (_14862_, _14861_, _03653_);
  or (_14863_, _14862_, _14859_);
  nor (_14864_, _13152_, _06883_);
  or (_14865_, _14769_, _04608_);
  or (_14866_, _14865_, _14864_);
  and (_14867_, _14866_, _04606_);
  and (_14868_, _14867_, _14863_);
  nor (_14869_, _13159_, _06883_);
  or (_14870_, _14869_, _14769_);
  and (_14871_, _14870_, _03786_);
  or (_14872_, _14871_, _03809_);
  or (_14873_, _14872_, _14868_);
  or (_14874_, _14781_, _04260_);
  and (_14875_, _14874_, _03206_);
  and (_14876_, _14875_, _14873_);
  and (_14877_, _14778_, _03205_);
  or (_14878_, _14877_, _03816_);
  or (_14879_, _14878_, _14876_);
  and (_14880_, _13217_, _05379_);
  or (_14881_, _14769_, _03820_);
  or (_14882_, _14881_, _14880_);
  and (_14883_, _14882_, _43227_);
  and (_14884_, _14883_, _14879_);
  or (_14885_, _14884_, _14768_);
  and (_43430_, _14885_, _41991_);
  nor (_14886_, _43227_, _07720_);
  nor (_14887_, _05379_, _07720_);
  nor (_14888_, _13356_, _06883_);
  or (_14889_, _14888_, _14887_);
  and (_14890_, _14889_, _03644_);
  nor (_14891_, _05442_, _06883_);
  or (_14892_, _14891_, _14887_);
  or (_14893_, _14892_, _06889_);
  nor (_14894_, _05992_, _07720_);
  and (_14895_, _13251_, _05992_);
  or (_14896_, _14895_, _14894_);
  and (_14897_, _14896_, _03511_);
  nor (_14898_, _13235_, _06883_);
  or (_14899_, _14898_, _14887_);
  or (_14900_, _14899_, _04515_);
  and (_14901_, _05379_, \oc8051_golden_model_1.ACC [6]);
  or (_14902_, _14901_, _14887_);
  and (_14903_, _14902_, _04499_);
  nor (_14904_, _04499_, _07720_);
  or (_14905_, _14904_, _03599_);
  or (_14906_, _14905_, _14903_);
  and (_14907_, _14906_, _03516_);
  and (_14908_, _14907_, _14900_);
  and (_14909_, _13266_, _05992_);
  or (_14910_, _14909_, _14894_);
  and (_14911_, _14910_, _03515_);
  or (_14912_, _14911_, _03597_);
  or (_14913_, _14912_, _14908_);
  or (_14914_, _14892_, _04524_);
  and (_14915_, _14914_, _14913_);
  or (_14916_, _14915_, _03603_);
  or (_14917_, _14902_, _03611_);
  and (_14918_, _14917_, _03512_);
  and (_14919_, _14918_, _14916_);
  or (_14920_, _14919_, _14897_);
  and (_14921_, _14920_, _03505_);
  or (_14922_, _14894_, _13281_);
  and (_14923_, _14922_, _03504_);
  and (_14924_, _14923_, _14910_);
  or (_14925_, _14924_, _06919_);
  or (_14926_, _14925_, _14921_);
  nor (_14927_, _07430_, _07418_);
  nor (_14928_, _14927_, _07431_);
  or (_14929_, _14928_, _06925_);
  and (_14930_, _14929_, _03501_);
  and (_14931_, _14930_, _14926_);
  nor (_14932_, _13249_, _07442_);
  or (_14933_, _14932_, _14894_);
  and (_14934_, _14933_, _03500_);
  or (_14935_, _14934_, _07441_);
  or (_14936_, _14935_, _14931_);
  and (_14937_, _14936_, _14893_);
  or (_14938_, _14937_, _05969_);
  and (_14939_, _06531_, _05379_);
  or (_14940_, _14887_, _05970_);
  or (_14941_, _14940_, _14939_);
  and (_14942_, _14941_, _03275_);
  and (_14943_, _14942_, _14938_);
  or (_14944_, _14943_, _14890_);
  and (_14945_, _14944_, _07805_);
  nor (_14946_, _14830_, _07736_);
  or (_14947_, _14946_, _07737_);
  or (_14948_, _14947_, _07793_);
  nand (_14949_, _14947_, _07793_);
  and (_14950_, _14949_, _14948_);
  or (_14951_, _14950_, _07803_);
  and (_14952_, _07726_, _07455_);
  or (_14953_, _14952_, _14834_);
  and (_14954_, _14953_, _14951_);
  or (_14955_, _14954_, _08861_);
  or (_14956_, _14955_, _14945_);
  and (_14957_, _13245_, _05379_);
  or (_14958_, _14887_, _04591_);
  or (_14959_, _14958_, _14957_);
  and (_14960_, _13363_, _05379_);
  or (_14961_, _14960_, _14887_);
  or (_14962_, _14961_, _04582_);
  and (_14963_, _14962_, _04589_);
  and (_14964_, _14963_, _14959_);
  and (_14965_, _14964_, _14956_);
  and (_14966_, _13374_, _05379_);
  or (_14967_, _14966_, _14887_);
  and (_14968_, _14967_, _03778_);
  or (_14969_, _14968_, _14965_);
  and (_14970_, _14969_, _04596_);
  or (_14971_, _14887_, _05491_);
  and (_14972_, _14961_, _03655_);
  and (_14973_, _14972_, _14971_);
  or (_14974_, _14973_, _14970_);
  and (_14975_, _14974_, _04594_);
  and (_14976_, _14902_, _03773_);
  and (_14977_, _14976_, _14971_);
  or (_14978_, _14977_, _03653_);
  or (_14979_, _14978_, _14975_);
  nor (_14980_, _13243_, _06883_);
  or (_14981_, _14887_, _04608_);
  or (_14982_, _14981_, _14980_);
  and (_14983_, _14982_, _04606_);
  and (_14984_, _14983_, _14979_);
  nor (_14985_, _13373_, _06883_);
  or (_14986_, _14985_, _14887_);
  and (_14987_, _14986_, _03786_);
  or (_14988_, _14987_, _03809_);
  or (_14989_, _14988_, _14984_);
  or (_14990_, _14899_, _04260_);
  and (_14991_, _14990_, _03206_);
  and (_14992_, _14991_, _14989_);
  and (_14993_, _14896_, _03205_);
  or (_14994_, _14993_, _03816_);
  or (_14995_, _14994_, _14992_);
  and (_14996_, _13425_, _05379_);
  or (_14997_, _14887_, _03820_);
  or (_14998_, _14997_, _14996_);
  and (_14999_, _14998_, _43227_);
  and (_15000_, _14999_, _14995_);
  or (_15001_, _15000_, _14886_);
  and (_43431_, _15001_, _41991_);
  nor (_15002_, _43227_, _03397_);
  and (_15003_, _08814_, \oc8051_golden_model_1.ACC [1]);
  nand (_15004_, _08769_, _06061_);
  and (_15005_, _06622_, _03397_);
  nor (_15006_, _08701_, _15005_);
  or (_15007_, _10369_, _15006_);
  nand (_15008_, _08524_, _10129_);
  not (_15009_, _03954_);
  nor (_15010_, _05744_, _07957_);
  nor (_15011_, _05371_, _03397_);
  and (_15012_, _05371_, _06366_);
  nor (_15013_, _15012_, _15011_);
  nor (_15014_, _15013_, _15010_);
  and (_15015_, _15014_, _03655_);
  and (_15016_, _12019_, _05371_);
  nor (_15017_, _15016_, _15011_);
  nand (_15018_, _15017_, _03649_);
  or (_15019_, _12145_, _03777_);
  and (_15020_, _15019_, _08473_);
  nand (_15021_, _04042_, _03313_);
  nor (_15022_, _12129_, _07957_);
  nor (_15023_, _15022_, _15011_);
  nor (_15024_, _15023_, _03275_);
  and (_15025_, _05371_, _04491_);
  nor (_15026_, _15025_, _15011_);
  nand (_15027_, _15026_, _07441_);
  nand (_15028_, _08032_, _08021_);
  or (_15029_, _08041_, _04491_);
  or (_15030_, _08048_, _04491_);
  nor (_15031_, _04063_, _03397_);
  and (_15032_, _04063_, _03397_);
  nor (_15033_, _15032_, _15031_);
  nand (_15034_, _15033_, _08048_);
  and (_15035_, _15034_, _08052_);
  and (_15036_, _15035_, _15030_);
  and (_15037_, _15036_, _06068_);
  or (_15038_, _15037_, _06836_);
  or (_15039_, _15036_, _08051_);
  and (_15040_, _15039_, _03262_);
  or (_15041_, _15040_, _04509_);
  and (_15042_, _15041_, _04515_);
  and (_15043_, _15042_, _15038_);
  nor (_15044_, _15011_, _15010_);
  nor (_15045_, _15044_, _04515_);
  or (_15046_, _15045_, _03515_);
  or (_15047_, _15046_, _15043_);
  nor (_15048_, _05983_, _03397_);
  and (_15049_, _12035_, _05983_);
  nor (_15050_, _15049_, _15048_);
  nand (_15051_, _15050_, _03515_);
  and (_15052_, _15051_, _04524_);
  and (_15053_, _15052_, _15047_);
  nor (_15054_, _15026_, _04524_);
  or (_15055_, _15054_, _08042_);
  or (_15056_, _15055_, _15053_);
  and (_15057_, _15056_, _15029_);
  or (_15058_, _15057_, _04529_);
  or (_15059_, _06836_, _08102_);
  and (_15060_, _15059_, _03611_);
  and (_15061_, _15060_, _15058_);
  nor (_15062_, _08238_, _03611_);
  or (_15063_, _15062_, _08106_);
  or (_15064_, _15063_, _15061_);
  nand (_15065_, _08106_, _07536_);
  and (_15066_, _15065_, _15064_);
  or (_15067_, _15066_, _03511_);
  or (_15068_, _15011_, _03512_);
  and (_15069_, _15068_, _03505_);
  and (_15070_, _15069_, _15067_);
  nor (_15071_, _15044_, _03505_);
  or (_15072_, _15071_, _06919_);
  or (_15073_, _15072_, _15070_);
  not (_15074_, _07379_);
  nand (_15075_, _15074_, _06919_);
  and (_15076_, _15075_, _15073_);
  or (_15077_, _15076_, _08034_);
  nor (_15078_, _08144_, _08036_);
  or (_15079_, _15078_, _08037_);
  and (_15080_, _15079_, _15077_);
  not (_15081_, _08144_);
  and (_15082_, _15081_, _08036_);
  or (_15083_, _15082_, _08032_);
  or (_15084_, _15083_, _15080_);
  and (_15085_, _15084_, _15028_);
  or (_15086_, _15085_, _03635_);
  nor (_15087_, _08313_, _03397_);
  nor (_15088_, _15087_, _08314_);
  nand (_15089_, _15088_, _03635_);
  and (_15090_, _15089_, _08161_);
  and (_15091_, _15090_, _15086_);
  nor (_15092_, _08380_, _08161_);
  or (_15093_, _15092_, _03371_);
  or (_15094_, _15093_, _15091_);
  nand (_15095_, _04042_, _03371_);
  and (_15096_, _15095_, _03501_);
  and (_15097_, _15096_, _15094_);
  nor (_15098_, _12066_, _08421_);
  nor (_15099_, _15098_, _15048_);
  nor (_15100_, _15099_, _03501_);
  or (_15101_, _15100_, _07441_);
  or (_15102_, _15101_, _15097_);
  and (_15103_, _15102_, _15027_);
  or (_15104_, _15103_, _05969_);
  and (_15105_, _06836_, _05371_);
  nor (_15106_, _15105_, _15011_);
  nand (_15107_, _15106_, _05969_);
  and (_15108_, _15107_, _03275_);
  and (_15109_, _15108_, _15104_);
  or (_15110_, _15109_, _15024_);
  and (_15111_, _15110_, _07805_);
  or (_15112_, _14834_, _03313_);
  or (_15113_, _15112_, _15111_);
  and (_15114_, _15113_, _15021_);
  or (_15115_, _15114_, _03650_);
  nand (_15116_, _15013_, _03650_);
  and (_15117_, _15116_, _08446_);
  and (_15118_, _15117_, _15115_);
  nor (_15119_, _08446_, _04042_);
  or (_15120_, _15119_, _08451_);
  or (_15121_, _15120_, _15118_);
  and (_15122_, _04510_, _03397_);
  nor (_15123_, _15122_, _08660_);
  not (_15124_, _11837_);
  and (_15125_, _15124_, _15123_);
  or (_15126_, _15125_, _11838_);
  and (_15127_, _15126_, _15121_);
  and (_15128_, _11837_, _15123_);
  or (_15129_, _15128_, _11839_);
  or (_15130_, _15129_, _15127_);
  and (_15131_, _03680_, _03230_);
  not (_15132_, _11839_);
  nor (_15133_, _15132_, _15123_);
  nor (_15134_, _15133_, _15131_);
  and (_15135_, _15134_, _15130_);
  and (_15136_, _15131_, _15006_);
  or (_15137_, _15136_, _15135_);
  and (_15138_, _15137_, _04185_);
  and (_15139_, _15006_, _04184_);
  or (_15140_, _15139_, _03776_);
  or (_15141_, _15140_, _15138_);
  and (_15142_, _15141_, _15020_);
  and (_15143_, _08472_, _10130_);
  or (_15144_, _15143_, _03649_);
  or (_15145_, _15144_, _15142_);
  and (_15146_, _15145_, _15018_);
  or (_15147_, _15146_, _03778_);
  or (_15148_, _15011_, _04589_);
  and (_15149_, _03237_, _03134_);
  not (_15150_, _15149_);
  and (_15151_, _15150_, _15148_);
  and (_15152_, _15151_, _15147_);
  and (_15153_, _15149_, _08660_);
  or (_15154_, _15153_, _04198_);
  or (_15155_, _15154_, _15152_);
  or (_15156_, _08701_, _07944_);
  and (_15157_, _15156_, _03772_);
  and (_15158_, _15157_, _15155_);
  or (_15159_, _12144_, _07942_);
  and (_15160_, _15159_, _11368_);
  or (_15161_, _15160_, _15158_);
  or (_15162_, _08787_, _08500_);
  and (_15163_, _15162_, _04596_);
  and (_15164_, _15163_, _15161_);
  or (_15165_, _15164_, _15015_);
  and (_15166_, _15165_, _15009_);
  nor (_15167_, _15122_, _15009_);
  or (_15168_, _15167_, _15166_);
  and (_15169_, _03567_, _03235_);
  not (_15170_, _15169_);
  and (_15171_, _15170_, _15168_);
  nor (_15172_, _15170_, _15122_);
  or (_15173_, _15172_, _04207_);
  or (_15174_, _15173_, _15171_);
  nand (_15175_, _15005_, _04207_);
  and (_15176_, _15175_, _03785_);
  and (_15177_, _15176_, _15174_);
  nand (_15178_, _12015_, _08525_);
  and (_15179_, _15178_, _11358_);
  or (_15180_, _15179_, _15177_);
  and (_15181_, _15180_, _15008_);
  or (_15182_, _15181_, _03653_);
  nor (_15183_, _12017_, _07957_);
  nor (_15184_, _15183_, _15011_);
  nand (_15185_, _15184_, _03653_);
  and (_15186_, _15185_, _07933_);
  and (_15187_, _15186_, _15182_);
  nor (_15188_, _08144_, _07933_);
  or (_15189_, _15188_, _08539_);
  or (_15190_, _15189_, _15187_);
  nand (_15191_, _08539_, _08021_);
  and (_15192_, _15191_, _15190_);
  or (_15193_, _15192_, _03782_);
  nand (_15194_, _15088_, _03782_);
  and (_15195_, _15194_, _08602_);
  and (_15196_, _15195_, _15193_);
  nor (_15197_, _08602_, _08380_);
  or (_15198_, _15197_, _08600_);
  or (_15199_, _15198_, _15196_);
  nand (_15200_, _08600_, _07911_);
  and (_15201_, _15200_, _09696_);
  and (_15202_, _15201_, _15199_);
  and (_15203_, _10362_, _15123_);
  or (_15204_, _15203_, _08679_);
  or (_15205_, _15204_, _15202_);
  and (_15206_, _15205_, _15007_);
  or (_15207_, _15206_, _03524_);
  nand (_15208_, _09943_, _03524_);
  and (_15209_, _15208_, _08771_);
  and (_15210_, _15209_, _15207_);
  and (_15211_, _08720_, _10130_);
  or (_15212_, _15211_, _08769_);
  or (_15213_, _15212_, _15210_);
  and (_15214_, _15213_, _15004_);
  or (_15215_, _15214_, _03809_);
  nand (_15216_, _15044_, _03809_);
  and (_15217_, _15216_, _08810_);
  and (_15218_, _15217_, _15215_);
  and (_15219_, _08809_, _03397_);
  or (_15220_, _15219_, _15218_);
  and (_15221_, _15220_, _09690_);
  or (_15222_, _15221_, _15003_);
  and (_15223_, _15222_, _03206_);
  and (_15224_, _15011_, _03205_);
  or (_15225_, _15224_, _03816_);
  or (_15226_, _15225_, _15223_);
  nand (_15227_, _15044_, _03816_);
  and (_15228_, _15227_, _08832_);
  and (_15229_, _15228_, _15226_);
  nor (_15230_, _08838_, _03397_);
  nor (_15231_, _15230_, _11974_);
  or (_15232_, _15231_, _15229_);
  nand (_15233_, _08838_, _03320_);
  and (_15234_, _15233_, _43227_);
  and (_15235_, _15234_, _15232_);
  or (_15236_, _15235_, _15002_);
  and (_43433_, _15236_, _41991_);
  nor (_15237_, _43227_, _03320_);
  nand (_15238_, _08600_, _03397_);
  nand (_15239_, _08524_, _08382_);
  nor (_15240_, _05371_, _03320_);
  and (_15241_, _12219_, _05371_);
  nor (_15242_, _15241_, _15240_);
  nor (_15243_, _15242_, _04596_);
  and (_15244_, _12220_, _05371_);
  nor (_15245_, _15244_, _15240_);
  nand (_15246_, _15245_, _03649_);
  nand (_15247_, _04434_, _03313_);
  and (_15248_, _05371_, _05898_);
  nor (_15249_, _15248_, _15240_);
  nand (_15250_, _15249_, _07441_);
  not (_15251_, _08385_);
  and (_15252_, _15251_, _06836_);
  nor (_15253_, _15252_, _08384_);
  and (_15254_, _15253_, _08700_);
  nor (_15255_, _15253_, _08700_);
  or (_15256_, _15255_, _15254_);
  or (_15257_, _15256_, _08128_);
  nor (_15258_, _08051_, _04509_);
  or (_15259_, _15258_, _06835_);
  and (_15260_, _08049_, _05898_);
  and (_15261_, _04063_, _03320_);
  nor (_15262_, _04063_, _03320_);
  or (_15263_, _15262_, _15261_);
  and (_15264_, _15263_, _08048_);
  or (_15265_, _15264_, _08051_);
  or (_15266_, _15265_, _15260_);
  and (_15267_, _15266_, _03262_);
  or (_15268_, _15267_, _04509_);
  and (_15269_, _15268_, _15259_);
  or (_15270_, _15269_, _03599_);
  nor (_15271_, _05371_, \oc8051_golden_model_1.ACC [1]);
  and (_15272_, _12234_, _05371_);
  nor (_15273_, _15272_, _15271_);
  or (_15274_, _15273_, _04515_);
  and (_15275_, _15274_, _15270_);
  or (_15276_, _15275_, _08063_);
  nor (_15277_, _08070_, \oc8051_golden_model_1.PSW [6]);
  nor (_15278_, _15277_, \oc8051_golden_model_1.ACC [1]);
  and (_15279_, _15277_, \oc8051_golden_model_1.ACC [1]);
  nor (_15280_, _15279_, _15278_);
  nand (_15281_, _15280_, _08063_);
  and (_15282_, _15281_, _03604_);
  and (_15283_, _15282_, _15276_);
  nor (_15284_, _05983_, _03320_);
  and (_15285_, _12238_, _05983_);
  nor (_15286_, _15285_, _15284_);
  nor (_15287_, _15286_, _03516_);
  nor (_15288_, _15249_, _04524_);
  or (_15289_, _15288_, _08042_);
  or (_15290_, _15289_, _15287_);
  or (_15291_, _15290_, _15283_);
  or (_15292_, _08041_, _05898_);
  and (_15293_, _15292_, _15291_);
  or (_15294_, _15293_, _04529_);
  or (_15295_, _06835_, _08102_);
  and (_15296_, _15295_, _03611_);
  and (_15297_, _15296_, _15294_);
  nor (_15298_, _08223_, _03611_);
  or (_15299_, _15298_, _08106_);
  or (_15300_, _15299_, _15297_);
  nand (_15301_, _08106_, _07530_);
  and (_15302_, _15301_, _15300_);
  or (_15303_, _15302_, _03511_);
  and (_15304_, _12224_, _05983_);
  nor (_15305_, _15304_, _15284_);
  nand (_15306_, _15305_, _03511_);
  and (_15307_, _15306_, _03505_);
  and (_15308_, _15307_, _15303_);
  and (_15309_, _15285_, _12253_);
  nor (_15310_, _15309_, _15284_);
  nor (_15311_, _15310_, _03505_);
  or (_15312_, _15311_, _06919_);
  or (_15313_, _15312_, _15308_);
  and (_15314_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_15315_, _15314_, _07765_);
  nor (_15316_, _15315_, _07380_);
  or (_15317_, _15316_, _06925_);
  and (_15318_, _15317_, _08037_);
  and (_15319_, _15318_, _15313_);
  and (_15320_, _15251_, _04491_);
  nor (_15321_, _15320_, _08384_);
  and (_15322_, _15321_, _08659_);
  nor (_15323_, _15321_, _08659_);
  or (_15324_, _15323_, _15322_);
  and (_15325_, _15324_, _08038_);
  or (_15326_, _15325_, _08032_);
  or (_15327_, _15326_, _15319_);
  and (_15328_, _15327_, _15257_);
  or (_15329_, _15328_, _03635_);
  nor (_15330_, _08238_, _08385_);
  nor (_15331_, _15330_, _08384_);
  and (_15332_, _15331_, _08746_);
  nor (_15333_, _15331_, _08746_);
  or (_15334_, _15333_, _15332_);
  nand (_15335_, _15334_, _03635_);
  and (_15336_, _15335_, _08161_);
  and (_15337_, _15336_, _15329_);
  nor (_15338_, _08390_, _08161_);
  or (_15339_, _15338_, _03371_);
  or (_15340_, _15339_, _15337_);
  nand (_15341_, _04434_, _03371_);
  and (_15342_, _15341_, _03501_);
  and (_15343_, _15342_, _15340_);
  nor (_15344_, _12270_, _08421_);
  nor (_15345_, _15344_, _15284_);
  nor (_15346_, _15345_, _03501_);
  or (_15347_, _15346_, _07441_);
  or (_15348_, _15347_, _15343_);
  and (_15349_, _15348_, _15250_);
  or (_15350_, _15349_, _05969_);
  and (_15351_, _06835_, _05371_);
  nor (_15352_, _15351_, _15240_);
  nand (_15353_, _15352_, _05969_);
  and (_15354_, _15353_, _03275_);
  and (_15355_, _15354_, _15350_);
  nor (_15356_, _12330_, _07957_);
  nor (_15357_, _15356_, _15240_);
  nor (_15358_, _15357_, _03275_);
  or (_15359_, _15358_, _07455_);
  or (_15360_, _15359_, _15355_);
  nand (_15361_, _07713_, _07455_);
  and (_15362_, _15361_, _15360_);
  or (_15363_, _15362_, _03313_);
  and (_15364_, _15363_, _15247_);
  or (_15365_, _15364_, _03650_);
  and (_15366_, _05371_, _04347_);
  nor (_15367_, _15366_, _15271_);
  or (_15368_, _15367_, _04582_);
  and (_15369_, _15368_, _08446_);
  and (_15370_, _15369_, _15365_);
  nor (_15371_, _08446_, _04434_);
  or (_15372_, _15371_, _08451_);
  or (_15373_, _15372_, _15370_);
  or (_15374_, _08452_, _08659_);
  nor (_15375_, _11837_, _08462_);
  and (_15376_, _15375_, _15374_);
  and (_15377_, _15376_, _15373_);
  and (_15378_, _11839_, _03170_);
  not (_15379_, _08659_);
  nor (_15380_, _15375_, _15379_);
  or (_15381_, _15380_, _15378_);
  or (_15382_, _15381_, _15377_);
  nand (_15383_, _15378_, _15379_);
  and (_15384_, _15383_, _07953_);
  and (_15385_, _15384_, _15382_);
  and (_15386_, _08700_, _07952_);
  or (_15387_, _15386_, _03776_);
  or (_15388_, _15387_, _15385_);
  or (_15389_, _12347_, _03777_);
  and (_15390_, _15389_, _08473_);
  and (_15391_, _15390_, _15388_);
  and (_15392_, _08472_, _08383_);
  or (_15393_, _15392_, _03649_);
  or (_15394_, _15393_, _15391_);
  and (_15395_, _15394_, _15246_);
  or (_15396_, _15395_, _03778_);
  nor (_15397_, _06886_, _04194_);
  not (_15398_, _15397_);
  or (_15399_, _15240_, _04589_);
  and (_15400_, _15399_, _15398_);
  and (_15401_, _15400_, _15396_);
  and (_15402_, _03568_, _03237_);
  or (_15403_, _15402_, _04200_);
  and (_15404_, _15397_, _08657_);
  or (_15405_, _15404_, _15403_);
  or (_15406_, _15405_, _15401_);
  not (_15407_, _15403_);
  or (_15408_, _15407_, _08657_);
  and (_15409_, _15408_, _15406_);
  or (_15410_, _15409_, _04198_);
  or (_15411_, _08698_, _07944_);
  and (_15412_, _15411_, _03772_);
  and (_15413_, _15412_, _15410_);
  or (_15414_, _12345_, _07942_);
  and (_15415_, _15414_, _11368_);
  or (_15416_, _15415_, _15413_);
  or (_15417_, _08381_, _08500_);
  and (_15418_, _15417_, _04596_);
  and (_15419_, _15418_, _15416_);
  or (_15420_, _15419_, _15243_);
  and (_15421_, _15420_, _15009_);
  nor (_15422_, _08658_, _15009_);
  or (_15423_, _15422_, _15421_);
  and (_15424_, _15423_, _15170_);
  nor (_15425_, _15170_, _08658_);
  or (_15426_, _15425_, _04207_);
  or (_15427_, _15426_, _15424_);
  nand (_15428_, _08699_, _04207_);
  and (_15429_, _15428_, _03785_);
  and (_15430_, _15429_, _15427_);
  nand (_15431_, _12346_, _08525_);
  and (_15432_, _15431_, _11358_);
  or (_15433_, _15432_, _15430_);
  and (_15434_, _15433_, _15239_);
  or (_15435_, _15434_, _03653_);
  nor (_15436_, _12218_, _07957_);
  or (_15437_, _15436_, _15240_);
  or (_15438_, _15437_, _04608_);
  and (_15439_, _15438_, _07933_);
  and (_15440_, _15439_, _15435_);
  and (_15441_, _07915_, _07910_);
  nor (_15442_, _15441_, _07916_);
  or (_15443_, _15442_, _08539_);
  and (_15444_, _15443_, _11898_);
  or (_15445_, _15444_, _15440_);
  and (_15446_, _08550_, _08019_);
  nor (_15447_, _15446_, _08551_);
  or (_15448_, _15447_, _08541_);
  and (_15449_, _15448_, _15445_);
  or (_15450_, _15449_, _03782_);
  and (_15451_, _08581_, _08579_);
  nor (_15452_, _15451_, _08582_);
  or (_15453_, _15452_, _03783_);
  and (_15454_, _15453_, _08602_);
  and (_15455_, _15454_, _15450_);
  and (_15456_, _08612_, _08610_);
  nor (_15457_, _15456_, _08613_);
  and (_15458_, _15457_, _08569_);
  or (_15459_, _15458_, _08600_);
  or (_15460_, _15459_, _15455_);
  and (_15461_, _15460_, _15238_);
  or (_15462_, _15461_, _10362_);
  nor (_15463_, _08660_, _08659_);
  nor (_15464_, _15463_, _08661_);
  or (_15465_, _15464_, _09696_);
  and (_15466_, _15465_, _10369_);
  and (_15467_, _15466_, _15462_);
  nor (_15468_, _08701_, _08700_);
  nor (_15469_, _15468_, _08702_);
  and (_15470_, _15469_, _08679_);
  or (_15471_, _15470_, _08722_);
  or (_15472_, _15471_, _15467_);
  and (_15473_, _08748_, _08746_);
  nor (_15474_, _15473_, _08749_);
  or (_15475_, _15474_, _03525_);
  nor (_15476_, _08787_, _08383_);
  nor (_15477_, _15476_, _08788_);
  or (_15478_, _15477_, _08771_);
  and (_15479_, _15478_, _08770_);
  and (_15480_, _15479_, _15475_);
  and (_15481_, _15480_, _15472_);
  and (_15482_, _08769_, \oc8051_golden_model_1.ACC [0]);
  or (_15483_, _15482_, _03809_);
  or (_15484_, _15483_, _15481_);
  or (_15485_, _15273_, _04260_);
  and (_15486_, _15485_, _08810_);
  and (_15487_, _15486_, _15484_);
  nor (_15488_, _08839_, _08815_);
  and (_15489_, _15488_, _09690_);
  nor (_15490_, _15489_, _11952_);
  or (_15491_, _15490_, _15487_);
  nand (_15492_, _08814_, _07634_);
  and (_15493_, _15492_, _03206_);
  and (_15494_, _15493_, _15491_);
  nor (_15495_, _15305_, _03206_);
  or (_15496_, _15495_, _03816_);
  or (_15497_, _15496_, _15494_);
  nor (_15498_, _15272_, _15240_);
  nand (_15499_, _15498_, _03816_);
  and (_15500_, _15499_, _08832_);
  and (_15501_, _15500_, _15497_);
  nor (_15502_, _15488_, _08838_);
  nor (_15503_, _15502_, _11974_);
  or (_15504_, _15503_, _15501_);
  nand (_15505_, _08838_, _07634_);
  and (_15506_, _15505_, _43227_);
  and (_15507_, _15506_, _15504_);
  or (_15508_, _15507_, _15237_);
  and (_43434_, _15508_, _41991_);
  nor (_15509_, _43227_, _07634_);
  nand (_15510_, _08769_, _03320_);
  nand (_15511_, _08600_, _03320_);
  nand (_15512_, _08524_, _08784_);
  nand (_15513_, _08654_, _03954_);
  and (_15514_, _15149_, _08653_);
  nor (_15515_, _05371_, _07634_);
  and (_15516_, _12538_, _05371_);
  nor (_15517_, _15516_, _15515_);
  nand (_15518_, _15517_, _03649_);
  and (_15519_, _15375_, _08452_);
  or (_15520_, _15519_, _08655_);
  nand (_15521_, _03898_, _03313_);
  nor (_15522_, _07957_, _05130_);
  nor (_15523_, _15522_, _15515_);
  nand (_15524_, _15523_, _07441_);
  nand (_15525_, _08042_, _05130_);
  or (_15526_, _15258_, _06839_);
  nand (_15527_, _08049_, _05130_);
  nor (_15528_, _04063_, _07634_);
  and (_15529_, _04063_, _07634_);
  nor (_15530_, _15529_, _15528_);
  nand (_15531_, _15530_, _08048_);
  and (_15532_, _15531_, _15527_);
  or (_15533_, _15532_, _08051_);
  and (_15534_, _15533_, _03262_);
  or (_15535_, _15534_, _04509_);
  and (_15536_, _15535_, _15526_);
  and (_15537_, _15536_, _04515_);
  nor (_15538_, _12430_, _07957_);
  nor (_15539_, _15538_, _15515_);
  nor (_15540_, _15539_, _04515_);
  or (_15541_, _15540_, _08063_);
  or (_15542_, _15541_, _15537_);
  nand (_15543_, _15277_, \oc8051_golden_model_1.ACC [2]);
  and (_15544_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_15545_, _15544_, _08069_);
  or (_15546_, _15545_, _15277_);
  and (_15547_, _15546_, _15543_);
  nand (_15548_, _15547_, _08063_);
  and (_15549_, _15548_, _03604_);
  and (_15550_, _15549_, _15542_);
  nor (_15551_, _05983_, _07634_);
  and (_15552_, _12416_, _05983_);
  nor (_15553_, _15552_, _15551_);
  nor (_15554_, _15553_, _03516_);
  nor (_15555_, _15523_, _04524_);
  or (_15556_, _15555_, _08042_);
  or (_15557_, _15556_, _15554_);
  or (_15558_, _15557_, _15550_);
  and (_15559_, _15558_, _15525_);
  or (_15560_, _15559_, _04529_);
  or (_15561_, _06839_, _08102_);
  and (_15562_, _15561_, _03611_);
  and (_15563_, _15562_, _15560_);
  nor (_15564_, _08208_, _03611_);
  or (_15565_, _15564_, _08106_);
  or (_15566_, _15565_, _15563_);
  nand (_15567_, _08106_, _07484_);
  and (_15568_, _15567_, _15566_);
  or (_15569_, _15568_, _03511_);
  and (_15570_, _12414_, _05983_);
  nor (_15571_, _15570_, _15551_);
  nand (_15572_, _15571_, _03511_);
  and (_15573_, _15572_, _03505_);
  and (_15574_, _15573_, _15569_);
  and (_15575_, _15552_, _12447_);
  nor (_15576_, _15575_, _15551_);
  nor (_15577_, _15576_, _03505_);
  or (_15578_, _15577_, _06919_);
  or (_15579_, _15578_, _15574_);
  nor (_15580_, _07382_, _07380_);
  nor (_15581_, _15580_, _07383_);
  or (_15582_, _15581_, _06925_);
  and (_15583_, _15582_, _15579_);
  or (_15584_, _15583_, _08038_);
  and (_15585_, _04699_, \oc8051_golden_model_1.ACC [1]);
  and (_15586_, _04491_, _03397_);
  nor (_15587_, _15586_, _08659_);
  nor (_15588_, _15587_, _15585_);
  nor (_15589_, _08655_, _15588_);
  and (_15590_, _08655_, _15588_);
  nor (_15591_, _15590_, _15589_);
  nor (_15592_, _15123_, _08659_);
  not (_15593_, _15592_);
  or (_15594_, _15593_, _15591_);
  and (_15595_, _15594_, \oc8051_golden_model_1.PSW [7]);
  nor (_15596_, _15591_, \oc8051_golden_model_1.PSW [7]);
  or (_15597_, _15596_, _15595_);
  nand (_15598_, _15593_, _15591_);
  and (_15599_, _15598_, _15597_);
  nor (_15600_, _15599_, _08032_);
  or (_15601_, _15600_, _11381_);
  and (_15602_, _15601_, _15584_);
  and (_15603_, _06577_, \oc8051_golden_model_1.ACC [1]);
  and (_15604_, _06836_, _03397_);
  nor (_15605_, _15604_, _08700_);
  nor (_15606_, _15605_, _15603_);
  nor (_15607_, _08696_, _15606_);
  and (_15608_, _08696_, _15606_);
  nor (_15609_, _15608_, _15607_);
  nor (_15610_, _15006_, _08700_);
  not (_15611_, _15610_);
  or (_15612_, _15611_, _15609_);
  and (_15614_, _15612_, \oc8051_golden_model_1.PSW [7]);
  nor (_15615_, _15609_, \oc8051_golden_model_1.PSW [7]);
  or (_15616_, _15615_, _15614_);
  nand (_15617_, _15611_, _15609_);
  and (_15618_, _15617_, _15616_);
  nor (_15619_, _15618_, _08128_);
  or (_15620_, _15619_, _03635_);
  or (_15621_, _15620_, _15602_);
  nor (_15622_, _09942_, _08744_);
  or (_15623_, _15622_, _08745_);
  and (_15625_, _08742_, _15623_);
  nor (_15626_, _08742_, _15623_);
  nor (_15627_, _15626_, _15625_);
  and (_15628_, _09944_, \oc8051_golden_model_1.PSW [7]);
  not (_15629_, _15628_);
  nor (_15630_, _15629_, _15627_);
  and (_15631_, _15629_, _15627_);
  nor (_15632_, _15631_, _15630_);
  nand (_15633_, _15632_, _03635_);
  and (_15634_, _15633_, _08161_);
  and (_15636_, _15634_, _15621_);
  nor (_15637_, _04042_, \oc8051_golden_model_1.ACC [0]);
  nor (_15638_, _15637_, _08383_);
  nor (_15639_, _15638_, _10100_);
  nor (_15640_, _08785_, _15639_);
  and (_15641_, _08785_, _15639_);
  nor (_15642_, _15641_, _15640_);
  not (_15643_, _10131_);
  or (_15644_, _15643_, _15642_);
  and (_15645_, _15644_, \oc8051_golden_model_1.PSW [7]);
  nor (_15647_, _15642_, \oc8051_golden_model_1.PSW [7]);
  or (_15648_, _15647_, _15645_);
  nand (_15649_, _15643_, _15642_);
  and (_15650_, _15649_, _15648_);
  nor (_15651_, _15650_, _08161_);
  or (_15652_, _15651_, _03371_);
  or (_15653_, _15652_, _15636_);
  nand (_15654_, _03898_, _03371_);
  and (_15655_, _15654_, _03501_);
  and (_15656_, _15655_, _15653_);
  nor (_15658_, _12465_, _08421_);
  nor (_15659_, _15658_, _15551_);
  nor (_15660_, _15659_, _03501_);
  or (_15661_, _15660_, _07441_);
  or (_15662_, _15661_, _15656_);
  and (_15663_, _15662_, _15524_);
  or (_15664_, _15663_, _05969_);
  and (_15665_, _06839_, _05371_);
  nor (_15666_, _15665_, _15515_);
  nand (_15667_, _15666_, _05969_);
  and (_15669_, _15667_, _03275_);
  and (_15670_, _15669_, _15664_);
  nor (_15671_, _12524_, _07957_);
  nor (_15672_, _15671_, _15515_);
  nor (_15673_, _15672_, _03275_);
  or (_15674_, _15673_, _07455_);
  or (_15675_, _15674_, _15670_);
  or (_15676_, _07648_, _07805_);
  and (_15677_, _15676_, _15675_);
  or (_15678_, _15677_, _03313_);
  and (_15680_, _15678_, _15521_);
  or (_15681_, _15680_, _03650_);
  and (_15682_, _05371_, _06414_);
  nor (_15683_, _15682_, _15515_);
  nand (_15684_, _15683_, _03650_);
  and (_15685_, _15684_, _08446_);
  and (_15686_, _15685_, _15681_);
  or (_15687_, _08446_, _03898_);
  nand (_15688_, _15687_, _15519_);
  or (_15689_, _15688_, _15686_);
  and (_15691_, _15689_, _15520_);
  or (_15692_, _15691_, _15378_);
  nand (_15693_, _15378_, _08656_);
  and (_15694_, _15693_, _07953_);
  and (_15695_, _15694_, _15692_);
  and (_15696_, _08696_, _07952_);
  or (_15697_, _15696_, _03776_);
  or (_15698_, _15697_, _15695_);
  or (_15699_, _12544_, _03777_);
  and (_15700_, _15699_, _08473_);
  and (_15702_, _15700_, _15698_);
  and (_15703_, _08472_, _08785_);
  or (_15704_, _15703_, _03649_);
  or (_15705_, _15704_, _15702_);
  and (_15706_, _15705_, _15518_);
  or (_15707_, _15706_, _03778_);
  or (_15708_, _15515_, _04589_);
  and (_15709_, _15708_, _15150_);
  and (_15710_, _15709_, _15707_);
  nor (_15711_, _15710_, _15514_);
  nor (_15713_, _15711_, _04198_);
  and (_15714_, _08694_, _04198_);
  or (_15715_, _15714_, _03771_);
  or (_15716_, _15715_, _15713_);
  or (_15717_, _12542_, _03772_);
  and (_15718_, _15717_, _08500_);
  and (_15719_, _15718_, _15716_);
  and (_15720_, _08783_, _07942_);
  or (_15721_, _15720_, _15719_);
  and (_15722_, _15721_, _04596_);
  or (_15724_, _15683_, _12543_);
  nor (_15725_, _15724_, _04596_);
  or (_15726_, _15725_, _03954_);
  or (_15727_, _15726_, _15722_);
  and (_15728_, _15727_, _15513_);
  and (_15729_, _15169_, _04562_);
  or (_15730_, _15729_, _15728_);
  nand (_15731_, _15729_, _08654_);
  and (_15732_, _15731_, _08518_);
  and (_15733_, _15732_, _15730_);
  nor (_15735_, _08654_, _08518_);
  or (_15736_, _15735_, _04207_);
  or (_15737_, _15736_, _15733_);
  nand (_15738_, _08695_, _04207_);
  and (_15739_, _15738_, _03785_);
  and (_15740_, _15739_, _15737_);
  nand (_15741_, _12543_, _08525_);
  and (_15742_, _15741_, _11358_);
  or (_15743_, _15742_, _15740_);
  and (_15744_, _15743_, _15512_);
  or (_15746_, _15744_, _03653_);
  nor (_15747_, _12537_, _07957_);
  nor (_15748_, _15747_, _15515_);
  nand (_15749_, _15748_, _03653_);
  and (_15750_, _15749_, _07933_);
  and (_15751_, _15750_, _15746_);
  and (_15752_, _07917_, _07903_);
  nor (_15753_, _15752_, _07918_);
  and (_15754_, _15753_, _08532_);
  or (_15755_, _15754_, _15751_);
  and (_15757_, _15755_, _08541_);
  and (_15758_, _08552_, _08002_);
  nor (_15759_, _15758_, _08553_);
  and (_15760_, _15759_, _08539_);
  or (_15761_, _15760_, _03782_);
  or (_15762_, _15761_, _15757_);
  and (_15763_, _08583_, _08306_);
  nor (_15764_, _15763_, _08584_);
  or (_15765_, _15764_, _03783_);
  and (_15766_, _15765_, _08602_);
  and (_15768_, _15766_, _15762_);
  and (_15769_, _08614_, _08372_);
  nor (_15770_, _15769_, _08615_);
  and (_15771_, _15770_, _08569_);
  or (_15772_, _15771_, _08600_);
  or (_15773_, _15772_, _15768_);
  nand (_15774_, _15773_, _15511_);
  and (_15775_, _15774_, _09696_);
  and (_15776_, _08662_, _08656_);
  nor (_15777_, _15776_, _08663_);
  nor (_15779_, _15777_, _09696_);
  or (_15780_, _15779_, _08679_);
  nor (_15781_, _15780_, _15775_);
  and (_15782_, _08703_, _08697_);
  nor (_15783_, _15782_, _08704_);
  nand (_15784_, _15783_, _08679_);
  nand (_15785_, _15784_, _03525_);
  or (_15786_, _15785_, _15781_);
  and (_15787_, _08750_, _08742_);
  nor (_15788_, _15787_, _08751_);
  or (_15789_, _15788_, _03525_);
  and (_15790_, _15789_, _08771_);
  and (_15791_, _15790_, _15786_);
  and (_15792_, _08789_, _08786_);
  nor (_15793_, _15792_, _08790_);
  and (_15794_, _15793_, _08720_);
  or (_15795_, _15794_, _08769_);
  or (_15796_, _15795_, _15791_);
  and (_15797_, _15796_, _15510_);
  or (_15798_, _15797_, _03809_);
  nand (_15800_, _15539_, _03809_);
  and (_15801_, _15800_, _08810_);
  and (_15802_, _15801_, _15798_);
  and (_15803_, _08069_, _03397_);
  nor (_15804_, _08815_, _07634_);
  or (_15805_, _15804_, _15803_);
  nor (_15806_, _15805_, _08814_);
  nor (_15807_, _15806_, _11952_);
  or (_15808_, _15807_, _15802_);
  nand (_15809_, _08814_, _07628_);
  and (_15811_, _15809_, _03206_);
  and (_15812_, _15811_, _15808_);
  nor (_15813_, _15571_, _03206_);
  or (_15814_, _15813_, _03816_);
  or (_15815_, _15814_, _15812_);
  and (_15816_, _12600_, _05371_);
  nor (_15817_, _15816_, _15515_);
  nand (_15818_, _15817_, _03816_);
  and (_15819_, _15818_, _08832_);
  and (_15820_, _15819_, _15815_);
  and (_15822_, _08839_, \oc8051_golden_model_1.ACC [2]);
  nor (_15823_, _08839_, \oc8051_golden_model_1.ACC [2]);
  nor (_15824_, _15823_, _15822_);
  nor (_15825_, _15824_, _08838_);
  nor (_15826_, _15825_, _11974_);
  or (_15827_, _15826_, _15820_);
  nand (_15828_, _08838_, _07628_);
  and (_15829_, _15828_, _43227_);
  and (_15830_, _15829_, _15827_);
  or (_15831_, _15830_, _15509_);
  and (_43435_, _15831_, _41991_);
  nor (_15833_, _43227_, _07628_);
  nor (_15834_, _08649_, _08651_);
  nor (_15835_, _08664_, _15834_);
  and (_15836_, _08664_, _15834_);
  nor (_15837_, _15836_, _15835_);
  nand (_15838_, _15837_, _10362_);
  and (_15839_, _07919_, _07897_);
  nor (_15840_, _15839_, _07920_);
  or (_15841_, _15840_, _07933_);
  nor (_15843_, _05371_, _07628_);
  and (_15844_, _05371_, _06347_);
  nor (_15845_, _15844_, _15843_);
  or (_15846_, _15845_, _12618_);
  nor (_15847_, _15846_, _04596_);
  and (_15848_, _15843_, _03778_);
  nand (_15849_, _03494_, _03313_);
  nor (_15850_, _07957_, _04944_);
  nor (_15851_, _15850_, _15843_);
  nand (_15852_, _15851_, _07441_);
  and (_15854_, _03898_, \oc8051_golden_model_1.ACC [2]);
  nor (_15855_, _15640_, _15854_);
  nor (_15856_, _10097_, _15855_);
  and (_15857_, _10097_, _15855_);
  nor (_15858_, _15857_, _15856_);
  and (_15859_, _15858_, \oc8051_golden_model_1.PSW [7]);
  nor (_15860_, _15858_, \oc8051_golden_model_1.PSW [7]);
  nor (_15861_, _15860_, _15859_);
  and (_15862_, _15861_, _15645_);
  nor (_15863_, _15861_, _15645_);
  or (_15865_, _15863_, _15862_);
  nand (_15866_, _15865_, _08160_);
  nor (_15867_, _05983_, _07628_);
  and (_15868_, _12638_, _05983_);
  and (_15869_, _15868_, _12653_);
  nor (_15870_, _15869_, _15867_);
  nor (_15871_, _15870_, _03505_);
  nand (_15872_, _08042_, _04944_);
  or (_15873_, _15258_, _06838_);
  nand (_15874_, _08049_, _04944_);
  nor (_15876_, _04063_, _07628_);
  and (_15877_, _04063_, _07628_);
  nor (_15878_, _15877_, _15876_);
  nand (_15879_, _15878_, _08048_);
  and (_15880_, _15879_, _15874_);
  or (_15881_, _15880_, _08051_);
  and (_15882_, _15881_, _03262_);
  or (_15883_, _15882_, _04509_);
  and (_15884_, _15883_, _04515_);
  and (_15885_, _15884_, _15873_);
  nor (_15887_, _12625_, _07957_);
  nor (_15888_, _15887_, _15843_);
  nor (_15889_, _15888_, _04515_);
  or (_15890_, _15889_, _08063_);
  or (_15891_, _15890_, _15885_);
  not (_15892_, \oc8051_golden_model_1.PSW [6]);
  nor (_15893_, _08069_, _15892_);
  nor (_15894_, _15893_, \oc8051_golden_model_1.ACC [3]);
  or (_15895_, _15894_, _08070_);
  nand (_15896_, _15895_, _08063_);
  and (_15898_, _15896_, _15891_);
  or (_15899_, _15898_, _03515_);
  nor (_15900_, _15868_, _15867_);
  nand (_15901_, _15900_, _03515_);
  and (_15902_, _15901_, _04524_);
  and (_15903_, _15902_, _15899_);
  nor (_15904_, _15851_, _04524_);
  or (_15905_, _15904_, _08042_);
  or (_15906_, _15905_, _15903_);
  and (_15907_, _15906_, _15872_);
  or (_15909_, _15907_, _04529_);
  or (_15910_, _06838_, _08102_);
  and (_15911_, _15910_, _03611_);
  and (_15912_, _15911_, _15909_);
  nor (_15913_, _08191_, _03611_);
  or (_15914_, _15913_, _08106_);
  or (_15915_, _15914_, _15912_);
  nand (_15916_, _08106_, _06061_);
  and (_15917_, _15916_, _15915_);
  or (_15918_, _15917_, _03511_);
  and (_15920_, _12622_, _05983_);
  nor (_15921_, _15920_, _15867_);
  nand (_15922_, _15921_, _03511_);
  and (_15923_, _15922_, _03505_);
  and (_15924_, _15923_, _15918_);
  or (_15925_, _15924_, _15871_);
  and (_15926_, _15925_, _06925_);
  nor (_15927_, _07385_, _07383_);
  nor (_15928_, _15927_, _07386_);
  nand (_15929_, _15928_, _06919_);
  nand (_15931_, _15929_, _08037_);
  or (_15932_, _15931_, _15926_);
  and (_15933_, _05130_, \oc8051_golden_model_1.ACC [2]);
  nor (_15934_, _15589_, _15933_);
  nor (_15935_, _15834_, _15934_);
  and (_15936_, _15834_, _15934_);
  nor (_15937_, _15936_, _15935_);
  and (_15938_, _15937_, \oc8051_golden_model_1.PSW [7]);
  nor (_15939_, _15937_, \oc8051_golden_model_1.PSW [7]);
  nor (_15940_, _15939_, _15938_);
  and (_15942_, _15940_, _15595_);
  nor (_15943_, _15940_, _15595_);
  or (_15944_, _15943_, _15942_);
  nand (_15945_, _15944_, _08038_);
  and (_15946_, _15945_, _15932_);
  or (_15947_, _15946_, _08032_);
  and (_15948_, _06714_, \oc8051_golden_model_1.ACC [2]);
  nor (_15949_, _15607_, _15948_);
  nor (_15950_, _08692_, _08693_);
  and (_15951_, _15950_, _15949_);
  nor (_15953_, _15950_, _15949_);
  or (_15954_, _15953_, _15951_);
  nor (_15955_, _15954_, _07911_);
  and (_15956_, _15954_, _07911_);
  nor (_15957_, _15956_, _15955_);
  and (_15958_, _15957_, _15614_);
  nor (_15959_, _15957_, _15614_);
  nor (_15960_, _15959_, _15958_);
  or (_15961_, _15960_, _08128_);
  and (_15962_, _15961_, _03640_);
  and (_15964_, _15962_, _15947_);
  and (_15965_, _09945_, \oc8051_golden_model_1.PSW [7]);
  nor (_15966_, _15625_, _08740_);
  nor (_15967_, _09919_, _15966_);
  and (_15968_, _09919_, _15966_);
  or (_15969_, _15968_, _15967_);
  not (_15970_, _15630_);
  and (_15971_, _15970_, _15969_);
  nor (_15972_, _15971_, _15965_);
  nand (_15973_, _15972_, _08161_);
  and (_15975_, _15973_, _11380_);
  or (_15976_, _15975_, _15964_);
  and (_15977_, _15976_, _15866_);
  or (_15978_, _15977_, _03371_);
  nand (_15979_, _03494_, _03371_);
  and (_15980_, _15979_, _03501_);
  and (_15981_, _15980_, _15978_);
  nor (_15982_, _12671_, _08421_);
  nor (_15983_, _15982_, _15867_);
  nor (_15984_, _15983_, _03501_);
  or (_15986_, _15984_, _07441_);
  or (_15987_, _15986_, _15981_);
  and (_15988_, _15987_, _15852_);
  or (_15989_, _15988_, _05969_);
  and (_15990_, _06838_, _05371_);
  nor (_15991_, _15990_, _15843_);
  nand (_15992_, _15991_, _05969_);
  and (_15993_, _15992_, _03275_);
  and (_15994_, _15993_, _15989_);
  nor (_15995_, _12731_, _07957_);
  nor (_15997_, _15995_, _15843_);
  nor (_15998_, _15997_, _03275_);
  or (_15999_, _15998_, _07455_);
  or (_16000_, _15999_, _15994_);
  or (_16001_, _07595_, _07805_);
  and (_16002_, _16001_, _16000_);
  or (_16003_, _16002_, _03313_);
  and (_16004_, _16003_, _15849_);
  or (_16005_, _16004_, _03650_);
  nand (_16006_, _15845_, _03650_);
  and (_16008_, _16006_, _08446_);
  and (_16009_, _16008_, _16005_);
  nor (_16010_, _08446_, _03494_);
  and (_16011_, _11838_, _15132_);
  not (_16012_, _16011_);
  or (_16013_, _16012_, _16010_);
  or (_16014_, _16013_, _16009_);
  or (_16015_, _16011_, _15834_);
  and (_16016_, _16015_, _07953_);
  and (_16017_, _16016_, _16014_);
  and (_16019_, _15950_, _07952_);
  or (_16020_, _16019_, _03776_);
  or (_16021_, _16020_, _16017_);
  or (_16022_, _12619_, _03777_);
  and (_16023_, _16022_, _08473_);
  and (_16024_, _16023_, _16021_);
  and (_16025_, _08472_, _10097_);
  or (_16026_, _16025_, _03649_);
  or (_16027_, _16026_, _16024_);
  and (_16028_, _12746_, _05371_);
  nor (_16030_, _16028_, _15843_);
  nand (_16031_, _16030_, _03649_);
  and (_16032_, _16031_, _04589_);
  and (_16033_, _16032_, _16027_);
  nor (_16034_, _16033_, _15848_);
  nor (_16035_, _16034_, _08486_);
  or (_16036_, _08651_, _04357_);
  and (_16037_, _16036_, _08490_);
  or (_16038_, _16037_, _16035_);
  nand (_16039_, _08652_, _04357_);
  and (_16041_, _16039_, _07945_);
  and (_16042_, _16041_, _16038_);
  and (_16043_, _08651_, _04200_);
  or (_16044_, _16043_, _04198_);
  or (_16045_, _16044_, _16042_);
  or (_16046_, _08692_, _07944_);
  and (_16047_, _16046_, _03772_);
  and (_16048_, _16047_, _16045_);
  or (_16049_, _12617_, _07942_);
  and (_16050_, _16049_, _11368_);
  or (_16052_, _16050_, _16048_);
  or (_16053_, _08781_, _08500_);
  and (_16054_, _16053_, _04596_);
  and (_16055_, _16054_, _16052_);
  or (_16056_, _16055_, _15847_);
  and (_16057_, _16056_, _15009_);
  nor (_16058_, _08649_, _15009_);
  or (_16059_, _16058_, _15729_);
  or (_16060_, _16059_, _16057_);
  nand (_16061_, _15729_, _08649_);
  and (_16063_, _16061_, _08518_);
  and (_16064_, _16063_, _16060_);
  nor (_16065_, _08649_, _08518_);
  or (_16066_, _16065_, _04207_);
  or (_16067_, _16066_, _16064_);
  nand (_16068_, _08693_, _04207_);
  and (_16069_, _16068_, _03785_);
  and (_16070_, _16069_, _16067_);
  nand (_16071_, _12618_, _08525_);
  and (_16072_, _16071_, _11358_);
  or (_16074_, _16072_, _16070_);
  nand (_16075_, _08524_, _08782_);
  and (_16076_, _16075_, _04608_);
  and (_16077_, _16076_, _16074_);
  nor (_16078_, _12745_, _07957_);
  nor (_16079_, _16078_, _15843_);
  nor (_16080_, _16079_, _04608_);
  or (_16081_, _16080_, _08532_);
  or (_16082_, _16081_, _16077_);
  and (_16083_, _16082_, _15841_);
  or (_16085_, _16083_, _08539_);
  and (_16086_, _08554_, _07997_);
  nor (_16087_, _16086_, _08555_);
  or (_16088_, _16087_, _08541_);
  and (_16089_, _16088_, _03783_);
  and (_16090_, _16089_, _16085_);
  and (_16091_, _08585_, _08301_);
  nor (_16092_, _16091_, _08586_);
  or (_16093_, _16092_, _08569_);
  and (_16094_, _16093_, _08571_);
  or (_16096_, _16094_, _16090_);
  and (_16097_, _08616_, _08367_);
  nor (_16098_, _16097_, _08617_);
  or (_16099_, _16098_, _08602_);
  and (_16100_, _16099_, _08601_);
  and (_16101_, _16100_, _16096_);
  and (_16102_, _08600_, \oc8051_golden_model_1.ACC [2]);
  or (_16103_, _16102_, _10362_);
  or (_16104_, _16103_, _16101_);
  and (_16105_, _16104_, _15838_);
  or (_16107_, _16105_, _08679_);
  nor (_16108_, _08705_, _15950_);
  and (_16109_, _08705_, _15950_);
  nor (_16110_, _16109_, _16108_);
  nand (_16111_, _16110_, _08679_);
  and (_16112_, _16111_, _03525_);
  and (_16113_, _16112_, _16107_);
  nor (_16114_, _08752_, _09919_);
  and (_16115_, _08752_, _09919_);
  nor (_16116_, _16115_, _16114_);
  or (_16118_, _16116_, _08720_);
  and (_16119_, _16118_, _08722_);
  or (_16120_, _16119_, _16113_);
  nor (_16121_, _08791_, _10097_);
  and (_16122_, _08791_, _10097_);
  nor (_16123_, _16122_, _16121_);
  nand (_16124_, _16123_, _08720_);
  and (_16125_, _16124_, _08770_);
  and (_16126_, _16125_, _16120_);
  and (_16127_, _08769_, \oc8051_golden_model_1.ACC [2]);
  or (_16129_, _16127_, _03809_);
  or (_16130_, _16129_, _16126_);
  nand (_16131_, _15888_, _03809_);
  and (_16132_, _16131_, _08810_);
  and (_16133_, _16132_, _16130_);
  nor (_16134_, _15803_, _07628_);
  or (_16135_, _16134_, _08816_);
  nor (_16136_, _16135_, _08814_);
  nor (_16137_, _16136_, _11952_);
  or (_16138_, _16137_, _16133_);
  nand (_16140_, _08814_, _07536_);
  and (_16141_, _16140_, _03206_);
  and (_16142_, _16141_, _16138_);
  nor (_16143_, _15921_, _03206_);
  or (_16144_, _16143_, _03816_);
  or (_16145_, _16144_, _16142_);
  and (_16146_, _12806_, _05371_);
  nor (_16147_, _16146_, _15843_);
  nand (_16148_, _16147_, _03816_);
  and (_16149_, _16148_, _08832_);
  and (_16151_, _16149_, _16145_);
  or (_16152_, _15822_, \oc8051_golden_model_1.ACC [3]);
  and (_16153_, _16152_, _08840_);
  and (_16154_, _16153_, _08831_);
  or (_16155_, _16154_, _08838_);
  or (_16156_, _16155_, _16151_);
  nand (_16157_, _08838_, _07536_);
  and (_16158_, _16157_, _43227_);
  and (_16159_, _16158_, _16156_);
  or (_16160_, _16159_, _15833_);
  and (_43436_, _16160_, _41991_);
  nor (_16162_, _43227_, _07536_);
  nand (_16163_, _08769_, _07628_);
  and (_16164_, _08600_, _07628_);
  nand (_16165_, _08524_, _08779_);
  nor (_16166_, _05371_, _07536_);
  and (_16167_, _12951_, _05371_);
  nor (_16168_, _16167_, _16166_);
  nand (_16169_, _16168_, _03649_);
  nand (_16170_, _04308_, _03313_);
  nor (_16172_, _05840_, _07957_);
  nor (_16173_, _16172_, _16166_);
  nand (_16174_, _16173_, _07441_);
  nor (_16175_, _15966_, _09917_);
  or (_16176_, _16175_, _09918_);
  and (_16177_, _08737_, _16176_);
  nor (_16178_, _08737_, _16176_);
  nor (_16179_, _16178_, _16177_);
  not (_16180_, _15965_);
  nor (_16181_, _16180_, _16179_);
  and (_16183_, _16180_, _16179_);
  nor (_16184_, _16183_, _16181_);
  nand (_16185_, _16184_, _03635_);
  and (_16186_, _16185_, _08161_);
  or (_16187_, _15958_, _15955_);
  and (_16188_, _06838_, _07628_);
  or (_16189_, _06838_, _07628_);
  and (_16190_, _16189_, _15949_);
  or (_16191_, _16190_, _16188_);
  nor (_16192_, _08691_, _16191_);
  and (_16194_, _08691_, _16191_);
  nor (_16195_, _16194_, _16192_);
  and (_16196_, _16195_, \oc8051_golden_model_1.PSW [7]);
  nor (_16197_, _16195_, \oc8051_golden_model_1.PSW [7]);
  nor (_16198_, _16197_, _16196_);
  and (_16199_, _16198_, _16187_);
  nor (_16200_, _16198_, _16187_);
  nor (_16201_, _16200_, _16199_);
  and (_16202_, _16201_, _08032_);
  nand (_16203_, _08042_, _05840_);
  or (_16205_, _08052_, _06843_);
  nand (_16206_, _08049_, _05840_);
  nor (_16207_, _04063_, _07536_);
  and (_16208_, _04063_, _07536_);
  nor (_16209_, _16208_, _16207_);
  nand (_16210_, _16209_, _08048_);
  and (_16211_, _16210_, _16206_);
  or (_16212_, _16211_, _08051_);
  and (_16213_, _16212_, _08061_);
  and (_16214_, _16213_, _16205_);
  nor (_16216_, _12820_, _07957_);
  nor (_16217_, _16216_, _16166_);
  nor (_16218_, _16217_, _04515_);
  or (_16219_, _16218_, _08063_);
  or (_16220_, _16219_, _16214_);
  nor (_16221_, _08070_, \oc8051_golden_model_1.ACC [4]);
  or (_16222_, _16221_, _08076_);
  nand (_16223_, _16222_, _08063_);
  and (_16224_, _16223_, _03604_);
  and (_16225_, _16224_, _16220_);
  nor (_16227_, _05983_, _07536_);
  and (_16228_, _12830_, _05983_);
  nor (_16229_, _16228_, _16227_);
  nor (_16230_, _16229_, _03516_);
  nor (_16231_, _16173_, _04524_);
  or (_16232_, _16231_, _08042_);
  or (_16233_, _16232_, _16230_);
  or (_16234_, _16233_, _16225_);
  and (_16235_, _16234_, _16203_);
  or (_16236_, _16235_, _04529_);
  or (_16238_, _06843_, _08102_);
  and (_16239_, _16238_, _03611_);
  and (_16240_, _16239_, _16236_);
  nor (_16241_, _08269_, _03611_);
  or (_16242_, _16241_, _08106_);
  or (_16243_, _16242_, _16240_);
  nand (_16244_, _08106_, _03397_);
  and (_16245_, _16244_, _16243_);
  or (_16246_, _16245_, _03511_);
  and (_16247_, _12853_, _05983_);
  nor (_16249_, _16247_, _16227_);
  nand (_16250_, _16249_, _03511_);
  and (_16251_, _16250_, _03505_);
  and (_16252_, _16251_, _16246_);
  and (_16253_, _16228_, _12860_);
  nor (_16254_, _16253_, _16227_);
  nor (_16255_, _16254_, _03505_);
  or (_16256_, _16255_, _06919_);
  or (_16257_, _16256_, _16252_);
  nor (_16258_, _07388_, _07386_);
  nor (_16260_, _16258_, _07389_);
  or (_16261_, _16260_, _06925_);
  and (_16262_, _16261_, _16257_);
  or (_16263_, _16262_, _08038_);
  or (_16264_, _15942_, _15938_);
  nor (_16265_, _04944_, \oc8051_golden_model_1.ACC [3]);
  nand (_16266_, _04944_, \oc8051_golden_model_1.ACC [3]);
  and (_16267_, _16266_, _15934_);
  or (_16268_, _16267_, _16265_);
  nor (_16269_, _08648_, _16268_);
  and (_16271_, _08648_, _16268_);
  nor (_16272_, _16271_, _16269_);
  and (_16273_, _16272_, \oc8051_golden_model_1.PSW [7]);
  nor (_16274_, _16272_, \oc8051_golden_model_1.PSW [7]);
  nor (_16275_, _16274_, _16273_);
  and (_16276_, _16275_, _16264_);
  nor (_16277_, _16275_, _16264_);
  nor (_16278_, _16277_, _16276_);
  or (_16279_, _16278_, _08037_);
  and (_16280_, _16279_, _08128_);
  and (_16282_, _16280_, _16263_);
  or (_16283_, _16282_, _03635_);
  or (_16284_, _16283_, _16202_);
  and (_16285_, _16284_, _16186_);
  or (_16286_, _15862_, _15859_);
  or (_16287_, _15855_, _10106_);
  and (_16288_, _16287_, _10105_);
  nor (_16289_, _08780_, _16288_);
  and (_16290_, _08780_, _16288_);
  nor (_16291_, _16290_, _16289_);
  and (_16293_, _16291_, \oc8051_golden_model_1.PSW [7]);
  nor (_16294_, _16291_, \oc8051_golden_model_1.PSW [7]);
  nor (_16295_, _16294_, _16293_);
  and (_16296_, _16295_, _16286_);
  nor (_16297_, _16295_, _16286_);
  nor (_16298_, _16297_, _16296_);
  and (_16299_, _16298_, _08160_);
  or (_16300_, _16299_, _03371_);
  or (_16301_, _16300_, _16285_);
  nand (_16302_, _04308_, _03371_);
  and (_16304_, _16302_, _03501_);
  and (_16305_, _16304_, _16301_);
  nor (_16306_, _12828_, _08421_);
  nor (_16307_, _16306_, _16227_);
  nor (_16308_, _16307_, _03501_);
  or (_16309_, _16308_, _07441_);
  or (_16310_, _16309_, _16305_);
  and (_16311_, _16310_, _16174_);
  or (_16312_, _16311_, _05969_);
  and (_16313_, _06843_, _05371_);
  nor (_16315_, _16313_, _16166_);
  nand (_16316_, _16315_, _05969_);
  and (_16317_, _16316_, _03275_);
  and (_16318_, _16317_, _16312_);
  nor (_16319_, _12936_, _07957_);
  nor (_16320_, _16319_, _16166_);
  nor (_16321_, _16320_, _03275_);
  or (_16322_, _16321_, _07455_);
  or (_16323_, _16322_, _16318_);
  or (_16324_, _07545_, _07805_);
  and (_16326_, _16324_, _16323_);
  or (_16327_, _16326_, _03313_);
  and (_16328_, _16327_, _16170_);
  or (_16329_, _16328_, _03650_);
  and (_16330_, _06375_, _05371_);
  nor (_16331_, _16330_, _16166_);
  nand (_16332_, _16331_, _03650_);
  and (_16333_, _16332_, _08446_);
  and (_16334_, _16333_, _16329_);
  nor (_16335_, _08446_, _04308_);
  or (_16337_, _16335_, _08451_);
  or (_16338_, _16337_, _16334_);
  or (_16339_, _08452_, _08648_);
  and (_16340_, _16339_, _15124_);
  and (_16341_, _16340_, _16338_);
  and (_16342_, _11837_, _08648_);
  or (_16343_, _16342_, _11839_);
  or (_16344_, _16343_, _16341_);
  or (_16345_, _15132_, _08648_);
  and (_16346_, _16345_, _07953_);
  and (_16348_, _16346_, _16344_);
  and (_16349_, _08691_, _07952_);
  or (_16350_, _16349_, _03776_);
  or (_16351_, _16350_, _16348_);
  or (_16352_, _12957_, _03777_);
  and (_16353_, _16352_, _08473_);
  and (_16354_, _16353_, _16351_);
  and (_16355_, _08472_, _08780_);
  or (_16356_, _16355_, _03649_);
  or (_16357_, _16356_, _16354_);
  and (_16359_, _16357_, _16169_);
  or (_16360_, _16359_, _03778_);
  or (_16361_, _16166_, _04589_);
  and (_16362_, _16361_, _15398_);
  and (_16363_, _16362_, _16360_);
  and (_16364_, _15397_, _08646_);
  or (_16365_, _16364_, _15403_);
  or (_16366_, _16365_, _16363_);
  or (_16367_, _15407_, _08646_);
  and (_16368_, _16367_, _16366_);
  or (_16370_, _16368_, _04198_);
  or (_16371_, _08689_, _07944_);
  and (_16372_, _16371_, _03772_);
  and (_16373_, _16372_, _16370_);
  or (_16374_, _12955_, _07942_);
  and (_16375_, _16374_, _11368_);
  or (_16376_, _16375_, _16373_);
  or (_16377_, _08778_, _08500_);
  and (_16378_, _16377_, _04596_);
  and (_16379_, _16378_, _16376_);
  or (_16381_, _16331_, _12956_);
  nor (_16382_, _16381_, _04596_);
  nand (_16383_, _03235_, _03134_);
  not (_16384_, _16383_);
  or (_16385_, _16384_, _16382_);
  or (_16386_, _16385_, _16379_);
  nand (_16387_, _16384_, _08647_);
  and (_16388_, _16387_, _16386_);
  or (_16389_, _16388_, _04207_);
  nand (_16390_, _08690_, _04207_);
  and (_16392_, _16390_, _03785_);
  and (_16393_, _16392_, _16389_);
  nand (_16394_, _12956_, _08525_);
  and (_16395_, _16394_, _11358_);
  or (_16396_, _16395_, _16393_);
  and (_16397_, _16396_, _16165_);
  or (_16398_, _16397_, _03653_);
  nor (_16399_, _12949_, _07957_);
  nor (_16400_, _16399_, _16166_);
  nand (_16401_, _16400_, _03653_);
  and (_16403_, _16401_, _07933_);
  and (_16404_, _16403_, _16398_);
  and (_16405_, _07921_, _07887_);
  nor (_16406_, _16405_, _07922_);
  or (_16407_, _16406_, _08539_);
  and (_16408_, _16407_, _11898_);
  or (_16409_, _16408_, _16404_);
  and (_16410_, _08556_, _07988_);
  nor (_16411_, _16410_, _08557_);
  or (_16412_, _16411_, _08541_);
  and (_16414_, _16412_, _16409_);
  or (_16415_, _16414_, _03782_);
  and (_16416_, _08587_, _08295_);
  nor (_16417_, _16416_, _08588_);
  or (_16418_, _16417_, _03783_);
  and (_16419_, _16418_, _08602_);
  nand (_16420_, _16419_, _16415_);
  and (_16421_, _08618_, _08360_);
  nor (_16422_, _16421_, _08619_);
  nand (_16423_, _16422_, _08569_);
  and (_16425_, _16423_, _08601_);
  and (_16426_, _16425_, _16420_);
  or (_16427_, _16426_, _16164_);
  and (_16428_, _16427_, _09696_);
  nor (_16429_, _08666_, _08648_);
  nor (_16430_, _16429_, _08667_);
  nor (_16431_, _16430_, _09696_);
  or (_16432_, _16431_, _08679_);
  nor (_16433_, _16432_, _16428_);
  nor (_16434_, _08707_, _08691_);
  nor (_16436_, _16434_, _08708_);
  nand (_16437_, _16436_, _08679_);
  nand (_16438_, _16437_, _03525_);
  or (_16439_, _16438_, _16433_);
  nor (_16440_, _08756_, _08738_);
  nor (_16441_, _16440_, _08757_);
  or (_16442_, _16441_, _03525_);
  and (_16443_, _16442_, _08771_);
  and (_16444_, _16443_, _16439_);
  nor (_16445_, _08793_, _08780_);
  nor (_16447_, _16445_, _08794_);
  and (_16448_, _16447_, _08720_);
  or (_16449_, _16448_, _08769_);
  or (_16450_, _16449_, _16444_);
  and (_16451_, _16450_, _16163_);
  or (_16452_, _16451_, _03809_);
  nand (_16453_, _16217_, _03809_);
  and (_16454_, _16453_, _08810_);
  and (_16455_, _16454_, _16452_);
  and (_16456_, _08816_, _07536_);
  nor (_16458_, _08816_, _07536_);
  nor (_16459_, _16458_, _16456_);
  not (_16460_, _16459_);
  and (_16461_, _16460_, _08809_);
  or (_16462_, _16461_, _08814_);
  or (_16463_, _16462_, _16455_);
  nand (_16464_, _08814_, _07530_);
  and (_16465_, _16464_, _03206_);
  and (_16466_, _16465_, _16463_);
  nor (_16467_, _16249_, _03206_);
  or (_16469_, _16467_, _03816_);
  or (_16470_, _16469_, _16466_);
  and (_16471_, _13013_, _05371_);
  nor (_16472_, _16471_, _16166_);
  nand (_16473_, _16472_, _03816_);
  and (_16474_, _16473_, _08832_);
  and (_16475_, _16474_, _16470_);
  and (_16476_, _08840_, _07536_);
  nor (_16477_, _16476_, _08841_);
  and (_16478_, _16477_, _08831_);
  or (_16480_, _16478_, _08838_);
  or (_16481_, _16480_, _16475_);
  nand (_16482_, _08838_, _07530_);
  and (_16483_, _16482_, _43227_);
  and (_16484_, _16483_, _16481_);
  or (_16485_, _16484_, _16162_);
  and (_43437_, _16485_, _41991_);
  nor (_16486_, _43227_, _07530_);
  and (_16487_, _08600_, \oc8051_golden_model_1.ACC [4]);
  nor (_16488_, _05371_, _07530_);
  nor (_16490_, _13152_, _07957_);
  nor (_16491_, _16490_, _16488_);
  nor (_16492_, _16491_, _04608_);
  nand (_16493_, _16384_, _08645_);
  or (_16494_, _08686_, _07944_);
  and (_16495_, _13154_, _05371_);
  nor (_16496_, _16495_, _16488_);
  nand (_16497_, _16496_, _03649_);
  nor (_16498_, _08644_, _08645_);
  or (_16499_, _11838_, _16498_);
  nand (_16501_, _03853_, _03313_);
  nor (_16502_, _05552_, _07957_);
  nor (_16503_, _16502_, _16488_);
  nand (_16504_, _16503_, _07441_);
  and (_16505_, _06806_, \oc8051_golden_model_1.ACC [4]);
  nor (_16506_, _16192_, _16505_);
  nor (_16507_, _08688_, _16506_);
  and (_16508_, _08688_, _16506_);
  nor (_16509_, _16508_, _16507_);
  nor (_16510_, _16509_, _07911_);
  and (_16512_, _16509_, _07911_);
  nor (_16513_, _16512_, _16510_);
  nor (_16514_, _16199_, _16196_);
  not (_16515_, _16514_);
  and (_16516_, _16515_, _16513_);
  nor (_16517_, _16515_, _16513_);
  nor (_16518_, _16517_, _16516_);
  or (_16519_, _16518_, _08128_);
  nor (_16520_, _07391_, _07389_);
  nor (_16521_, _16520_, _07392_);
  and (_16523_, _16521_, _06919_);
  nor (_16524_, _05983_, _07530_);
  and (_16525_, _13051_, _05983_);
  and (_16526_, _16525_, _13066_);
  nor (_16527_, _16526_, _16524_);
  nor (_16528_, _16527_, _03505_);
  nand (_16529_, _08042_, _05552_);
  or (_16530_, _08052_, _06842_);
  nand (_16531_, _08049_, _05552_);
  nor (_16532_, _04063_, _07530_);
  and (_16534_, _04063_, _07530_);
  nor (_16535_, _16534_, _16532_);
  nand (_16536_, _16535_, _08048_);
  and (_16537_, _16536_, _16531_);
  or (_16538_, _16537_, _08051_);
  and (_16539_, _16538_, _08061_);
  and (_16540_, _16539_, _16530_);
  nor (_16541_, _13035_, _07957_);
  nor (_16542_, _16541_, _16488_);
  nor (_16543_, _16542_, _04515_);
  or (_16546_, _16543_, _08063_);
  or (_16547_, _16546_, _16540_);
  and (_16548_, _09963_, _08078_);
  nor (_16549_, _09963_, _08078_);
  nor (_16550_, _16549_, _16548_);
  nand (_16551_, _16550_, _08063_);
  and (_16552_, _16551_, _03604_);
  and (_16553_, _16552_, _16547_);
  nor (_16554_, _16525_, _16524_);
  nor (_16555_, _16554_, _03516_);
  nor (_16557_, _16503_, _04524_);
  or (_16558_, _16557_, _08042_);
  or (_16559_, _16558_, _16555_);
  or (_16560_, _16559_, _16553_);
  and (_16561_, _16560_, _16529_);
  or (_16562_, _16561_, _04529_);
  or (_16563_, _06842_, _08102_);
  and (_16564_, _16563_, _03611_);
  and (_16565_, _16564_, _16562_);
  nor (_16566_, _08255_, _03611_);
  or (_16568_, _16566_, _08106_);
  or (_16569_, _16568_, _16565_);
  nand (_16570_, _08106_, _03320_);
  and (_16571_, _16570_, _16569_);
  or (_16572_, _16571_, _03511_);
  and (_16573_, _13032_, _05983_);
  nor (_16574_, _16573_, _16524_);
  nand (_16575_, _16574_, _03511_);
  and (_16576_, _16575_, _03505_);
  and (_16577_, _16576_, _16572_);
  or (_16579_, _16577_, _16528_);
  and (_16580_, _16579_, _06925_);
  or (_16581_, _16580_, _16523_);
  and (_16582_, _16581_, _08037_);
  and (_16583_, _05840_, \oc8051_golden_model_1.ACC [4]);
  nor (_16584_, _16269_, _16583_);
  not (_16585_, _16498_);
  and (_16586_, _16585_, _16584_);
  nor (_16587_, _16585_, _16584_);
  nor (_16588_, _16587_, _16586_);
  nor (_16590_, _16588_, _07911_);
  and (_16591_, _16588_, _07911_);
  nor (_16592_, _16591_, _16590_);
  nor (_16593_, _16276_, _16273_);
  not (_16594_, _16593_);
  and (_16595_, _16594_, _16592_);
  nor (_16596_, _16594_, _16592_);
  nor (_16597_, _16596_, _16595_);
  and (_16598_, _16597_, _08038_);
  or (_16599_, _16598_, _08032_);
  or (_16601_, _16599_, _16582_);
  and (_16602_, _16601_, _16519_);
  or (_16603_, _16602_, _03635_);
  nor (_16604_, _16177_, _08735_);
  nor (_16605_, _08733_, _16604_);
  and (_16606_, _08733_, _16604_);
  or (_16607_, _16606_, _16605_);
  not (_16608_, _16181_);
  nor (_16609_, _16608_, _16607_);
  and (_16610_, _16608_, _16607_);
  nor (_16612_, _16610_, _16609_);
  nand (_16613_, _16612_, _03635_);
  and (_16614_, _16613_, _08161_);
  and (_16615_, _16614_, _16603_);
  and (_16616_, _04308_, \oc8051_golden_model_1.ACC [4]);
  nor (_16617_, _16289_, _16616_);
  and (_16618_, _10112_, _16617_);
  nor (_16619_, _10112_, _16617_);
  nor (_16620_, _16619_, _16618_);
  and (_16621_, _16620_, \oc8051_golden_model_1.PSW [7]);
  nor (_16623_, _16620_, \oc8051_golden_model_1.PSW [7]);
  nor (_16624_, _16623_, _16621_);
  nor (_16625_, _16296_, _16293_);
  not (_16626_, _16625_);
  and (_16627_, _16626_, _16624_);
  nor (_16628_, _16626_, _16624_);
  nor (_16629_, _16628_, _16627_);
  and (_16630_, _16629_, _08160_);
  or (_16631_, _16630_, _03371_);
  or (_16632_, _16631_, _16615_);
  nand (_16634_, _03853_, _03371_);
  and (_16635_, _16634_, _03501_);
  and (_16636_, _16635_, _16632_);
  nor (_16637_, _13030_, _08421_);
  nor (_16638_, _16637_, _16524_);
  nor (_16639_, _16638_, _03501_);
  or (_16640_, _16639_, _07441_);
  or (_16641_, _16640_, _16636_);
  and (_16642_, _16641_, _16504_);
  or (_16643_, _16642_, _05969_);
  and (_16645_, _06842_, _05371_);
  nor (_16646_, _16645_, _16488_);
  nand (_16647_, _16646_, _05969_);
  and (_16648_, _16647_, _03275_);
  and (_16649_, _16648_, _16643_);
  nor (_16650_, _13139_, _07957_);
  nor (_16651_, _16650_, _16488_);
  nor (_16652_, _16651_, _03275_);
  or (_16653_, _16652_, _07455_);
  or (_16654_, _16653_, _16649_);
  or (_16656_, _07515_, _07805_);
  and (_16657_, _16656_, _16654_);
  or (_16658_, _16657_, _03313_);
  and (_16659_, _16658_, _16501_);
  or (_16660_, _16659_, _03650_);
  and (_16661_, _06358_, _05371_);
  nor (_16662_, _16661_, _16488_);
  nand (_16663_, _16662_, _03650_);
  and (_16664_, _16663_, _08446_);
  and (_16665_, _16664_, _16660_);
  or (_16667_, _08446_, _03853_);
  nand (_16668_, _16667_, _11838_);
  or (_16669_, _16668_, _16665_);
  and (_16670_, _16669_, _16499_);
  or (_16671_, _16670_, _11839_);
  or (_16672_, _15132_, _16498_);
  and (_16673_, _16672_, _07953_);
  and (_16674_, _16673_, _16671_);
  nor (_16675_, _08688_, _07953_);
  or (_16676_, _16675_, _03776_);
  or (_16678_, _16676_, _16674_);
  or (_16679_, _13160_, _03777_);
  and (_16680_, _16679_, _08473_);
  and (_16681_, _16680_, _16678_);
  nor (_16682_, _08473_, _10111_);
  or (_16683_, _16682_, _03649_);
  or (_16684_, _16683_, _16681_);
  and (_16685_, _16684_, _16497_);
  or (_16686_, _16685_, _03778_);
  or (_16687_, _16488_, _04589_);
  and (_16689_, _16687_, _15150_);
  and (_16690_, _16689_, _16686_);
  and (_16691_, _15149_, _08644_);
  or (_16692_, _16691_, _04198_);
  or (_16693_, _16692_, _16690_);
  and (_16694_, _16693_, _16494_);
  or (_16695_, _16694_, _03771_);
  or (_16696_, _13158_, _03772_);
  and (_16697_, _16696_, _08500_);
  and (_16698_, _16697_, _16695_);
  and (_16700_, _08776_, _07942_);
  or (_16701_, _16700_, _16698_);
  and (_16702_, _16701_, _04596_);
  or (_16703_, _16662_, _13159_);
  nor (_16704_, _16703_, _04596_);
  or (_16705_, _16704_, _16384_);
  or (_16706_, _16705_, _16702_);
  and (_16707_, _16706_, _16493_);
  or (_16708_, _16707_, _04207_);
  nand (_16709_, _08687_, _04207_);
  and (_16711_, _16709_, _03785_);
  and (_16712_, _16711_, _16708_);
  nand (_16713_, _13159_, _08525_);
  and (_16714_, _16713_, _11358_);
  or (_16715_, _16714_, _16712_);
  nand (_16716_, _08524_, _08777_);
  and (_16717_, _16716_, _04608_);
  and (_16718_, _16717_, _16715_);
  or (_16719_, _16718_, _16492_);
  and (_16720_, _16719_, _07933_);
  and (_16722_, _07923_, _07881_);
  nor (_16723_, _16722_, _07924_);
  and (_16724_, _16723_, _08532_);
  or (_16725_, _16724_, _08539_);
  or (_16726_, _16725_, _16720_);
  and (_16727_, _08558_, _07986_);
  nor (_16728_, _16727_, _08559_);
  or (_16729_, _16728_, _08541_);
  and (_16730_, _16729_, _03783_);
  and (_16731_, _16730_, _16726_);
  and (_16733_, _08589_, _08290_);
  nor (_16734_, _16733_, _08590_);
  and (_16735_, _16734_, _03782_);
  or (_16736_, _16735_, _08569_);
  or (_16737_, _16736_, _16731_);
  and (_16738_, _08620_, _08355_);
  nor (_16739_, _16738_, _08621_);
  or (_16740_, _16739_, _08602_);
  and (_16741_, _16740_, _08601_);
  and (_16742_, _16741_, _16737_);
  or (_16744_, _16742_, _16487_);
  and (_16745_, _16744_, _09696_);
  and (_16746_, _08668_, _16585_);
  nor (_16747_, _08668_, _16585_);
  nor (_16748_, _16747_, _16746_);
  and (_16749_, _16748_, _10362_);
  or (_16750_, _16749_, _08679_);
  or (_16751_, _16750_, _16745_);
  and (_16752_, _08709_, _08688_);
  nor (_16753_, _16752_, _08710_);
  or (_16755_, _16753_, _10369_);
  and (_16756_, _16755_, _03525_);
  and (_16757_, _16756_, _16751_);
  and (_16758_, _08758_, _08733_);
  nor (_16759_, _16758_, _08759_);
  or (_16760_, _16759_, _08720_);
  and (_16761_, _16760_, _08722_);
  or (_16762_, _16761_, _16757_);
  nor (_16763_, _08795_, _10111_);
  and (_16764_, _08795_, _10111_);
  nor (_16766_, _16764_, _16763_);
  or (_16767_, _16766_, _08771_);
  and (_16768_, _16767_, _08770_);
  and (_16769_, _16768_, _16762_);
  and (_16770_, _08769_, \oc8051_golden_model_1.ACC [4]);
  or (_16771_, _16770_, _03809_);
  or (_16772_, _16771_, _16769_);
  nand (_16773_, _16542_, _03809_);
  and (_16774_, _16773_, _08810_);
  and (_16775_, _16774_, _16772_);
  nor (_16777_, _16456_, _07530_);
  or (_16778_, _16777_, _08817_);
  and (_16779_, _16778_, _08809_);
  or (_16780_, _16779_, _08814_);
  or (_16781_, _16780_, _16775_);
  nand (_16782_, _08814_, _07484_);
  and (_16783_, _16782_, _03206_);
  and (_16784_, _16783_, _16781_);
  nor (_16785_, _16574_, _03206_);
  or (_16786_, _16785_, _03816_);
  or (_16788_, _16786_, _16784_);
  and (_16789_, _13217_, _05371_);
  nor (_16790_, _16789_, _16488_);
  nand (_16791_, _16790_, _03816_);
  and (_16792_, _16791_, _08832_);
  and (_16793_, _16792_, _16788_);
  nor (_16794_, _08841_, \oc8051_golden_model_1.ACC [5]);
  nor (_16795_, _16794_, _08842_);
  and (_16796_, _16795_, _08831_);
  or (_16797_, _16796_, _08838_);
  or (_16799_, _16797_, _16793_);
  nand (_16800_, _08838_, _07484_);
  and (_16801_, _16800_, _43227_);
  and (_16802_, _16801_, _16799_);
  or (_16803_, _16802_, _16486_);
  and (_43438_, _16803_, _41991_);
  nor (_16804_, _43227_, _07484_);
  nand (_16805_, _08769_, _07530_);
  and (_16806_, _08760_, _08729_);
  nor (_16807_, _16806_, _08761_);
  or (_16809_, _16807_, _03525_);
  and (_16810_, _16809_, _08771_);
  nor (_16811_, _05371_, _07484_);
  nor (_16812_, _13243_, _07957_);
  nor (_16813_, _16812_, _16811_);
  nand (_16814_, _16813_, _03653_);
  nand (_16815_, _08684_, _04207_);
  not (_16816_, _08506_);
  nand (_16817_, _16816_, _08642_);
  nor (_16818_, _05080_, _04194_);
  nor (_16820_, _16818_, _15397_);
  not (_16821_, _16820_);
  and (_16822_, _16821_, _08641_);
  and (_16823_, _16811_, _03778_);
  nand (_16824_, _03556_, _03313_);
  nor (_16825_, _05442_, _07957_);
  nor (_16826_, _16825_, _16811_);
  nand (_16827_, _16826_, _07441_);
  nor (_16828_, _16604_, _08731_);
  or (_16829_, _16828_, _08732_);
  and (_16831_, _16829_, _08729_);
  nor (_16832_, _16829_, _08729_);
  nor (_16833_, _16832_, _16831_);
  not (_16834_, _16609_);
  nor (_16835_, _16834_, _16833_);
  and (_16836_, _16834_, _16833_);
  nor (_16837_, _16836_, _16835_);
  nand (_16838_, _16837_, _03635_);
  and (_16839_, _16838_, _08161_);
  or (_16840_, _06842_, _07530_);
  and (_16842_, _06842_, _07530_);
  or (_16843_, _16506_, _16842_);
  and (_16844_, _16843_, _16840_);
  nor (_16845_, _16844_, _08685_);
  and (_16846_, _16844_, _08685_);
  nor (_16847_, _16846_, _16845_);
  nor (_16848_, _16516_, _16510_);
  and (_16849_, _16848_, \oc8051_golden_model_1.PSW [7]);
  nor (_16850_, _16849_, _16847_);
  and (_16851_, _16849_, _16847_);
  nor (_16853_, _16851_, _16850_);
  and (_16854_, _16853_, _08032_);
  nand (_16855_, _08042_, _05442_);
  nor (_16856_, _13235_, _07957_);
  nor (_16857_, _16856_, _16811_);
  nor (_16858_, _16857_, _04515_);
  or (_16859_, _08052_, _06531_);
  nor (_16860_, _08048_, _05442_);
  and (_16861_, _04063_, _07484_);
  nor (_16862_, _04063_, _07484_);
  or (_16864_, _16862_, _16861_);
  and (_16865_, _16864_, _08048_);
  or (_16866_, _16865_, _08051_);
  or (_16867_, _16866_, _16860_);
  and (_16868_, _16867_, _08061_);
  and (_16869_, _16868_, _16859_);
  or (_16870_, _16869_, _16858_);
  and (_16871_, _16870_, _09952_);
  not (_16872_, _08080_);
  nor (_16873_, _16549_, _16872_);
  and (_16875_, _09962_, _08081_);
  nor (_16876_, _16875_, _16873_);
  nor (_16877_, _16876_, _09952_);
  or (_16878_, _16877_, _03515_);
  or (_16879_, _16878_, _16871_);
  nor (_16880_, _05983_, _07484_);
  and (_16881_, _13266_, _05983_);
  nor (_16882_, _16881_, _16880_);
  nand (_16883_, _16882_, _03515_);
  and (_16884_, _16883_, _04524_);
  and (_16886_, _16884_, _16879_);
  nor (_16887_, _16826_, _04524_);
  or (_16888_, _16887_, _08042_);
  or (_16889_, _16888_, _16886_);
  and (_16890_, _16889_, _16855_);
  or (_16891_, _16890_, _04529_);
  or (_16892_, _06531_, _08102_);
  and (_16893_, _16892_, _03611_);
  and (_16894_, _16893_, _16891_);
  nor (_16895_, _08173_, _03611_);
  or (_16897_, _16895_, _08106_);
  or (_16898_, _16897_, _16894_);
  nand (_16899_, _08106_, _07634_);
  and (_16900_, _16899_, _16898_);
  or (_16901_, _16900_, _03511_);
  and (_16902_, _13251_, _05983_);
  nor (_16903_, _16902_, _16880_);
  nand (_16904_, _16903_, _03511_);
  and (_16905_, _16904_, _03505_);
  and (_16906_, _16905_, _16901_);
  and (_16908_, _16881_, _13281_);
  nor (_16909_, _16908_, _16880_);
  nor (_16910_, _16909_, _03505_);
  or (_16911_, _16910_, _06919_);
  or (_16912_, _16911_, _16906_);
  nor (_16913_, _07394_, _07392_);
  nor (_16914_, _16913_, _07395_);
  or (_16915_, _16914_, _06925_);
  and (_16916_, _16915_, _16912_);
  or (_16917_, _16916_, _08038_);
  nand (_16919_, _05552_, \oc8051_golden_model_1.ACC [5]);
  nor (_16920_, _05552_, \oc8051_golden_model_1.ACC [5]);
  or (_16921_, _16584_, _16920_);
  and (_16922_, _16921_, _16919_);
  nor (_16923_, _16922_, _08643_);
  and (_16924_, _16922_, _08643_);
  nor (_16925_, _16924_, _16923_);
  nor (_16926_, _16595_, _16590_);
  and (_16927_, _16926_, \oc8051_golden_model_1.PSW [7]);
  nor (_16928_, _16927_, _16925_);
  and (_16930_, _16927_, _16925_);
  nor (_16931_, _16930_, _16928_);
  or (_16932_, _16931_, _08037_);
  and (_16933_, _16932_, _08128_);
  and (_16934_, _16933_, _16917_);
  or (_16935_, _16934_, _03635_);
  or (_16936_, _16935_, _16854_);
  and (_16937_, _16936_, _16839_);
  or (_16938_, _16617_, _10118_);
  and (_16939_, _16938_, _10117_);
  nor (_16941_, _16939_, _08775_);
  and (_16942_, _16939_, _08775_);
  nor (_16943_, _16942_, _16941_);
  nor (_16944_, _16627_, _16621_);
  and (_16945_, _16944_, \oc8051_golden_model_1.PSW [7]);
  or (_16946_, _16945_, _16943_);
  nand (_16947_, _16945_, _16943_);
  and (_16948_, _16947_, _16946_);
  and (_16949_, _16948_, _08160_);
  or (_16950_, _16949_, _03371_);
  or (_16952_, _16950_, _16937_);
  nand (_16953_, _03556_, _03371_);
  and (_16954_, _16953_, _03501_);
  and (_16955_, _16954_, _16952_);
  nor (_16956_, _13249_, _08421_);
  nor (_16957_, _16956_, _16880_);
  nor (_16958_, _16957_, _03501_);
  or (_16959_, _16958_, _07441_);
  or (_16960_, _16959_, _16955_);
  and (_16961_, _16960_, _16827_);
  or (_16963_, _16961_, _05969_);
  and (_16964_, _06531_, _05371_);
  nor (_16965_, _16964_, _16811_);
  nand (_16966_, _16965_, _05969_);
  and (_16967_, _16966_, _03275_);
  and (_16968_, _16967_, _16963_);
  nor (_16969_, _13356_, _07957_);
  nor (_16970_, _16969_, _16811_);
  nor (_16971_, _16970_, _03275_);
  or (_16972_, _16971_, _07455_);
  or (_16974_, _16972_, _16968_);
  not (_16975_, _07485_);
  and (_16976_, _07489_, _16975_);
  or (_16977_, _16976_, _07805_);
  and (_16978_, _16977_, _16974_);
  or (_16979_, _16978_, _03313_);
  and (_16980_, _16979_, _16824_);
  or (_16981_, _16980_, _03650_);
  and (_16982_, _13363_, _05371_);
  nor (_16983_, _16982_, _16811_);
  nand (_16985_, _16983_, _03650_);
  and (_16986_, _16985_, _08446_);
  and (_16987_, _16986_, _16981_);
  nor (_16988_, _08446_, _03556_);
  or (_16989_, _16988_, _08451_);
  or (_16990_, _16989_, _16987_);
  or (_16991_, _08452_, _08643_);
  and (_16992_, _16991_, _15124_);
  and (_16993_, _16992_, _16990_);
  and (_16994_, _11837_, _08643_);
  or (_16996_, _16994_, _11839_);
  or (_16997_, _16996_, _16993_);
  or (_16998_, _15132_, _08643_);
  and (_16999_, _16998_, _07953_);
  and (_17000_, _16999_, _16997_);
  and (_17001_, _08685_, _07952_);
  or (_17002_, _17001_, _03776_);
  or (_17003_, _17002_, _17000_);
  or (_17004_, _13374_, _03777_);
  and (_17005_, _17004_, _08473_);
  and (_17007_, _17005_, _17003_);
  nor (_17008_, _08473_, _08774_);
  or (_17009_, _17008_, _03649_);
  or (_17010_, _17009_, _17007_);
  and (_17011_, _13245_, _05371_);
  nor (_17012_, _17011_, _16811_);
  nand (_17013_, _17012_, _03649_);
  and (_17014_, _17013_, _04589_);
  and (_17015_, _17014_, _17010_);
  or (_17016_, _17015_, _16823_);
  and (_17018_, _17016_, _16820_);
  nor (_17019_, _17018_, _16822_);
  or (_17020_, _17019_, _04201_);
  and (_17021_, _08641_, _04201_);
  nor (_17022_, _17021_, _04198_);
  nand (_17023_, _17022_, _17020_);
  or (_17024_, _08683_, _07944_);
  and (_17025_, _17024_, _03772_);
  and (_17026_, _17025_, _17023_);
  or (_17027_, _13372_, _07942_);
  and (_17029_, _17027_, _11368_);
  or (_17030_, _17029_, _17026_);
  or (_17031_, _08772_, _08500_);
  and (_17032_, _17031_, _04596_);
  and (_17033_, _17032_, _17030_);
  or (_17034_, _16983_, _13373_);
  nor (_17035_, _17034_, _04596_);
  or (_17036_, _17035_, _16816_);
  or (_17037_, _17036_, _17033_);
  and (_17038_, _17037_, _16817_);
  or (_17040_, _17038_, _08508_);
  nor (_17041_, _08642_, _08514_);
  or (_17042_, _17041_, _08513_);
  and (_17043_, _17042_, _17040_);
  nor (_17044_, _08642_, _08518_);
  or (_17045_, _17044_, _04207_);
  or (_17046_, _17045_, _17043_);
  and (_17047_, _17046_, _16815_);
  or (_17048_, _17047_, _03784_);
  nand (_17049_, _13373_, _03784_);
  and (_17051_, _17049_, _08525_);
  and (_17052_, _17051_, _17048_);
  nor (_17053_, _08525_, _08773_);
  or (_17054_, _17053_, _03653_);
  or (_17055_, _17054_, _17052_);
  and (_17056_, _17055_, _16814_);
  or (_17057_, _17056_, _08532_);
  and (_17058_, _07925_, _07870_);
  nor (_17059_, _17058_, _07926_);
  and (_17060_, _17059_, _08541_);
  or (_17062_, _17060_, _11355_);
  and (_17063_, _17062_, _17057_);
  and (_17064_, _08560_, _08543_);
  nor (_17065_, _17064_, _08561_);
  and (_17066_, _17065_, _08539_);
  or (_17067_, _17066_, _03782_);
  or (_17068_, _17067_, _17063_);
  and (_17069_, _08591_, _08573_);
  nor (_17070_, _17069_, _08592_);
  or (_17071_, _17070_, _03783_);
  and (_17073_, _17071_, _08602_);
  and (_17074_, _17073_, _17068_);
  and (_17075_, _08622_, _08604_);
  nor (_17076_, _17075_, _08623_);
  and (_17077_, _17076_, _08569_);
  or (_17078_, _17077_, _08600_);
  or (_17079_, _17078_, _17074_);
  nor (_17080_, _03988_, _03950_);
  nand (_17081_, _04354_, _03689_);
  and (_17082_, _17081_, _17080_);
  nand (_17084_, _08600_, _07530_);
  and (_17085_, _17084_, _17082_);
  and (_17086_, _17085_, _17079_);
  nor (_17087_, _04236_, _08638_);
  nor (_17088_, _08670_, _08643_);
  nor (_17089_, _17088_, _08671_);
  not (_17090_, _17089_);
  or (_17091_, _17090_, _17082_);
  nand (_17092_, _17091_, _17087_);
  or (_17093_, _17092_, _17086_);
  or (_17095_, _17089_, _17087_);
  and (_17096_, _17095_, _10369_);
  and (_17097_, _17096_, _17093_);
  nor (_17098_, _08711_, _08685_);
  nor (_17099_, _17098_, _08712_);
  and (_17100_, _17099_, _08679_);
  or (_17101_, _17100_, _03524_);
  or (_17102_, _17101_, _17097_);
  and (_17103_, _17102_, _16810_);
  nor (_17104_, _08797_, _08775_);
  nor (_17106_, _17104_, _08798_);
  and (_17107_, _17106_, _08720_);
  or (_17108_, _17107_, _08769_);
  or (_17109_, _17108_, _17103_);
  and (_17110_, _17109_, _16805_);
  or (_17111_, _17110_, _03809_);
  nand (_17112_, _16857_, _03809_);
  and (_17113_, _17112_, _08810_);
  and (_17114_, _17113_, _17111_);
  nor (_17115_, _08817_, _07484_);
  or (_17117_, _17115_, _08818_);
  nor (_17118_, _17117_, _08814_);
  nor (_17119_, _17118_, _11952_);
  or (_17120_, _17119_, _17114_);
  nand (_17121_, _08814_, _06061_);
  and (_17122_, _17121_, _03206_);
  and (_17123_, _17122_, _17120_);
  nor (_17124_, _16903_, _03206_);
  or (_17125_, _17124_, _03816_);
  or (_17126_, _17125_, _17123_);
  and (_17128_, _13425_, _05371_);
  nor (_17129_, _17128_, _16811_);
  nand (_17130_, _17129_, _03816_);
  and (_17131_, _17130_, _08832_);
  and (_17132_, _17131_, _17126_);
  nor (_17133_, _08842_, \oc8051_golden_model_1.ACC [6]);
  nor (_17134_, _17133_, _08843_);
  nor (_17135_, _17134_, _08838_);
  nor (_17136_, _17135_, _11974_);
  or (_17137_, _17136_, _17132_);
  nand (_17139_, _08838_, _06061_);
  and (_17140_, _17139_, _43227_);
  and (_17141_, _17140_, _17137_);
  or (_17142_, _17141_, _16804_);
  and (_43439_, _17142_, _41991_);
  not (_17143_, \oc8051_golden_model_1.DPL [0]);
  nor (_17144_, _43227_, _17143_);
  nor (_17145_, _05319_, _17143_);
  and (_17146_, _05319_, _04491_);
  or (_17147_, _17146_, _17145_);
  or (_17149_, _17147_, _06889_);
  and (_17150_, _05319_, \oc8051_golden_model_1.ACC [0]);
  or (_17151_, _17150_, _17145_);
  or (_17152_, _17151_, _03611_);
  nor (_17153_, _05744_, _08857_);
  or (_17154_, _17153_, _17145_);
  or (_17155_, _17154_, _04515_);
  and (_17156_, _17151_, _04499_);
  nor (_17157_, _04499_, _17143_);
  or (_17158_, _17157_, _03599_);
  or (_17160_, _17158_, _17156_);
  and (_17161_, _17160_, _04524_);
  and (_17162_, _17161_, _17155_);
  and (_17163_, _17147_, _03597_);
  or (_17164_, _17163_, _03603_);
  or (_17165_, _17164_, _17162_);
  and (_17166_, _17165_, _17152_);
  or (_17167_, _17166_, _08880_);
  nand (_17168_, _08880_, \oc8051_golden_model_1.DPL [0]);
  and (_17169_, _17168_, _08865_);
  and (_17171_, _17169_, _17167_);
  nor (_17172_, _04172_, _08865_);
  or (_17173_, _17172_, _07441_);
  or (_17174_, _17173_, _17171_);
  and (_17175_, _17174_, _17149_);
  or (_17176_, _17175_, _05969_);
  and (_17177_, _06836_, _05319_);
  or (_17178_, _17145_, _05970_);
  or (_17179_, _17178_, _17177_);
  and (_17180_, _17179_, _17176_);
  or (_17182_, _17180_, _03644_);
  nor (_17183_, _12129_, _08857_);
  or (_17184_, _17183_, _17145_);
  or (_17185_, _17184_, _03275_);
  and (_17186_, _17185_, _04582_);
  and (_17187_, _17186_, _17182_);
  and (_17188_, _05319_, _06366_);
  or (_17189_, _17188_, _17145_);
  and (_17190_, _17189_, _03650_);
  or (_17191_, _17190_, _03649_);
  or (_17193_, _17191_, _17187_);
  and (_17194_, _12019_, _05319_);
  or (_17195_, _17194_, _17145_);
  or (_17196_, _17195_, _04591_);
  and (_17197_, _17196_, _17193_);
  or (_17198_, _17197_, _03778_);
  and (_17199_, _12145_, _05319_);
  or (_17200_, _17199_, _17145_);
  or (_17201_, _17200_, _04589_);
  and (_17202_, _17201_, _04596_);
  and (_17204_, _17202_, _17198_);
  nand (_17205_, _17189_, _03655_);
  nor (_17206_, _17205_, _17153_);
  or (_17207_, _17206_, _17204_);
  and (_17208_, _17207_, _04594_);
  or (_17209_, _17145_, _05744_);
  and (_17210_, _17151_, _03773_);
  and (_17211_, _17210_, _17209_);
  or (_17212_, _17211_, _03653_);
  or (_17213_, _17212_, _17208_);
  nor (_17215_, _12017_, _08857_);
  or (_17216_, _17145_, _04608_);
  or (_17217_, _17216_, _17215_);
  and (_17218_, _17217_, _04606_);
  and (_17219_, _17218_, _17213_);
  not (_17220_, _03907_);
  nor (_17221_, _12015_, _08857_);
  or (_17222_, _17221_, _17145_);
  and (_17223_, _17222_, _03786_);
  or (_17224_, _17223_, _17220_);
  or (_17226_, _17224_, _17219_);
  or (_17227_, _17154_, _03907_);
  and (_17228_, _17227_, _43227_);
  and (_17229_, _17228_, _17226_);
  or (_17230_, _17229_, _17144_);
  and (_43440_, _17230_, _41991_);
  not (_17231_, \oc8051_golden_model_1.DPL [1]);
  nor (_17232_, _43227_, _17231_);
  and (_17233_, _06835_, _05319_);
  nor (_17234_, _05319_, _17231_);
  or (_17236_, _17234_, _17233_);
  and (_17237_, _17236_, _05969_);
  nor (_17238_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_17239_, _17238_, _08885_);
  and (_17240_, _17239_, _08880_);
  or (_17241_, _05319_, \oc8051_golden_model_1.DPL [1]);
  and (_17242_, _12234_, _05319_);
  not (_17243_, _17242_);
  and (_17244_, _17243_, _17241_);
  or (_17245_, _17244_, _04515_);
  nand (_17247_, _05319_, _03320_);
  and (_17248_, _17247_, _17241_);
  and (_17249_, _17248_, _04499_);
  nor (_17250_, _04499_, _17231_);
  or (_17251_, _17250_, _03599_);
  or (_17252_, _17251_, _17249_);
  and (_17253_, _17252_, _04524_);
  and (_17254_, _17253_, _17245_);
  and (_17255_, _05319_, _05898_);
  or (_17256_, _17255_, _17234_);
  and (_17257_, _17256_, _03597_);
  or (_17258_, _17257_, _03603_);
  or (_17259_, _17258_, _17254_);
  or (_17260_, _17248_, _03611_);
  and (_17261_, _17260_, _08881_);
  and (_17262_, _17261_, _17259_);
  or (_17263_, _17262_, _17240_);
  and (_17264_, _17263_, _08865_);
  nor (_17265_, _04347_, _08865_);
  or (_17266_, _17265_, _07441_);
  or (_17269_, _17266_, _17264_);
  or (_17270_, _17256_, _06889_);
  and (_17271_, _17270_, _05970_);
  and (_17272_, _17271_, _17269_);
  or (_17273_, _17272_, _17237_);
  and (_17274_, _17273_, _03275_);
  nand (_17275_, _12330_, _05319_);
  and (_17276_, _17241_, _03644_);
  and (_17277_, _17276_, _17275_);
  or (_17278_, _17277_, _17274_);
  and (_17279_, _17278_, _03651_);
  nand (_17280_, _05319_, _04347_);
  and (_17281_, _17241_, _03650_);
  and (_17282_, _17281_, _17280_);
  or (_17283_, _12220_, _08857_);
  and (_17284_, _17241_, _03649_);
  and (_17285_, _17284_, _17283_);
  or (_17286_, _17285_, _17282_);
  or (_17287_, _17286_, _17279_);
  and (_17288_, _17287_, _04589_);
  or (_17291_, _12347_, _08857_);
  and (_17292_, _17241_, _03778_);
  and (_17293_, _17292_, _17291_);
  or (_17294_, _17293_, _17288_);
  and (_17295_, _17294_, _04596_);
  or (_17296_, _12219_, _08857_);
  and (_17297_, _17241_, _03655_);
  and (_17298_, _17297_, _17296_);
  or (_17299_, _17298_, _17295_);
  and (_17300_, _17299_, _04594_);
  or (_17302_, _17234_, _05699_);
  and (_17303_, _17248_, _03773_);
  and (_17304_, _17303_, _17302_);
  or (_17305_, _17304_, _17300_);
  and (_17306_, _17305_, _03787_);
  or (_17307_, _17280_, _05699_);
  and (_17308_, _17241_, _03653_);
  and (_17309_, _17308_, _17307_);
  or (_17310_, _17247_, _05699_);
  and (_17311_, _17241_, _03786_);
  and (_17313_, _17311_, _17310_);
  or (_17314_, _17313_, _03809_);
  or (_17315_, _17314_, _17309_);
  or (_17316_, _17315_, _17306_);
  or (_17317_, _17244_, _04260_);
  and (_17318_, _17317_, _17316_);
  or (_17319_, _17318_, _03816_);
  or (_17320_, _17234_, _03820_);
  or (_17321_, _17320_, _17242_);
  and (_17322_, _17321_, _43227_);
  and (_17324_, _17322_, _17319_);
  or (_17325_, _17324_, _17232_);
  and (_43441_, _17325_, _41991_);
  not (_17326_, \oc8051_golden_model_1.DPL [2]);
  nor (_17327_, _43227_, _17326_);
  nor (_17328_, _05319_, _17326_);
  nor (_17329_, _12543_, _08857_);
  or (_17330_, _17329_, _17328_);
  and (_17331_, _17330_, _03786_);
  and (_17332_, _12544_, _05319_);
  or (_17334_, _17332_, _17328_);
  and (_17335_, _17334_, _03778_);
  nor (_17336_, _08857_, _05130_);
  or (_17337_, _17336_, _17328_);
  or (_17338_, _17337_, _06889_);
  nor (_17339_, _08885_, \oc8051_golden_model_1.DPL [2]);
  nor (_17340_, _17339_, _08886_);
  and (_17341_, _17340_, _08880_);
  nor (_17342_, _12430_, _08857_);
  or (_17343_, _17342_, _17328_);
  or (_17345_, _17343_, _04515_);
  and (_17346_, _05319_, \oc8051_golden_model_1.ACC [2]);
  or (_17347_, _17346_, _17328_);
  and (_17348_, _17347_, _04499_);
  nor (_17349_, _04499_, _17326_);
  or (_17350_, _17349_, _03599_);
  or (_17351_, _17350_, _17348_);
  and (_17352_, _17351_, _04524_);
  and (_17353_, _17352_, _17345_);
  and (_17354_, _17337_, _03597_);
  or (_17356_, _17354_, _03603_);
  or (_17357_, _17356_, _17353_);
  or (_17358_, _17347_, _03611_);
  and (_17359_, _17358_, _08881_);
  and (_17360_, _17359_, _17357_);
  or (_17361_, _17360_, _17341_);
  and (_17362_, _17361_, _08865_);
  nor (_17363_, _03943_, _08865_);
  or (_17364_, _17363_, _07441_);
  or (_17365_, _17364_, _17362_);
  and (_17367_, _17365_, _17338_);
  or (_17368_, _17367_, _05969_);
  and (_17369_, _06839_, _05319_);
  or (_17370_, _17328_, _05970_);
  or (_17371_, _17370_, _17369_);
  and (_17372_, _17371_, _03275_);
  and (_17373_, _17372_, _17368_);
  nor (_17374_, _12524_, _08857_);
  or (_17375_, _17374_, _17328_);
  and (_17376_, _17375_, _03644_);
  or (_17378_, _17376_, _17373_);
  or (_17379_, _17378_, _08861_);
  and (_17380_, _12538_, _05319_);
  or (_17381_, _17328_, _04591_);
  or (_17382_, _17381_, _17380_);
  and (_17383_, _05319_, _06414_);
  or (_17384_, _17383_, _17328_);
  or (_17385_, _17384_, _04582_);
  and (_17386_, _17385_, _04589_);
  and (_17387_, _17386_, _17382_);
  and (_17389_, _17387_, _17379_);
  or (_17390_, _17389_, _17335_);
  and (_17391_, _17390_, _04596_);
  or (_17392_, _17328_, _05793_);
  and (_17393_, _17384_, _03655_);
  and (_17394_, _17393_, _17392_);
  or (_17395_, _17394_, _17391_);
  and (_17396_, _17395_, _04594_);
  and (_17397_, _17347_, _03773_);
  and (_17398_, _17397_, _17392_);
  or (_17400_, _17398_, _03653_);
  or (_17401_, _17400_, _17396_);
  nor (_17402_, _12537_, _08857_);
  or (_17403_, _17328_, _04608_);
  or (_17404_, _17403_, _17402_);
  and (_17405_, _17404_, _04606_);
  and (_17406_, _17405_, _17401_);
  or (_17407_, _17406_, _17331_);
  and (_17408_, _17407_, _04260_);
  and (_17409_, _17343_, _03809_);
  or (_17411_, _17409_, _03816_);
  or (_17412_, _17411_, _17408_);
  and (_17413_, _12600_, _05319_);
  or (_17414_, _17328_, _03820_);
  or (_17415_, _17414_, _17413_);
  and (_17416_, _17415_, _43227_);
  and (_17417_, _17416_, _17412_);
  or (_17418_, _17417_, _17327_);
  and (_43442_, _17418_, _41991_);
  not (_17419_, \oc8051_golden_model_1.DPL [3]);
  nor (_17421_, _43227_, _17419_);
  nor (_17422_, _05319_, _17419_);
  nor (_17423_, _12618_, _08857_);
  or (_17424_, _17423_, _17422_);
  and (_17425_, _17424_, _03786_);
  and (_17426_, _12619_, _05319_);
  or (_17427_, _17426_, _17422_);
  and (_17428_, _17427_, _03778_);
  nor (_17429_, _08886_, \oc8051_golden_model_1.DPL [3]);
  nor (_17430_, _17429_, _08887_);
  and (_17432_, _17430_, _08880_);
  nor (_17433_, _12625_, _08857_);
  or (_17434_, _17433_, _17422_);
  or (_17435_, _17434_, _04515_);
  and (_17436_, _05319_, \oc8051_golden_model_1.ACC [3]);
  or (_17437_, _17436_, _17422_);
  and (_17438_, _17437_, _04499_);
  nor (_17439_, _04499_, _17419_);
  or (_17440_, _17439_, _03599_);
  or (_17441_, _17440_, _17438_);
  and (_17443_, _17441_, _04524_);
  and (_17444_, _17443_, _17435_);
  nor (_17445_, _08857_, _04944_);
  or (_17446_, _17445_, _17422_);
  and (_17447_, _17446_, _03597_);
  or (_17448_, _17447_, _03603_);
  or (_17449_, _17448_, _17444_);
  or (_17450_, _17437_, _03611_);
  and (_17451_, _17450_, _08881_);
  and (_17452_, _17451_, _17449_);
  or (_17454_, _17452_, _17432_);
  and (_17455_, _17454_, _08865_);
  nor (_17456_, _03766_, _08865_);
  or (_17457_, _17456_, _07441_);
  or (_17458_, _17457_, _17455_);
  or (_17459_, _17446_, _06889_);
  and (_17460_, _17459_, _17458_);
  or (_17461_, _17460_, _05969_);
  and (_17462_, _06838_, _05319_);
  or (_17463_, _17422_, _05970_);
  or (_17465_, _17463_, _17462_);
  and (_17466_, _17465_, _03275_);
  and (_17467_, _17466_, _17461_);
  nor (_17468_, _12731_, _08857_);
  or (_17469_, _17468_, _17422_);
  and (_17470_, _17469_, _03644_);
  or (_17471_, _17470_, _08861_);
  or (_17472_, _17471_, _17467_);
  and (_17473_, _12746_, _05319_);
  or (_17474_, _17422_, _04591_);
  or (_17476_, _17474_, _17473_);
  and (_17477_, _05319_, _06347_);
  or (_17478_, _17477_, _17422_);
  or (_17479_, _17478_, _04582_);
  and (_17480_, _17479_, _04589_);
  and (_17481_, _17480_, _17476_);
  and (_17482_, _17481_, _17472_);
  or (_17483_, _17482_, _17428_);
  and (_17484_, _17483_, _04596_);
  or (_17485_, _17422_, _05650_);
  and (_17487_, _17478_, _03655_);
  and (_17488_, _17487_, _17485_);
  or (_17489_, _17488_, _17484_);
  and (_17490_, _17489_, _04594_);
  and (_17491_, _17437_, _03773_);
  and (_17492_, _17491_, _17485_);
  or (_17493_, _17492_, _03653_);
  or (_17494_, _17493_, _17490_);
  nor (_17495_, _12745_, _08857_);
  or (_17496_, _17422_, _04608_);
  or (_17498_, _17496_, _17495_);
  and (_17499_, _17498_, _04606_);
  and (_17500_, _17499_, _17494_);
  or (_17501_, _17500_, _17425_);
  and (_17502_, _17501_, _04260_);
  and (_17503_, _17434_, _03809_);
  or (_17504_, _17503_, _03816_);
  or (_17505_, _17504_, _17502_);
  and (_17506_, _12806_, _05319_);
  or (_17507_, _17422_, _03820_);
  or (_17509_, _17507_, _17506_);
  and (_17510_, _17509_, _43227_);
  and (_17511_, _17510_, _17505_);
  or (_17512_, _17511_, _17421_);
  and (_43443_, _17512_, _41991_);
  not (_17513_, \oc8051_golden_model_1.DPL [4]);
  nor (_17514_, _43227_, _17513_);
  nor (_17515_, _05319_, _17513_);
  nor (_17516_, _12956_, _08857_);
  or (_17517_, _17516_, _17515_);
  and (_17519_, _17517_, _03786_);
  nor (_17520_, _05840_, _08857_);
  or (_17521_, _17520_, _17515_);
  or (_17522_, _17521_, _06889_);
  nor (_17523_, _12820_, _08857_);
  or (_17524_, _17523_, _17515_);
  or (_17525_, _17524_, _04515_);
  and (_17526_, _05319_, \oc8051_golden_model_1.ACC [4]);
  or (_17527_, _17526_, _17515_);
  and (_17528_, _17527_, _04499_);
  nor (_17530_, _04499_, _17513_);
  or (_17531_, _17530_, _03599_);
  or (_17532_, _17531_, _17528_);
  and (_17533_, _17532_, _04524_);
  and (_17534_, _17533_, _17525_);
  and (_17535_, _17521_, _03597_);
  or (_17536_, _17535_, _03603_);
  or (_17537_, _17536_, _17534_);
  or (_17538_, _17527_, _03611_);
  and (_17539_, _17538_, _08881_);
  and (_17541_, _17539_, _17537_);
  nor (_17542_, _08887_, \oc8051_golden_model_1.DPL [4]);
  nor (_17543_, _17542_, _08888_);
  and (_17544_, _17543_, _08880_);
  or (_17545_, _17544_, _17541_);
  and (_17546_, _17545_, _08865_);
  nor (_17547_, _06344_, _08865_);
  or (_17548_, _17547_, _07441_);
  or (_17549_, _17548_, _17546_);
  and (_17550_, _17549_, _17522_);
  or (_17552_, _17550_, _05969_);
  and (_17553_, _06843_, _05319_);
  or (_17554_, _17515_, _05970_);
  or (_17555_, _17554_, _17553_);
  and (_17556_, _17555_, _03275_);
  and (_17557_, _17556_, _17552_);
  nor (_17558_, _12936_, _08857_);
  or (_17559_, _17558_, _17515_);
  and (_17560_, _17559_, _03644_);
  or (_17561_, _17560_, _17557_);
  or (_17563_, _17561_, _08861_);
  and (_17564_, _12951_, _05319_);
  or (_17565_, _17515_, _04591_);
  or (_17566_, _17565_, _17564_);
  and (_17567_, _06375_, _05319_);
  or (_17568_, _17567_, _17515_);
  or (_17569_, _17568_, _04582_);
  and (_17570_, _17569_, _04589_);
  and (_17571_, _17570_, _17566_);
  and (_17572_, _17571_, _17563_);
  and (_17574_, _12957_, _05319_);
  or (_17575_, _17574_, _17515_);
  and (_17576_, _17575_, _03778_);
  or (_17577_, _17576_, _17572_);
  and (_17578_, _17577_, _04596_);
  or (_17579_, _17515_, _05889_);
  and (_17580_, _17568_, _03655_);
  and (_17581_, _17580_, _17579_);
  or (_17582_, _17581_, _17578_);
  and (_17583_, _17582_, _04594_);
  and (_17585_, _17527_, _03773_);
  and (_17586_, _17585_, _17579_);
  or (_17587_, _17586_, _03653_);
  or (_17588_, _17587_, _17583_);
  nor (_17589_, _12949_, _08857_);
  or (_17590_, _17515_, _04608_);
  or (_17591_, _17590_, _17589_);
  and (_17592_, _17591_, _04606_);
  and (_17593_, _17592_, _17588_);
  or (_17594_, _17593_, _17519_);
  and (_17596_, _17594_, _04260_);
  and (_17597_, _17524_, _03809_);
  or (_17598_, _17597_, _03816_);
  or (_17599_, _17598_, _17596_);
  and (_17600_, _13013_, _05319_);
  or (_17601_, _17515_, _03820_);
  or (_17602_, _17601_, _17600_);
  and (_17603_, _17602_, _43227_);
  and (_17604_, _17603_, _17599_);
  or (_17605_, _17604_, _17514_);
  and (_43444_, _17605_, _41991_);
  not (_17607_, \oc8051_golden_model_1.DPL [5]);
  nor (_17608_, _43227_, _17607_);
  nor (_17609_, _05319_, _17607_);
  nor (_17610_, _13159_, _08857_);
  or (_17611_, _17610_, _17609_);
  and (_17612_, _17611_, _03786_);
  nor (_17613_, _05552_, _08857_);
  or (_17614_, _17613_, _17609_);
  or (_17615_, _17614_, _06889_);
  nor (_17617_, _13035_, _08857_);
  or (_17618_, _17617_, _17609_);
  or (_17619_, _17618_, _04515_);
  and (_17620_, _05319_, \oc8051_golden_model_1.ACC [5]);
  or (_17621_, _17620_, _17609_);
  and (_17622_, _17621_, _04499_);
  nor (_17623_, _04499_, _17607_);
  or (_17624_, _17623_, _03599_);
  or (_17625_, _17624_, _17622_);
  and (_17626_, _17625_, _04524_);
  and (_17628_, _17626_, _17619_);
  and (_17629_, _17614_, _03597_);
  or (_17630_, _17629_, _03603_);
  or (_17631_, _17630_, _17628_);
  or (_17632_, _17621_, _03611_);
  and (_17633_, _17632_, _08881_);
  and (_17634_, _17633_, _17631_);
  nor (_17635_, _08888_, \oc8051_golden_model_1.DPL [5]);
  nor (_17636_, _17635_, _08889_);
  and (_17637_, _17636_, _08880_);
  or (_17639_, _17637_, _17634_);
  and (_17640_, _17639_, _08865_);
  nor (_17641_, _06313_, _08865_);
  or (_17642_, _17641_, _07441_);
  or (_17643_, _17642_, _17640_);
  and (_17644_, _17643_, _17615_);
  or (_17645_, _17644_, _05969_);
  and (_17646_, _06842_, _05319_);
  or (_17647_, _17609_, _05970_);
  or (_17648_, _17647_, _17646_);
  and (_17650_, _17648_, _03275_);
  and (_17651_, _17650_, _17645_);
  nor (_17652_, _13139_, _08857_);
  or (_17653_, _17652_, _17609_);
  and (_17654_, _17653_, _03644_);
  or (_17655_, _17654_, _17651_);
  or (_17656_, _17655_, _08861_);
  and (_17657_, _13154_, _05319_);
  or (_17658_, _17609_, _04591_);
  or (_17659_, _17658_, _17657_);
  and (_17661_, _06358_, _05319_);
  or (_17662_, _17661_, _17609_);
  or (_17663_, _17662_, _04582_);
  and (_17664_, _17663_, _04589_);
  and (_17665_, _17664_, _17659_);
  and (_17666_, _17665_, _17656_);
  and (_17667_, _13160_, _05319_);
  or (_17668_, _17667_, _17609_);
  and (_17669_, _17668_, _03778_);
  or (_17670_, _17669_, _17666_);
  and (_17672_, _17670_, _04596_);
  or (_17673_, _17609_, _05601_);
  and (_17674_, _17662_, _03655_);
  and (_17675_, _17674_, _17673_);
  or (_17676_, _17675_, _17672_);
  and (_17677_, _17676_, _04594_);
  and (_17678_, _17621_, _03773_);
  and (_17679_, _17678_, _17673_);
  or (_17680_, _17679_, _03653_);
  or (_17681_, _17680_, _17677_);
  nor (_17683_, _13152_, _08857_);
  or (_17684_, _17609_, _04608_);
  or (_17685_, _17684_, _17683_);
  and (_17686_, _17685_, _04606_);
  and (_17687_, _17686_, _17681_);
  or (_17688_, _17687_, _17612_);
  and (_17689_, _17688_, _04260_);
  and (_17690_, _17618_, _03809_);
  or (_17691_, _17690_, _03816_);
  or (_17692_, _17691_, _17689_);
  and (_17694_, _13217_, _05319_);
  or (_17695_, _17609_, _03820_);
  or (_17696_, _17695_, _17694_);
  and (_17697_, _17696_, _43227_);
  and (_17698_, _17697_, _17692_);
  or (_17699_, _17698_, _17608_);
  and (_43447_, _17699_, _41991_);
  not (_17700_, \oc8051_golden_model_1.DPL [6]);
  nor (_17701_, _43227_, _17700_);
  nor (_17702_, _05319_, _17700_);
  nor (_17704_, _13373_, _08857_);
  or (_17705_, _17704_, _17702_);
  and (_17706_, _17705_, _03786_);
  nor (_17707_, _05442_, _08857_);
  or (_17708_, _17707_, _17702_);
  or (_17709_, _17708_, _06889_);
  nor (_17710_, _13235_, _08857_);
  or (_17711_, _17710_, _17702_);
  or (_17712_, _17711_, _04515_);
  and (_17713_, _05319_, \oc8051_golden_model_1.ACC [6]);
  or (_17715_, _17713_, _17702_);
  and (_17716_, _17715_, _04499_);
  nor (_17717_, _04499_, _17700_);
  or (_17718_, _17717_, _03599_);
  or (_17719_, _17718_, _17716_);
  and (_17720_, _17719_, _04524_);
  and (_17721_, _17720_, _17712_);
  and (_17722_, _17708_, _03597_);
  or (_17723_, _17722_, _03603_);
  or (_17724_, _17723_, _17721_);
  or (_17726_, _17715_, _03611_);
  and (_17727_, _17726_, _08881_);
  and (_17728_, _17727_, _17724_);
  nor (_17729_, _08889_, \oc8051_golden_model_1.DPL [6]);
  nor (_17730_, _17729_, _08890_);
  and (_17731_, _17730_, _08880_);
  or (_17732_, _17731_, _17728_);
  and (_17733_, _17732_, _08865_);
  nor (_17734_, _06281_, _08865_);
  or (_17735_, _17734_, _07441_);
  or (_17737_, _17735_, _17733_);
  and (_17738_, _17737_, _17709_);
  or (_17739_, _17738_, _05969_);
  and (_17740_, _06531_, _05319_);
  or (_17741_, _17702_, _05970_);
  or (_17742_, _17741_, _17740_);
  and (_17743_, _17742_, _03275_);
  and (_17744_, _17743_, _17739_);
  nor (_17745_, _13356_, _08857_);
  or (_17746_, _17745_, _17702_);
  and (_17748_, _17746_, _03644_);
  or (_17749_, _17748_, _17744_);
  or (_17750_, _17749_, _08861_);
  and (_17751_, _13245_, _05319_);
  or (_17752_, _17702_, _04591_);
  or (_17753_, _17752_, _17751_);
  and (_17754_, _13363_, _05319_);
  or (_17755_, _17754_, _17702_);
  or (_17756_, _17755_, _04582_);
  and (_17757_, _17756_, _04589_);
  and (_17759_, _17757_, _17753_);
  and (_17760_, _17759_, _17750_);
  and (_17761_, _13374_, _05319_);
  or (_17762_, _17761_, _17702_);
  and (_17763_, _17762_, _03778_);
  or (_17764_, _17763_, _17760_);
  and (_17765_, _17764_, _04596_);
  or (_17766_, _17702_, _05491_);
  and (_17767_, _17755_, _03655_);
  and (_17768_, _17767_, _17766_);
  or (_17770_, _17768_, _17765_);
  and (_17771_, _17770_, _04594_);
  and (_17772_, _17715_, _03773_);
  and (_17773_, _17772_, _17766_);
  or (_17774_, _17773_, _03653_);
  or (_17775_, _17774_, _17771_);
  nor (_17776_, _13243_, _08857_);
  or (_17777_, _17702_, _04608_);
  or (_17778_, _17777_, _17776_);
  and (_17779_, _17778_, _04606_);
  and (_17781_, _17779_, _17775_);
  or (_17782_, _17781_, _17706_);
  and (_17783_, _17782_, _04260_);
  and (_17784_, _17711_, _03809_);
  or (_17785_, _17784_, _03816_);
  or (_17786_, _17785_, _17783_);
  and (_17787_, _13425_, _05319_);
  or (_17788_, _17702_, _03820_);
  or (_17789_, _17788_, _17787_);
  and (_17790_, _17789_, _43227_);
  and (_17792_, _17790_, _17786_);
  or (_17793_, _17792_, _17701_);
  and (_43448_, _17793_, _41991_);
  not (_17794_, \oc8051_golden_model_1.DPH [0]);
  nor (_17795_, _43227_, _17794_);
  and (_17796_, _08892_, \oc8051_golden_model_1.DPH [0]);
  nor (_17797_, _08892_, \oc8051_golden_model_1.DPH [0]);
  nor (_17798_, _17797_, _17796_);
  and (_17799_, _17798_, _08880_);
  nor (_17800_, _05297_, _17794_);
  nor (_17802_, _05744_, _08958_);
  or (_17803_, _17802_, _17800_);
  or (_17804_, _17803_, _04515_);
  and (_17805_, _05297_, \oc8051_golden_model_1.ACC [0]);
  or (_17806_, _17805_, _17800_);
  and (_17807_, _17806_, _04499_);
  nor (_17808_, _04499_, _17794_);
  or (_17809_, _17808_, _03599_);
  or (_17810_, _17809_, _17807_);
  and (_17811_, _17810_, _04524_);
  and (_17813_, _17811_, _17804_);
  and (_17814_, _05297_, _04491_);
  or (_17815_, _17814_, _17800_);
  and (_17816_, _17815_, _03597_);
  or (_17817_, _17816_, _03603_);
  or (_17818_, _17817_, _17813_);
  or (_17819_, _17806_, _03611_);
  and (_17820_, _17819_, _08881_);
  and (_17821_, _17820_, _17818_);
  or (_17822_, _17821_, _17799_);
  and (_17824_, _17822_, _08865_);
  nor (_17825_, _04042_, _08865_);
  or (_17826_, _17825_, _07441_);
  or (_17827_, _17826_, _17824_);
  or (_17828_, _17815_, _06889_);
  and (_17829_, _17828_, _17827_);
  or (_17830_, _17829_, _05969_);
  and (_17831_, _06836_, _05297_);
  or (_17832_, _17800_, _05970_);
  or (_17833_, _17832_, _17831_);
  and (_17835_, _17833_, _17830_);
  or (_17836_, _17835_, _03644_);
  nor (_17837_, _12129_, _08958_);
  or (_17838_, _17837_, _17800_);
  or (_17839_, _17838_, _03275_);
  and (_17840_, _17839_, _04582_);
  and (_17841_, _17840_, _17836_);
  and (_17842_, _05297_, _06366_);
  or (_17843_, _17842_, _17800_);
  and (_17844_, _17843_, _03650_);
  or (_17846_, _17844_, _03649_);
  or (_17847_, _17846_, _17841_);
  and (_17848_, _12019_, _05297_);
  or (_17849_, _17848_, _17800_);
  or (_17850_, _17849_, _04591_);
  and (_17851_, _17850_, _17847_);
  or (_17852_, _17851_, _03778_);
  and (_17853_, _12145_, _05297_);
  or (_17854_, _17853_, _17800_);
  or (_17855_, _17854_, _04589_);
  and (_17857_, _17855_, _04596_);
  and (_17858_, _17857_, _17852_);
  nand (_17859_, _17843_, _03655_);
  nor (_17860_, _17859_, _17802_);
  or (_17861_, _17860_, _17858_);
  and (_17862_, _17861_, _04594_);
  or (_17863_, _17800_, _05744_);
  and (_17864_, _17806_, _03773_);
  and (_17865_, _17864_, _17863_);
  or (_17866_, _17865_, _03653_);
  or (_17868_, _17866_, _17862_);
  nor (_17869_, _12017_, _08958_);
  or (_17870_, _17800_, _04608_);
  or (_17871_, _17870_, _17869_);
  and (_17872_, _17871_, _04606_);
  and (_17873_, _17872_, _17868_);
  nor (_17874_, _12015_, _08958_);
  or (_17875_, _17874_, _17800_);
  and (_17876_, _17875_, _03786_);
  or (_17877_, _17876_, _17220_);
  or (_17879_, _17877_, _17873_);
  or (_17880_, _17803_, _03907_);
  and (_17881_, _17880_, _43227_);
  and (_17882_, _17881_, _17879_);
  or (_17883_, _17882_, _17795_);
  and (_43449_, _17883_, _41991_);
  not (_17884_, \oc8051_golden_model_1.DPH [1]);
  nor (_17885_, _43227_, _17884_);
  or (_17886_, _06835_, _08958_);
  or (_17887_, _05297_, \oc8051_golden_model_1.DPH [1]);
  and (_17889_, _17887_, _05969_);
  and (_17890_, _17889_, _17886_);
  and (_17891_, _12234_, _05297_);
  not (_17892_, _17891_);
  and (_17893_, _17892_, _17887_);
  or (_17894_, _17893_, _04515_);
  nand (_17895_, _05297_, _03320_);
  and (_17896_, _17895_, _17887_);
  and (_17897_, _17896_, _04499_);
  nor (_17898_, _04499_, _17884_);
  or (_17900_, _17898_, _03599_);
  or (_17901_, _17900_, _17897_);
  and (_17902_, _17901_, _04524_);
  and (_17903_, _17902_, _17894_);
  or (_17904_, _08958_, _05898_);
  and (_17905_, _17904_, _17887_);
  and (_17906_, _17905_, _03597_);
  or (_17907_, _17906_, _03603_);
  or (_17908_, _17907_, _17903_);
  or (_17909_, _17896_, _03611_);
  and (_17911_, _17909_, _08881_);
  and (_17912_, _17911_, _17908_);
  nor (_17913_, _17796_, \oc8051_golden_model_1.DPH [1]);
  nor (_17914_, _17913_, _08985_);
  and (_17915_, _17914_, _08880_);
  or (_17916_, _17915_, _17912_);
  and (_17917_, _17916_, _08865_);
  nor (_17918_, _04434_, _08865_);
  or (_17919_, _17918_, _07441_);
  or (_17920_, _17919_, _17917_);
  or (_17922_, _17905_, _06889_);
  and (_17923_, _17922_, _05970_);
  and (_17924_, _17923_, _17920_);
  or (_17925_, _17924_, _17890_);
  and (_17926_, _17925_, _03275_);
  nand (_17927_, _12330_, _05297_);
  and (_17928_, _17887_, _03644_);
  and (_17929_, _17928_, _17927_);
  or (_17930_, _17929_, _17926_);
  and (_17931_, _17930_, _03651_);
  or (_17933_, _12220_, _08958_);
  and (_17934_, _17933_, _03649_);
  nand (_17935_, _05297_, _04347_);
  and (_17936_, _17935_, _03650_);
  or (_17937_, _17936_, _17934_);
  and (_17938_, _17937_, _17887_);
  or (_17939_, _17938_, _17931_);
  and (_17940_, _17939_, _04589_);
  or (_17941_, _12347_, _08958_);
  and (_17942_, _17887_, _03778_);
  and (_17944_, _17942_, _17941_);
  or (_17945_, _17944_, _17940_);
  and (_17946_, _17945_, _04596_);
  or (_17947_, _12219_, _08958_);
  and (_17948_, _17887_, _03655_);
  and (_17949_, _17948_, _17947_);
  or (_17950_, _17949_, _17946_);
  and (_17951_, _17950_, _04594_);
  nor (_17952_, _05297_, _17884_);
  or (_17953_, _17952_, _05699_);
  and (_17955_, _17896_, _03773_);
  and (_17956_, _17955_, _17953_);
  or (_17957_, _17956_, _17951_);
  and (_17958_, _17957_, _03787_);
  or (_17959_, _17935_, _05699_);
  and (_17960_, _17887_, _03653_);
  and (_17961_, _17960_, _17959_);
  or (_17962_, _17895_, _05699_);
  and (_17963_, _17887_, _03786_);
  and (_17964_, _17963_, _17962_);
  or (_17966_, _17964_, _03809_);
  or (_17967_, _17966_, _17961_);
  or (_17968_, _17967_, _17958_);
  or (_17969_, _17893_, _04260_);
  and (_17970_, _17969_, _17968_);
  or (_17971_, _17970_, _03816_);
  or (_17972_, _17952_, _03820_);
  or (_17973_, _17972_, _17891_);
  and (_17974_, _17973_, _43227_);
  and (_17975_, _17974_, _17971_);
  or (_17977_, _17975_, _17885_);
  and (_43452_, _17977_, _41991_);
  not (_17978_, \oc8051_golden_model_1.DPH [2]);
  nor (_17979_, _43227_, _17978_);
  nor (_17980_, _05297_, _17978_);
  nor (_17981_, _12543_, _08958_);
  or (_17982_, _17981_, _17980_);
  and (_17983_, _17982_, _03786_);
  and (_17984_, _12544_, _05297_);
  or (_17985_, _17984_, _17980_);
  and (_17987_, _17985_, _03778_);
  nor (_17988_, _08958_, _05130_);
  or (_17989_, _17988_, _17980_);
  or (_17990_, _17989_, _06889_);
  nor (_17991_, _12430_, _08958_);
  or (_17992_, _17991_, _17980_);
  or (_17993_, _17992_, _04515_);
  and (_17994_, _05297_, \oc8051_golden_model_1.ACC [2]);
  or (_17995_, _17994_, _17980_);
  and (_17996_, _17995_, _04499_);
  nor (_17998_, _04499_, _17978_);
  or (_17999_, _17998_, _03599_);
  or (_18000_, _17999_, _17996_);
  and (_18001_, _18000_, _04524_);
  and (_18002_, _18001_, _17993_);
  and (_18003_, _17989_, _03597_);
  or (_18004_, _18003_, _03603_);
  or (_18005_, _18004_, _18002_);
  or (_18006_, _17995_, _03611_);
  and (_18007_, _18006_, _08881_);
  and (_18009_, _18007_, _18005_);
  or (_18010_, _08985_, \oc8051_golden_model_1.DPH [2]);
  nor (_18011_, _08987_, _08881_);
  and (_18012_, _18011_, _18010_);
  or (_18013_, _18012_, _18009_);
  and (_18014_, _18013_, _08865_);
  nor (_18015_, _03898_, _08865_);
  or (_18016_, _18015_, _07441_);
  or (_18017_, _18016_, _18014_);
  and (_18018_, _18017_, _17990_);
  or (_18020_, _18018_, _05969_);
  and (_18021_, _06839_, _05297_);
  or (_18022_, _17980_, _05970_);
  or (_18023_, _18022_, _18021_);
  and (_18024_, _18023_, _03275_);
  and (_18025_, _18024_, _18020_);
  nor (_18026_, _12524_, _08958_);
  or (_18027_, _18026_, _17980_);
  and (_18028_, _18027_, _03644_);
  or (_18029_, _18028_, _18025_);
  or (_18031_, _18029_, _08861_);
  and (_18032_, _12538_, _05297_);
  or (_18033_, _17980_, _04591_);
  or (_18034_, _18033_, _18032_);
  and (_18035_, _05297_, _06414_);
  or (_18036_, _18035_, _17980_);
  or (_18037_, _18036_, _04582_);
  and (_18038_, _18037_, _04589_);
  and (_18039_, _18038_, _18034_);
  and (_18040_, _18039_, _18031_);
  or (_18042_, _18040_, _17987_);
  and (_18043_, _18042_, _04596_);
  or (_18044_, _17980_, _05793_);
  and (_18045_, _18036_, _03655_);
  and (_18046_, _18045_, _18044_);
  or (_18047_, _18046_, _18043_);
  and (_18048_, _18047_, _04594_);
  and (_18049_, _17995_, _03773_);
  and (_18050_, _18049_, _18044_);
  or (_18051_, _18050_, _03653_);
  or (_18053_, _18051_, _18048_);
  nor (_18054_, _12537_, _08958_);
  or (_18055_, _17980_, _04608_);
  or (_18056_, _18055_, _18054_);
  and (_18057_, _18056_, _04606_);
  and (_18058_, _18057_, _18053_);
  or (_18059_, _18058_, _17983_);
  and (_18060_, _18059_, _04260_);
  and (_18061_, _17992_, _03809_);
  or (_18062_, _18061_, _03816_);
  or (_18064_, _18062_, _18060_);
  and (_18065_, _12600_, _05297_);
  or (_18066_, _17980_, _03820_);
  or (_18067_, _18066_, _18065_);
  and (_18068_, _18067_, _43227_);
  and (_18069_, _18068_, _18064_);
  or (_18070_, _18069_, _17979_);
  and (_43453_, _18070_, _41991_);
  not (_18071_, \oc8051_golden_model_1.DPH [3]);
  nor (_18072_, _43227_, _18071_);
  nor (_18074_, _05297_, _18071_);
  nor (_18075_, _12618_, _08958_);
  or (_18076_, _18075_, _18074_);
  and (_18077_, _18076_, _03786_);
  and (_18078_, _12619_, _05297_);
  or (_18079_, _18078_, _18074_);
  and (_18080_, _18079_, _03778_);
  nor (_18081_, _12625_, _08958_);
  or (_18082_, _18081_, _18074_);
  or (_18083_, _18082_, _04515_);
  and (_18085_, _05297_, \oc8051_golden_model_1.ACC [3]);
  or (_18086_, _18085_, _18074_);
  and (_18087_, _18086_, _04499_);
  nor (_18088_, _04499_, _18071_);
  or (_18089_, _18088_, _03599_);
  or (_18090_, _18089_, _18087_);
  and (_18091_, _18090_, _04524_);
  and (_18092_, _18091_, _18083_);
  nor (_18093_, _08958_, _04944_);
  or (_18094_, _18093_, _18074_);
  and (_18096_, _18094_, _03597_);
  or (_18097_, _18096_, _03603_);
  or (_18098_, _18097_, _18092_);
  or (_18099_, _18086_, _03611_);
  and (_18100_, _18099_, _08881_);
  and (_18101_, _18100_, _18098_);
  or (_18102_, _08987_, \oc8051_golden_model_1.DPH [3]);
  nor (_18103_, _08988_, _08881_);
  and (_18104_, _18103_, _18102_);
  or (_18105_, _18104_, _18101_);
  and (_18107_, _18105_, _08865_);
  nor (_18108_, _08865_, _03494_);
  or (_18109_, _18108_, _07441_);
  or (_18110_, _18109_, _18107_);
  or (_18111_, _18094_, _06889_);
  and (_18112_, _18111_, _18110_);
  or (_18113_, _18112_, _05969_);
  and (_18114_, _06838_, _05297_);
  or (_18115_, _18074_, _05970_);
  or (_18116_, _18115_, _18114_);
  and (_18118_, _18116_, _03275_);
  and (_18119_, _18118_, _18113_);
  nor (_18120_, _12731_, _08958_);
  or (_18121_, _18120_, _18074_);
  and (_18122_, _18121_, _03644_);
  or (_18123_, _18122_, _08861_);
  or (_18124_, _18123_, _18119_);
  and (_18125_, _12746_, _05297_);
  or (_18126_, _18074_, _04591_);
  or (_18127_, _18126_, _18125_);
  and (_18129_, _05297_, _06347_);
  or (_18130_, _18129_, _18074_);
  or (_18131_, _18130_, _04582_);
  and (_18132_, _18131_, _04589_);
  and (_18133_, _18132_, _18127_);
  and (_18134_, _18133_, _18124_);
  or (_18135_, _18134_, _18080_);
  and (_18136_, _18135_, _04596_);
  or (_18137_, _18074_, _05650_);
  and (_18138_, _18130_, _03655_);
  and (_18140_, _18138_, _18137_);
  or (_18141_, _18140_, _18136_);
  and (_18142_, _18141_, _04594_);
  and (_18143_, _18086_, _03773_);
  and (_18144_, _18143_, _18137_);
  or (_18145_, _18144_, _03653_);
  or (_18146_, _18145_, _18142_);
  nor (_18147_, _12745_, _08958_);
  or (_18148_, _18074_, _04608_);
  or (_18149_, _18148_, _18147_);
  and (_18151_, _18149_, _04606_);
  and (_18152_, _18151_, _18146_);
  or (_18153_, _18152_, _18077_);
  and (_18154_, _18153_, _04260_);
  and (_18155_, _18082_, _03809_);
  or (_18156_, _18155_, _03816_);
  or (_18157_, _18156_, _18154_);
  and (_18158_, _12806_, _05297_);
  or (_18159_, _18074_, _03820_);
  or (_18160_, _18159_, _18158_);
  and (_18162_, _18160_, _43227_);
  and (_18163_, _18162_, _18157_);
  or (_18164_, _18163_, _18072_);
  and (_43454_, _18164_, _41991_);
  not (_18165_, \oc8051_golden_model_1.DPH [4]);
  nor (_18166_, _43227_, _18165_);
  nor (_18167_, _05297_, _18165_);
  nor (_18168_, _12956_, _08958_);
  or (_18169_, _18168_, _18167_);
  and (_18170_, _18169_, _03786_);
  nor (_18172_, _05840_, _08958_);
  or (_18173_, _18172_, _18167_);
  or (_18174_, _18173_, _06889_);
  nor (_18175_, _12820_, _08958_);
  or (_18176_, _18175_, _18167_);
  or (_18177_, _18176_, _04515_);
  and (_18178_, _05297_, \oc8051_golden_model_1.ACC [4]);
  or (_18179_, _18178_, _18167_);
  and (_18180_, _18179_, _04499_);
  nor (_18181_, _04499_, _18165_);
  or (_18183_, _18181_, _03599_);
  or (_18184_, _18183_, _18180_);
  and (_18185_, _18184_, _04524_);
  and (_18186_, _18185_, _18177_);
  and (_18187_, _18173_, _03597_);
  or (_18188_, _18187_, _03603_);
  or (_18189_, _18188_, _18186_);
  or (_18190_, _18179_, _03611_);
  and (_18191_, _18190_, _08881_);
  and (_18192_, _18191_, _18189_);
  or (_18194_, _08988_, \oc8051_golden_model_1.DPH [4]);
  nor (_18195_, _08989_, _08881_);
  and (_18196_, _18195_, _18194_);
  or (_18197_, _18196_, _18192_);
  and (_18198_, _18197_, _08865_);
  nor (_18199_, _04308_, _08865_);
  or (_18200_, _18199_, _07441_);
  or (_18201_, _18200_, _18198_);
  and (_18202_, _18201_, _18174_);
  or (_18203_, _18202_, _05969_);
  and (_18205_, _06843_, _05297_);
  or (_18206_, _18167_, _05970_);
  or (_18207_, _18206_, _18205_);
  and (_18208_, _18207_, _03275_);
  and (_18209_, _18208_, _18203_);
  nor (_18210_, _12936_, _08958_);
  or (_18211_, _18210_, _18167_);
  and (_18212_, _18211_, _03644_);
  or (_18213_, _18212_, _18209_);
  or (_18214_, _18213_, _08861_);
  and (_18216_, _12951_, _05297_);
  or (_18217_, _18167_, _04591_);
  or (_18218_, _18217_, _18216_);
  and (_18219_, _06375_, _05297_);
  or (_18220_, _18219_, _18167_);
  or (_18221_, _18220_, _04582_);
  and (_18222_, _18221_, _04589_);
  and (_18223_, _18222_, _18218_);
  and (_18224_, _18223_, _18214_);
  and (_18225_, _12957_, _05297_);
  or (_18227_, _18225_, _18167_);
  and (_18228_, _18227_, _03778_);
  or (_18229_, _18228_, _18224_);
  and (_18230_, _18229_, _04596_);
  or (_18231_, _18167_, _05889_);
  and (_18232_, _18220_, _03655_);
  and (_18233_, _18232_, _18231_);
  or (_18234_, _18233_, _18230_);
  and (_18235_, _18234_, _04594_);
  and (_18236_, _18179_, _03773_);
  and (_18238_, _18236_, _18231_);
  or (_18239_, _18238_, _03653_);
  or (_18240_, _18239_, _18235_);
  nor (_18241_, _12949_, _08958_);
  or (_18242_, _18167_, _04608_);
  or (_18243_, _18242_, _18241_);
  and (_18244_, _18243_, _04606_);
  and (_18245_, _18244_, _18240_);
  or (_18246_, _18245_, _18170_);
  and (_18247_, _18246_, _04260_);
  and (_18249_, _18176_, _03809_);
  or (_18250_, _18249_, _03816_);
  or (_18251_, _18250_, _18247_);
  and (_18252_, _13013_, _05297_);
  or (_18253_, _18167_, _03820_);
  or (_18254_, _18253_, _18252_);
  and (_18255_, _18254_, _43227_);
  and (_18256_, _18255_, _18251_);
  or (_18257_, _18256_, _18166_);
  and (_43455_, _18257_, _41991_);
  not (_18259_, \oc8051_golden_model_1.DPH [5]);
  nor (_18260_, _43227_, _18259_);
  nor (_18261_, _05297_, _18259_);
  nor (_18262_, _13159_, _08958_);
  or (_18263_, _18262_, _18261_);
  and (_18264_, _18263_, _03786_);
  nor (_18265_, _05552_, _08958_);
  or (_18266_, _18265_, _18261_);
  or (_18267_, _18266_, _06889_);
  nor (_18268_, _13035_, _08958_);
  or (_18270_, _18268_, _18261_);
  or (_18271_, _18270_, _04515_);
  and (_18272_, _05297_, \oc8051_golden_model_1.ACC [5]);
  or (_18273_, _18272_, _18261_);
  and (_18274_, _18273_, _04499_);
  nor (_18275_, _04499_, _18259_);
  or (_18276_, _18275_, _03599_);
  or (_18277_, _18276_, _18274_);
  and (_18278_, _18277_, _04524_);
  and (_18279_, _18278_, _18271_);
  and (_18281_, _18266_, _03597_);
  or (_18282_, _18281_, _03603_);
  or (_18283_, _18282_, _18279_);
  or (_18284_, _18273_, _03611_);
  and (_18285_, _18284_, _08881_);
  and (_18286_, _18285_, _18283_);
  or (_18287_, _08989_, \oc8051_golden_model_1.DPH [5]);
  nor (_18288_, _08990_, _08881_);
  and (_18289_, _18288_, _18287_);
  or (_18290_, _18289_, _18286_);
  and (_18292_, _18290_, _08865_);
  nor (_18293_, _03853_, _08865_);
  or (_18294_, _18293_, _07441_);
  or (_18295_, _18294_, _18292_);
  and (_18296_, _18295_, _18267_);
  or (_18297_, _18296_, _05969_);
  and (_18298_, _06842_, _05297_);
  or (_18299_, _18261_, _05970_);
  or (_18300_, _18299_, _18298_);
  and (_18301_, _18300_, _03275_);
  and (_18303_, _18301_, _18297_);
  nor (_18304_, _13139_, _08958_);
  or (_18305_, _18304_, _18261_);
  and (_18306_, _18305_, _03644_);
  or (_18307_, _18306_, _18303_);
  or (_18308_, _18307_, _08861_);
  and (_18309_, _13154_, _05297_);
  or (_18310_, _18261_, _04591_);
  or (_18311_, _18310_, _18309_);
  and (_18312_, _06358_, _05297_);
  or (_18314_, _18312_, _18261_);
  or (_18315_, _18314_, _04582_);
  and (_18316_, _18315_, _04589_);
  and (_18317_, _18316_, _18311_);
  and (_18318_, _18317_, _18308_);
  and (_18319_, _13160_, _05297_);
  or (_18320_, _18319_, _18261_);
  and (_18321_, _18320_, _03778_);
  or (_18322_, _18321_, _18318_);
  and (_18323_, _18322_, _04596_);
  or (_18325_, _18261_, _05601_);
  and (_18326_, _18314_, _03655_);
  and (_18327_, _18326_, _18325_);
  or (_18328_, _18327_, _18323_);
  and (_18329_, _18328_, _04594_);
  and (_18330_, _18273_, _03773_);
  and (_18331_, _18330_, _18325_);
  or (_18332_, _18331_, _03653_);
  or (_18333_, _18332_, _18329_);
  nor (_18334_, _13152_, _08958_);
  or (_18336_, _18261_, _04608_);
  or (_18337_, _18336_, _18334_);
  and (_18338_, _18337_, _04606_);
  and (_18339_, _18338_, _18333_);
  or (_18340_, _18339_, _18264_);
  and (_18341_, _18340_, _04260_);
  and (_18342_, _18270_, _03809_);
  or (_18343_, _18342_, _03816_);
  or (_18344_, _18343_, _18341_);
  and (_18345_, _13217_, _05297_);
  or (_18347_, _18261_, _03820_);
  or (_18348_, _18347_, _18345_);
  and (_18349_, _18348_, _43227_);
  and (_18350_, _18349_, _18344_);
  or (_18351_, _18350_, _18260_);
  and (_43456_, _18351_, _41991_);
  not (_18352_, \oc8051_golden_model_1.DPH [6]);
  nor (_18353_, _43227_, _18352_);
  nor (_18354_, _05297_, _18352_);
  nor (_18355_, _13373_, _08958_);
  or (_18357_, _18355_, _18354_);
  and (_18358_, _18357_, _03786_);
  nor (_18359_, _05442_, _08958_);
  or (_18360_, _18359_, _18354_);
  or (_18361_, _18360_, _06889_);
  nor (_18362_, _13235_, _08958_);
  or (_18363_, _18362_, _18354_);
  or (_18364_, _18363_, _04515_);
  and (_18365_, _05297_, \oc8051_golden_model_1.ACC [6]);
  or (_18366_, _18365_, _18354_);
  and (_18368_, _18366_, _04499_);
  nor (_18369_, _04499_, _18352_);
  or (_18370_, _18369_, _03599_);
  or (_18371_, _18370_, _18368_);
  and (_18372_, _18371_, _04524_);
  and (_18373_, _18372_, _18364_);
  and (_18374_, _18360_, _03597_);
  or (_18375_, _18374_, _03603_);
  or (_18376_, _18375_, _18373_);
  or (_18377_, _18366_, _03611_);
  and (_18379_, _18377_, _08881_);
  and (_18380_, _18379_, _18376_);
  or (_18381_, _08990_, \oc8051_golden_model_1.DPH [6]);
  and (_18382_, _08991_, _08880_);
  and (_18383_, _18382_, _18381_);
  or (_18384_, _18383_, _18380_);
  and (_18385_, _18384_, _08865_);
  nor (_18386_, _08865_, _03556_);
  or (_18387_, _18386_, _07441_);
  or (_18388_, _18387_, _18385_);
  and (_18390_, _18388_, _18361_);
  or (_18391_, _18390_, _05969_);
  and (_18392_, _06531_, _05297_);
  or (_18393_, _18354_, _05970_);
  or (_18394_, _18393_, _18392_);
  and (_18395_, _18394_, _03275_);
  and (_18396_, _18395_, _18391_);
  nor (_18397_, _13356_, _08958_);
  or (_18398_, _18397_, _18354_);
  and (_18399_, _18398_, _03644_);
  or (_18401_, _18399_, _18396_);
  or (_18402_, _18401_, _08861_);
  and (_18403_, _13245_, _05297_);
  or (_18404_, _18354_, _04591_);
  or (_18405_, _18404_, _18403_);
  and (_18406_, _13363_, _05297_);
  or (_18407_, _18406_, _18354_);
  or (_18408_, _18407_, _04582_);
  and (_18409_, _18408_, _04589_);
  and (_18410_, _18409_, _18405_);
  and (_18412_, _18410_, _18402_);
  and (_18413_, _13374_, _05297_);
  or (_18414_, _18413_, _18354_);
  and (_18415_, _18414_, _03778_);
  or (_18416_, _18415_, _18412_);
  and (_18417_, _18416_, _04596_);
  or (_18418_, _18354_, _05491_);
  and (_18419_, _18407_, _03655_);
  and (_18420_, _18419_, _18418_);
  or (_18421_, _18420_, _18417_);
  and (_18423_, _18421_, _04594_);
  and (_18424_, _18366_, _03773_);
  and (_18425_, _18424_, _18418_);
  or (_18426_, _18425_, _03653_);
  or (_18427_, _18426_, _18423_);
  nor (_18428_, _13243_, _08958_);
  or (_18429_, _18354_, _04608_);
  or (_18430_, _18429_, _18428_);
  and (_18431_, _18430_, _04606_);
  and (_18432_, _18431_, _18427_);
  or (_18434_, _18432_, _18358_);
  and (_18435_, _18434_, _04260_);
  and (_18436_, _18363_, _03809_);
  or (_18437_, _18436_, _03816_);
  or (_18438_, _18437_, _18435_);
  and (_18439_, _13425_, _05297_);
  or (_18440_, _18354_, _03820_);
  or (_18441_, _18440_, _18439_);
  and (_18442_, _18441_, _43227_);
  and (_18443_, _18442_, _18438_);
  or (_18445_, _18443_, _18353_);
  and (_43457_, _18445_, _41991_);
  not (_18446_, \oc8051_golden_model_1.IE [0]);
  nor (_18447_, _05337_, _18446_);
  and (_18448_, _12145_, _05337_);
  nor (_18449_, _18448_, _18447_);
  nor (_18450_, _18449_, _04589_);
  and (_18451_, _05337_, _06366_);
  nor (_18452_, _18451_, _18447_);
  and (_18453_, _18452_, _03650_);
  and (_18455_, _05337_, _04491_);
  nor (_18456_, _18455_, _18447_);
  and (_18457_, _18456_, _07441_);
  and (_18458_, _05337_, \oc8051_golden_model_1.ACC [0]);
  nor (_18459_, _18458_, _18447_);
  nor (_18460_, _18459_, _04500_);
  nor (_18461_, _04499_, _18446_);
  or (_18462_, _18461_, _18460_);
  and (_18463_, _18462_, _04515_);
  nor (_18464_, _05744_, _09054_);
  nor (_18466_, _18464_, _18447_);
  nor (_18467_, _18466_, _04515_);
  or (_18468_, _18467_, _18463_);
  and (_18469_, _18468_, _03516_);
  nor (_18470_, _05979_, _18446_);
  and (_18471_, _12035_, _05979_);
  nor (_18472_, _18471_, _18470_);
  nor (_18473_, _18472_, _03516_);
  nor (_18474_, _18473_, _18469_);
  nor (_18475_, _18474_, _03597_);
  nor (_18477_, _18456_, _04524_);
  or (_18478_, _18477_, _18475_);
  and (_18479_, _18478_, _03611_);
  nor (_18480_, _18459_, _03611_);
  or (_18481_, _18480_, _18479_);
  and (_18482_, _18481_, _03512_);
  and (_18483_, _18447_, _03511_);
  or (_18484_, _18483_, _18482_);
  and (_18485_, _18484_, _03505_);
  nor (_18486_, _18466_, _03505_);
  or (_18488_, _18486_, _18485_);
  and (_18489_, _18488_, _03501_);
  nor (_18490_, _12066_, _09091_);
  nor (_18491_, _18490_, _18470_);
  nor (_18492_, _18491_, _03501_);
  or (_18493_, _18492_, _07441_);
  nor (_18494_, _18493_, _18489_);
  nor (_18495_, _18494_, _18457_);
  nor (_18496_, _18495_, _05969_);
  and (_18497_, _06836_, _05337_);
  nor (_18499_, _18447_, _05970_);
  not (_18500_, _18499_);
  nor (_18501_, _18500_, _18497_);
  or (_18502_, _18501_, _03644_);
  nor (_18503_, _18502_, _18496_);
  nor (_18504_, _12129_, _09054_);
  nor (_18505_, _18504_, _18447_);
  nor (_18506_, _18505_, _03275_);
  or (_18507_, _18506_, _03650_);
  nor (_18508_, _18507_, _18503_);
  nor (_18510_, _18508_, _18453_);
  or (_18511_, _18510_, _03649_);
  and (_18512_, _12019_, _05337_);
  or (_18513_, _18512_, _18447_);
  or (_18514_, _18513_, _04591_);
  and (_18515_, _18514_, _04589_);
  and (_18516_, _18515_, _18511_);
  nor (_18517_, _18516_, _18450_);
  nor (_18518_, _18517_, _03655_);
  or (_18519_, _18452_, _04596_);
  nor (_18521_, _18519_, _18464_);
  nor (_18522_, _18521_, _18518_);
  nor (_18523_, _18522_, _03773_);
  and (_18524_, _12144_, _05337_);
  or (_18525_, _18524_, _18447_);
  and (_18526_, _18525_, _03773_);
  or (_18527_, _18526_, _18523_);
  and (_18528_, _18527_, _04608_);
  nor (_18529_, _12017_, _09054_);
  nor (_18530_, _18529_, _18447_);
  nor (_18532_, _18530_, _04608_);
  or (_18533_, _18532_, _18528_);
  and (_18534_, _18533_, _04606_);
  nor (_18535_, _12015_, _09054_);
  nor (_18536_, _18535_, _18447_);
  nor (_18537_, _18536_, _04606_);
  or (_18538_, _18537_, _18534_);
  and (_18539_, _18538_, _04260_);
  nor (_18540_, _18466_, _04260_);
  or (_18541_, _18540_, _18539_);
  and (_18543_, _18541_, _03206_);
  and (_18544_, _18447_, _03205_);
  nor (_18545_, _18544_, _18543_);
  or (_18546_, _18545_, _03816_);
  or (_18547_, _18466_, _03820_);
  and (_18548_, _18547_, _18546_);
  nand (_18549_, _18548_, _43227_);
  or (_18550_, _43227_, \oc8051_golden_model_1.IE [0]);
  and (_18551_, _18550_, _41991_);
  and (_43458_, _18551_, _18549_);
  not (_18553_, _03787_);
  not (_18554_, \oc8051_golden_model_1.IE [1]);
  nor (_18555_, _05337_, _18554_);
  and (_18556_, _06835_, _05337_);
  or (_18557_, _18556_, _18555_);
  and (_18558_, _18557_, _05969_);
  nor (_18559_, _05337_, \oc8051_golden_model_1.IE [1]);
  and (_18560_, _05337_, _03320_);
  nor (_18561_, _18560_, _18559_);
  and (_18562_, _18561_, _04499_);
  nor (_18564_, _04499_, _18554_);
  or (_18565_, _18564_, _18562_);
  and (_18566_, _18565_, _04515_);
  and (_18567_, _12234_, _05337_);
  nor (_18568_, _18567_, _18559_);
  and (_18569_, _18568_, _03599_);
  or (_18570_, _18569_, _18566_);
  and (_18571_, _18570_, _03516_);
  nor (_18572_, _05979_, _18554_);
  and (_18573_, _12238_, _05979_);
  nor (_18575_, _18573_, _18572_);
  nor (_18576_, _18575_, _03516_);
  or (_18577_, _18576_, _18571_);
  and (_18578_, _18577_, _04524_);
  and (_18579_, _05337_, _05898_);
  nor (_18580_, _18579_, _18555_);
  nor (_18581_, _18580_, _04524_);
  or (_18582_, _18581_, _18578_);
  and (_18583_, _18582_, _03611_);
  and (_18584_, _18561_, _03603_);
  or (_18586_, _18584_, _18583_);
  and (_18587_, _18586_, _03512_);
  and (_18588_, _12224_, _05979_);
  nor (_18589_, _18588_, _18572_);
  nor (_18590_, _18589_, _03512_);
  or (_18591_, _18590_, _03504_);
  or (_18592_, _18591_, _18587_);
  and (_18593_, _18573_, _12253_);
  or (_18594_, _18572_, _03505_);
  or (_18595_, _18594_, _18593_);
  and (_18597_, _18595_, _18592_);
  and (_18598_, _18597_, _03501_);
  nor (_18599_, _12270_, _09091_);
  nor (_18600_, _18572_, _18599_);
  nor (_18601_, _18600_, _03501_);
  or (_18602_, _18601_, _07441_);
  nor (_18603_, _18602_, _18598_);
  and (_18604_, _18580_, _07441_);
  or (_18605_, _18604_, _05969_);
  nor (_18606_, _18605_, _18603_);
  or (_18608_, _18606_, _18558_);
  and (_18609_, _18608_, _03275_);
  nor (_18610_, _12330_, _09054_);
  nor (_18611_, _18610_, _18555_);
  nor (_18612_, _18611_, _03275_);
  nor (_18613_, _18612_, _18609_);
  nor (_18614_, _18613_, _08861_);
  not (_18615_, _18559_);
  nor (_18616_, _12220_, _09054_);
  nor (_18617_, _18616_, _04591_);
  and (_18619_, _05337_, _04347_);
  nor (_18620_, _18619_, _04582_);
  or (_18621_, _18620_, _18617_);
  and (_18622_, _18621_, _18615_);
  nor (_18623_, _18622_, _18614_);
  nor (_18624_, _18623_, _03778_);
  nor (_18625_, _12347_, _09054_);
  nor (_18626_, _18625_, _04589_);
  and (_18627_, _18626_, _18615_);
  nor (_18628_, _18627_, _18624_);
  nor (_18630_, _18628_, _03655_);
  nor (_18631_, _12219_, _09054_);
  nor (_18632_, _18631_, _04596_);
  and (_18633_, _18632_, _18615_);
  nor (_18634_, _18633_, _18630_);
  nor (_18635_, _18634_, _03773_);
  nor (_18636_, _18555_, _05699_);
  nor (_18637_, _18636_, _04594_);
  and (_18638_, _18637_, _18561_);
  nor (_18639_, _18638_, _18635_);
  or (_18641_, _18639_, _18553_);
  and (_18642_, _18619_, _05698_);
  nor (_18643_, _18642_, _04608_);
  and (_18644_, _18643_, _18615_);
  and (_18645_, _18560_, _05698_);
  or (_18646_, _18559_, _04606_);
  nor (_18647_, _18646_, _18645_);
  or (_18648_, _18647_, _03809_);
  nor (_18649_, _18648_, _18644_);
  and (_18650_, _18649_, _18641_);
  nor (_18652_, _18568_, _04260_);
  or (_18653_, _18652_, _03205_);
  nor (_18654_, _18653_, _18650_);
  nor (_18655_, _18589_, _03206_);
  or (_18656_, _18655_, _03816_);
  nor (_18657_, _18656_, _18654_);
  or (_18658_, _18555_, _03820_);
  nor (_18659_, _18658_, _18567_);
  nor (_18660_, _18659_, _18657_);
  or (_18661_, _18660_, _43231_);
  or (_18663_, _43227_, \oc8051_golden_model_1.IE [1]);
  and (_18664_, _18663_, _41991_);
  and (_43459_, _18664_, _18661_);
  not (_18665_, \oc8051_golden_model_1.IE [2]);
  nor (_18666_, _05337_, _18665_);
  and (_18667_, _05337_, _06414_);
  nor (_18668_, _18667_, _18666_);
  and (_18669_, _18668_, _03650_);
  nor (_18670_, _09054_, _05130_);
  nor (_18671_, _18670_, _18666_);
  and (_18673_, _18671_, _07441_);
  nor (_18674_, _18671_, _04524_);
  nor (_18675_, _05979_, _18665_);
  and (_18676_, _12416_, _05979_);
  nor (_18677_, _18676_, _18675_);
  and (_18678_, _18677_, _03515_);
  nor (_18679_, _12430_, _09054_);
  nor (_18680_, _18679_, _18666_);
  nor (_18681_, _18680_, _04515_);
  nor (_18682_, _04499_, _18665_);
  and (_18684_, _05337_, \oc8051_golden_model_1.ACC [2]);
  nor (_18685_, _18684_, _18666_);
  nor (_18686_, _18685_, _04500_);
  nor (_18687_, _18686_, _18682_);
  nor (_18688_, _18687_, _03599_);
  or (_18689_, _18688_, _03515_);
  nor (_18690_, _18689_, _18681_);
  nor (_18691_, _18690_, _18678_);
  and (_18692_, _18691_, _04524_);
  or (_18693_, _18692_, _18674_);
  and (_18695_, _18693_, _03611_);
  nor (_18696_, _18685_, _03611_);
  or (_18697_, _18696_, _18695_);
  and (_18698_, _18697_, _03512_);
  and (_18699_, _12414_, _05979_);
  nor (_18700_, _18699_, _18675_);
  nor (_18701_, _18700_, _03512_);
  or (_18702_, _18701_, _03504_);
  or (_18703_, _18702_, _18698_);
  nor (_18704_, _18675_, _12447_);
  nor (_18706_, _18704_, _18677_);
  or (_18707_, _18706_, _03505_);
  and (_18708_, _18707_, _03501_);
  and (_18709_, _18708_, _18703_);
  nor (_18710_, _12465_, _09091_);
  nor (_18711_, _18710_, _18675_);
  nor (_18712_, _18711_, _03501_);
  nor (_18713_, _18712_, _07441_);
  not (_18714_, _18713_);
  nor (_18715_, _18714_, _18709_);
  nor (_18717_, _18715_, _18673_);
  nor (_18718_, _18717_, _05969_);
  and (_18719_, _06839_, _05337_);
  nor (_18720_, _18666_, _05970_);
  not (_18721_, _18720_);
  nor (_18722_, _18721_, _18719_);
  or (_18723_, _18722_, _03644_);
  nor (_18724_, _18723_, _18718_);
  nor (_18725_, _12524_, _09054_);
  nor (_18726_, _18666_, _18725_);
  nor (_18728_, _18726_, _03275_);
  or (_18729_, _18728_, _03650_);
  nor (_18730_, _18729_, _18724_);
  nor (_18731_, _18730_, _18669_);
  or (_18732_, _18731_, _03649_);
  and (_18733_, _12538_, _05337_);
  or (_18734_, _18733_, _18666_);
  or (_18735_, _18734_, _04591_);
  and (_18736_, _18735_, _04589_);
  and (_18737_, _18736_, _18732_);
  and (_18739_, _12544_, _05337_);
  nor (_18740_, _18739_, _18666_);
  nor (_18741_, _18740_, _04589_);
  nor (_18742_, _18741_, _18737_);
  nor (_18743_, _18742_, _03655_);
  nor (_18744_, _18666_, _05793_);
  not (_18745_, _18744_);
  nor (_18746_, _18668_, _04596_);
  and (_18747_, _18746_, _18745_);
  nor (_18748_, _18747_, _18743_);
  nor (_18750_, _18748_, _03773_);
  nor (_18751_, _18685_, _04594_);
  and (_18752_, _18751_, _18745_);
  or (_18753_, _18752_, _18750_);
  and (_18754_, _18753_, _04608_);
  nor (_18755_, _12537_, _09054_);
  nor (_18756_, _18755_, _18666_);
  nor (_18757_, _18756_, _04608_);
  or (_18758_, _18757_, _18754_);
  and (_18759_, _18758_, _04606_);
  nor (_18761_, _12543_, _09054_);
  nor (_18762_, _18761_, _18666_);
  nor (_18763_, _18762_, _04606_);
  or (_18764_, _18763_, _18759_);
  and (_18765_, _18764_, _04260_);
  nor (_18766_, _18680_, _04260_);
  or (_18767_, _18766_, _18765_);
  and (_18768_, _18767_, _03206_);
  nor (_18769_, _18700_, _03206_);
  or (_18770_, _18769_, _18768_);
  and (_18772_, _18770_, _03820_);
  and (_18773_, _12600_, _05337_);
  nor (_18774_, _18773_, _18666_);
  nor (_18775_, _18774_, _03820_);
  or (_18776_, _18775_, _18772_);
  or (_18777_, _18776_, _43231_);
  or (_18778_, _43227_, \oc8051_golden_model_1.IE [2]);
  and (_18779_, _18778_, _41991_);
  and (_43460_, _18779_, _18777_);
  not (_18780_, \oc8051_golden_model_1.IE [3]);
  nor (_18782_, _05337_, _18780_);
  and (_18783_, _05337_, _06347_);
  nor (_18784_, _18783_, _18782_);
  and (_18785_, _18784_, _03650_);
  nor (_18786_, _09054_, _04944_);
  nor (_18787_, _18786_, _18782_);
  and (_18788_, _18787_, _07441_);
  and (_18789_, _05337_, \oc8051_golden_model_1.ACC [3]);
  nor (_18790_, _18789_, _18782_);
  nor (_18791_, _18790_, _04500_);
  nor (_18793_, _04499_, _18780_);
  or (_18794_, _18793_, _18791_);
  and (_18795_, _18794_, _04515_);
  nor (_18796_, _12625_, _09054_);
  nor (_18797_, _18796_, _18782_);
  nor (_18798_, _18797_, _04515_);
  or (_18799_, _18798_, _18795_);
  and (_18800_, _18799_, _03516_);
  nor (_18801_, _05979_, _18780_);
  and (_18802_, _12638_, _05979_);
  nor (_18804_, _18802_, _18801_);
  nor (_18805_, _18804_, _03516_);
  or (_18806_, _18805_, _03597_);
  or (_18807_, _18806_, _18800_);
  nand (_18808_, _18787_, _03597_);
  and (_18809_, _18808_, _18807_);
  and (_18810_, _18809_, _03611_);
  nor (_18811_, _18790_, _03611_);
  or (_18812_, _18811_, _18810_);
  and (_18813_, _18812_, _03512_);
  and (_18815_, _12622_, _05979_);
  nor (_18816_, _18815_, _18801_);
  nor (_18817_, _18816_, _03512_);
  or (_18818_, _18817_, _03504_);
  or (_18819_, _18818_, _18813_);
  nor (_18820_, _18801_, _12653_);
  nor (_18821_, _18820_, _18804_);
  or (_18822_, _18821_, _03505_);
  and (_18823_, _18822_, _03501_);
  and (_18824_, _18823_, _18819_);
  nor (_18826_, _12671_, _09091_);
  nor (_18827_, _18826_, _18801_);
  nor (_18828_, _18827_, _03501_);
  nor (_18829_, _18828_, _07441_);
  not (_18830_, _18829_);
  nor (_18831_, _18830_, _18824_);
  nor (_18832_, _18831_, _18788_);
  nor (_18833_, _18832_, _05969_);
  and (_18834_, _06838_, _05337_);
  nor (_18835_, _18782_, _05970_);
  not (_18837_, _18835_);
  nor (_18838_, _18837_, _18834_);
  or (_18839_, _18838_, _03644_);
  nor (_18840_, _18839_, _18833_);
  nor (_18841_, _12731_, _09054_);
  nor (_18842_, _18782_, _18841_);
  nor (_18843_, _18842_, _03275_);
  or (_18844_, _18843_, _03650_);
  nor (_18845_, _18844_, _18840_);
  nor (_18846_, _18845_, _18785_);
  or (_18848_, _18846_, _03649_);
  and (_18849_, _12746_, _05337_);
  or (_18850_, _18849_, _18782_);
  or (_18851_, _18850_, _04591_);
  and (_18852_, _18851_, _04589_);
  and (_18853_, _18852_, _18848_);
  and (_18854_, _12619_, _05337_);
  nor (_18855_, _18854_, _18782_);
  nor (_18856_, _18855_, _04589_);
  nor (_18857_, _18856_, _18853_);
  nor (_18859_, _18857_, _03655_);
  nor (_18860_, _18782_, _05650_);
  not (_18861_, _18860_);
  nor (_18862_, _18784_, _04596_);
  and (_18863_, _18862_, _18861_);
  nor (_18864_, _18863_, _18859_);
  nor (_18865_, _18864_, _03773_);
  nor (_18866_, _18790_, _04594_);
  and (_18867_, _18866_, _18861_);
  nor (_18868_, _18867_, _03653_);
  not (_18870_, _18868_);
  nor (_18871_, _18870_, _18865_);
  nor (_18872_, _12745_, _09054_);
  or (_18873_, _18782_, _04608_);
  nor (_18874_, _18873_, _18872_);
  or (_18875_, _18874_, _03786_);
  nor (_18876_, _18875_, _18871_);
  nor (_18877_, _12618_, _09054_);
  nor (_18878_, _18877_, _18782_);
  nor (_18879_, _18878_, _04606_);
  or (_18881_, _18879_, _18876_);
  and (_18882_, _18881_, _04260_);
  nor (_18883_, _18797_, _04260_);
  or (_18884_, _18883_, _18882_);
  and (_18885_, _18884_, _03206_);
  nor (_18886_, _18816_, _03206_);
  or (_18887_, _18886_, _18885_);
  and (_18888_, _18887_, _03820_);
  and (_18889_, _12806_, _05337_);
  nor (_18890_, _18889_, _18782_);
  nor (_18892_, _18890_, _03820_);
  or (_18893_, _18892_, _18888_);
  or (_18894_, _18893_, _43231_);
  or (_18895_, _43227_, \oc8051_golden_model_1.IE [3]);
  and (_18896_, _18895_, _41991_);
  and (_43461_, _18896_, _18894_);
  not (_18897_, \oc8051_golden_model_1.IE [4]);
  nor (_18898_, _05337_, _18897_);
  nor (_18899_, _05840_, _09054_);
  nor (_18900_, _18899_, _18898_);
  and (_18902_, _18900_, _07441_);
  nor (_18903_, _05979_, _18897_);
  and (_18904_, _12853_, _05979_);
  nor (_18905_, _18904_, _18903_);
  nor (_18906_, _18905_, _03512_);
  and (_18907_, _05337_, \oc8051_golden_model_1.ACC [4]);
  nor (_18908_, _18907_, _18898_);
  nor (_18909_, _18908_, _04500_);
  nor (_18910_, _04499_, _18897_);
  or (_18911_, _18910_, _18909_);
  and (_18913_, _18911_, _04515_);
  nor (_18914_, _12820_, _09054_);
  nor (_18915_, _18914_, _18898_);
  nor (_18916_, _18915_, _04515_);
  or (_18917_, _18916_, _18913_);
  and (_18918_, _18917_, _03516_);
  and (_18919_, _12830_, _05979_);
  nor (_18920_, _18919_, _18903_);
  nor (_18921_, _18920_, _03516_);
  or (_18922_, _18921_, _03597_);
  or (_18924_, _18922_, _18918_);
  nand (_18925_, _18900_, _03597_);
  and (_18926_, _18925_, _18924_);
  and (_18927_, _18926_, _03611_);
  nor (_18928_, _18908_, _03611_);
  or (_18929_, _18928_, _18927_);
  and (_18930_, _18929_, _03512_);
  nor (_18931_, _18930_, _18906_);
  nor (_18932_, _18931_, _03504_);
  and (_18933_, _12861_, _05979_);
  nor (_18935_, _18933_, _18903_);
  nor (_18936_, _18935_, _03505_);
  nor (_18937_, _18936_, _18932_);
  nor (_18938_, _18937_, _03500_);
  nor (_18939_, _12828_, _09091_);
  nor (_18940_, _18939_, _18903_);
  nor (_18941_, _18940_, _03501_);
  nor (_18942_, _18941_, _07441_);
  not (_18943_, _18942_);
  nor (_18944_, _18943_, _18938_);
  nor (_18946_, _18944_, _18902_);
  nor (_18947_, _18946_, _05969_);
  and (_18948_, _06843_, _05337_);
  nor (_18949_, _18898_, _05970_);
  not (_18950_, _18949_);
  nor (_18951_, _18950_, _18948_);
  nor (_18952_, _18951_, _03644_);
  not (_18953_, _18952_);
  nor (_18954_, _18953_, _18947_);
  nor (_18955_, _12936_, _09054_);
  nor (_18957_, _18955_, _18898_);
  nor (_18958_, _18957_, _03275_);
  or (_18959_, _18958_, _08861_);
  or (_18960_, _18959_, _18954_);
  and (_18961_, _12951_, _05337_);
  or (_18962_, _18898_, _04591_);
  or (_18963_, _18962_, _18961_);
  and (_18964_, _06375_, _05337_);
  nor (_18965_, _18964_, _18898_);
  and (_18966_, _18965_, _03650_);
  nor (_18968_, _18966_, _03778_);
  and (_18969_, _18968_, _18963_);
  and (_18970_, _18969_, _18960_);
  and (_18971_, _12957_, _05337_);
  nor (_18972_, _18971_, _18898_);
  nor (_18973_, _18972_, _04589_);
  nor (_18974_, _18973_, _18970_);
  nor (_18975_, _18974_, _03655_);
  nor (_18976_, _18898_, _05889_);
  not (_18977_, _18976_);
  nor (_18979_, _18965_, _04596_);
  and (_18980_, _18979_, _18977_);
  nor (_18981_, _18980_, _18975_);
  nor (_18982_, _18981_, _03773_);
  nor (_18983_, _18908_, _04594_);
  and (_18984_, _18983_, _18977_);
  or (_18985_, _18984_, _18982_);
  and (_18986_, _18985_, _04608_);
  nor (_18987_, _12949_, _09054_);
  nor (_18988_, _18987_, _18898_);
  nor (_18990_, _18988_, _04608_);
  or (_18991_, _18990_, _18986_);
  and (_18992_, _18991_, _04606_);
  nor (_18993_, _12956_, _09054_);
  nor (_18994_, _18993_, _18898_);
  nor (_18995_, _18994_, _04606_);
  or (_18996_, _18995_, _18992_);
  and (_18997_, _18996_, _04260_);
  nor (_18998_, _18915_, _04260_);
  or (_18999_, _18998_, _18997_);
  and (_19001_, _18999_, _03206_);
  nor (_19002_, _18905_, _03206_);
  or (_19003_, _19002_, _19001_);
  and (_19004_, _19003_, _03820_);
  and (_19005_, _13013_, _05337_);
  nor (_19006_, _19005_, _18898_);
  nor (_19007_, _19006_, _03820_);
  or (_19008_, _19007_, _19004_);
  or (_19009_, _19008_, _43231_);
  or (_19010_, _43227_, \oc8051_golden_model_1.IE [4]);
  and (_19012_, _19010_, _41991_);
  and (_43462_, _19012_, _19009_);
  not (_19013_, \oc8051_golden_model_1.IE [5]);
  nor (_19014_, _05337_, _19013_);
  and (_19015_, _06842_, _05337_);
  or (_19016_, _19015_, _19014_);
  and (_19017_, _19016_, _05969_);
  and (_19018_, _05337_, \oc8051_golden_model_1.ACC [5]);
  nor (_19019_, _19018_, _19014_);
  nor (_19020_, _19019_, _04500_);
  nor (_19022_, _04499_, _19013_);
  or (_19023_, _19022_, _19020_);
  and (_19024_, _19023_, _04515_);
  nor (_19025_, _13035_, _09054_);
  nor (_19026_, _19025_, _19014_);
  nor (_19027_, _19026_, _04515_);
  or (_19028_, _19027_, _19024_);
  and (_19029_, _19028_, _03516_);
  nor (_19030_, _05979_, _19013_);
  and (_19031_, _13051_, _05979_);
  nor (_19033_, _19031_, _19030_);
  nor (_19034_, _19033_, _03516_);
  or (_19035_, _19034_, _03597_);
  or (_19036_, _19035_, _19029_);
  nor (_19037_, _05552_, _09054_);
  nor (_19038_, _19037_, _19014_);
  nand (_19039_, _19038_, _03597_);
  and (_19040_, _19039_, _19036_);
  and (_19041_, _19040_, _03611_);
  nor (_19042_, _19019_, _03611_);
  or (_19044_, _19042_, _19041_);
  and (_19045_, _19044_, _03512_);
  and (_19046_, _13032_, _05979_);
  nor (_19047_, _19046_, _19030_);
  nor (_19048_, _19047_, _03512_);
  or (_19049_, _19048_, _03504_);
  or (_19050_, _19049_, _19045_);
  nor (_19051_, _19030_, _13066_);
  nor (_19052_, _19051_, _19033_);
  or (_19053_, _19052_, _03505_);
  and (_19055_, _19053_, _03501_);
  and (_19056_, _19055_, _19050_);
  nor (_19057_, _13030_, _09091_);
  nor (_19058_, _19057_, _19030_);
  nor (_19059_, _19058_, _03501_);
  nor (_19060_, _19059_, _07441_);
  not (_19061_, _19060_);
  nor (_19062_, _19061_, _19056_);
  and (_19063_, _19038_, _07441_);
  or (_19064_, _19063_, _05969_);
  nor (_19066_, _19064_, _19062_);
  or (_19067_, _19066_, _19017_);
  and (_19068_, _19067_, _03275_);
  nor (_19069_, _13139_, _09054_);
  nor (_19070_, _19069_, _19014_);
  nor (_19071_, _19070_, _03275_);
  or (_19072_, _19071_, _08861_);
  or (_19073_, _19072_, _19068_);
  and (_19074_, _13154_, _05337_);
  or (_19075_, _19014_, _04591_);
  or (_19077_, _19075_, _19074_);
  and (_19078_, _06358_, _05337_);
  nor (_19079_, _19078_, _19014_);
  and (_19080_, _19079_, _03650_);
  nor (_19081_, _19080_, _03778_);
  and (_19082_, _19081_, _19077_);
  and (_19083_, _19082_, _19073_);
  and (_19084_, _13160_, _05337_);
  nor (_19085_, _19084_, _19014_);
  nor (_19086_, _19085_, _04589_);
  nor (_19088_, _19086_, _19083_);
  nor (_19089_, _19088_, _03655_);
  nor (_19090_, _19014_, _05601_);
  not (_19091_, _19090_);
  nor (_19092_, _19079_, _04596_);
  and (_19093_, _19092_, _19091_);
  nor (_19094_, _19093_, _19089_);
  nor (_19095_, _19094_, _03773_);
  nor (_19096_, _19019_, _04594_);
  and (_19097_, _19096_, _19091_);
  or (_19099_, _19097_, _19095_);
  and (_19100_, _19099_, _04608_);
  nor (_19101_, _13152_, _09054_);
  nor (_19102_, _19101_, _19014_);
  nor (_19103_, _19102_, _04608_);
  or (_19104_, _19103_, _19100_);
  and (_19105_, _19104_, _04606_);
  nor (_19106_, _13159_, _09054_);
  nor (_19107_, _19106_, _19014_);
  nor (_19108_, _19107_, _04606_);
  or (_19110_, _19108_, _19105_);
  and (_19111_, _19110_, _04260_);
  nor (_19112_, _19026_, _04260_);
  or (_19113_, _19112_, _19111_);
  and (_19114_, _19113_, _03206_);
  nor (_19115_, _19047_, _03206_);
  or (_19116_, _19115_, _19114_);
  and (_19117_, _19116_, _03820_);
  and (_19118_, _13217_, _05337_);
  nor (_19119_, _19118_, _19014_);
  nor (_19121_, _19119_, _03820_);
  or (_19122_, _19121_, _19117_);
  or (_19123_, _19122_, _43231_);
  or (_19124_, _43227_, \oc8051_golden_model_1.IE [5]);
  and (_19125_, _19124_, _41991_);
  and (_43463_, _19125_, _19123_);
  not (_19126_, \oc8051_golden_model_1.IE [6]);
  nor (_19127_, _05337_, _19126_);
  and (_19128_, _06531_, _05337_);
  or (_19129_, _19128_, _19127_);
  and (_19131_, _19129_, _05969_);
  and (_19132_, _05337_, \oc8051_golden_model_1.ACC [6]);
  nor (_19133_, _19132_, _19127_);
  nor (_19134_, _19133_, _04500_);
  nor (_19135_, _04499_, _19126_);
  or (_19136_, _19135_, _19134_);
  and (_19137_, _19136_, _04515_);
  nor (_19138_, _13235_, _09054_);
  nor (_19139_, _19138_, _19127_);
  nor (_19140_, _19139_, _04515_);
  or (_19142_, _19140_, _19137_);
  and (_19143_, _19142_, _03516_);
  nor (_19144_, _05979_, _19126_);
  and (_19145_, _13266_, _05979_);
  nor (_19146_, _19145_, _19144_);
  nor (_19147_, _19146_, _03516_);
  or (_19148_, _19147_, _03597_);
  or (_19149_, _19148_, _19143_);
  nor (_19150_, _05442_, _09054_);
  nor (_19151_, _19150_, _19127_);
  nand (_19153_, _19151_, _03597_);
  and (_19154_, _19153_, _19149_);
  and (_19155_, _19154_, _03611_);
  nor (_19156_, _19133_, _03611_);
  or (_19157_, _19156_, _19155_);
  and (_19158_, _19157_, _03512_);
  and (_19159_, _13251_, _05979_);
  nor (_19160_, _19159_, _19144_);
  nor (_19161_, _19160_, _03512_);
  or (_19162_, _19161_, _19158_);
  and (_19164_, _19162_, _03505_);
  nor (_19165_, _19144_, _13281_);
  nor (_19166_, _19165_, _19146_);
  and (_19167_, _19166_, _03504_);
  or (_19168_, _19167_, _19164_);
  and (_19169_, _19168_, _03501_);
  nor (_19170_, _13249_, _09091_);
  nor (_19171_, _19170_, _19144_);
  nor (_19172_, _19171_, _03501_);
  nor (_19173_, _19172_, _07441_);
  not (_19175_, _19173_);
  nor (_19176_, _19175_, _19169_);
  and (_19177_, _19151_, _07441_);
  or (_19178_, _19177_, _05969_);
  nor (_19179_, _19178_, _19176_);
  or (_19180_, _19179_, _19131_);
  and (_19181_, _19180_, _03275_);
  nor (_19182_, _13356_, _09054_);
  nor (_19183_, _19182_, _19127_);
  nor (_19184_, _19183_, _03275_);
  or (_19186_, _19184_, _08861_);
  or (_19187_, _19186_, _19181_);
  and (_19188_, _13245_, _05337_);
  or (_19189_, _19127_, _04591_);
  or (_19190_, _19189_, _19188_);
  and (_19191_, _13363_, _05337_);
  nor (_19192_, _19191_, _19127_);
  and (_19193_, _19192_, _03650_);
  nor (_19194_, _19193_, _03778_);
  and (_19195_, _19194_, _19190_);
  and (_19197_, _19195_, _19187_);
  and (_19198_, _13374_, _05337_);
  nor (_19199_, _19198_, _19127_);
  nor (_19200_, _19199_, _04589_);
  nor (_19201_, _19200_, _19197_);
  nor (_19202_, _19201_, _03655_);
  nor (_19203_, _19127_, _05491_);
  not (_19204_, _19203_);
  nor (_19205_, _19192_, _04596_);
  and (_19206_, _19205_, _19204_);
  nor (_19208_, _19206_, _19202_);
  nor (_19209_, _19208_, _03773_);
  nor (_19210_, _19133_, _04594_);
  and (_19211_, _19210_, _19204_);
  nor (_19212_, _19211_, _03653_);
  not (_19213_, _19212_);
  nor (_19214_, _19213_, _19209_);
  nor (_19215_, _13243_, _09054_);
  or (_19216_, _19127_, _04608_);
  nor (_19217_, _19216_, _19215_);
  or (_19219_, _19217_, _03786_);
  nor (_19220_, _19219_, _19214_);
  nor (_19221_, _13373_, _09054_);
  nor (_19222_, _19221_, _19127_);
  nor (_19223_, _19222_, _04606_);
  or (_19224_, _19223_, _19220_);
  and (_19225_, _19224_, _04260_);
  nor (_19226_, _19139_, _04260_);
  or (_19227_, _19226_, _19225_);
  and (_19228_, _19227_, _03206_);
  nor (_19230_, _19160_, _03206_);
  or (_19231_, _19230_, _19228_);
  and (_19232_, _19231_, _03820_);
  and (_19233_, _13425_, _05337_);
  nor (_19234_, _19233_, _19127_);
  nor (_19235_, _19234_, _03820_);
  or (_19236_, _19235_, _19232_);
  or (_19237_, _19236_, _43231_);
  or (_19238_, _43227_, \oc8051_golden_model_1.IE [6]);
  and (_19239_, _19238_, _41991_);
  and (_43464_, _19239_, _19237_);
  not (_19241_, \oc8051_golden_model_1.IP [0]);
  nor (_19242_, _05376_, _19241_);
  and (_19243_, _12145_, _05376_);
  nor (_19244_, _19243_, _19242_);
  nor (_19245_, _19244_, _04589_);
  and (_19246_, _05376_, _06366_);
  nor (_19247_, _19246_, _19242_);
  and (_19248_, _19247_, _03650_);
  and (_19249_, _05376_, _04491_);
  nor (_19251_, _19249_, _19242_);
  and (_19252_, _19251_, _07441_);
  and (_19253_, _05376_, \oc8051_golden_model_1.ACC [0]);
  nor (_19254_, _19253_, _19242_);
  nor (_19255_, _19254_, _04500_);
  nor (_19256_, _04499_, _19241_);
  or (_19257_, _19256_, _19255_);
  and (_19258_, _19257_, _04515_);
  nor (_19259_, _05744_, _09161_);
  nor (_19260_, _19259_, _19242_);
  nor (_19262_, _19260_, _04515_);
  or (_19263_, _19262_, _19258_);
  and (_19264_, _19263_, _03516_);
  nor (_19265_, _05989_, _19241_);
  and (_19266_, _12035_, _05989_);
  nor (_19267_, _19266_, _19265_);
  nor (_19268_, _19267_, _03516_);
  nor (_19269_, _19268_, _19264_);
  nor (_19270_, _19269_, _03597_);
  nor (_19271_, _19251_, _04524_);
  or (_19273_, _19271_, _19270_);
  and (_19274_, _19273_, _03611_);
  nor (_19275_, _19254_, _03611_);
  or (_19276_, _19275_, _19274_);
  and (_19277_, _19276_, _03512_);
  and (_19278_, _19242_, _03511_);
  or (_19279_, _19278_, _19277_);
  and (_19280_, _19279_, _03505_);
  nor (_19281_, _19260_, _03505_);
  or (_19282_, _19281_, _19280_);
  and (_19284_, _19282_, _03501_);
  nor (_19285_, _12066_, _09198_);
  nor (_19286_, _19285_, _19265_);
  nor (_19287_, _19286_, _03501_);
  or (_19288_, _19287_, _07441_);
  nor (_19289_, _19288_, _19284_);
  nor (_19290_, _19289_, _19252_);
  nor (_19291_, _19290_, _05969_);
  and (_19292_, _06836_, _05376_);
  nor (_19293_, _19242_, _05970_);
  not (_19295_, _19293_);
  nor (_19296_, _19295_, _19292_);
  or (_19297_, _19296_, _03644_);
  nor (_19298_, _19297_, _19291_);
  nor (_19299_, _12129_, _09161_);
  nor (_19300_, _19299_, _19242_);
  nor (_19301_, _19300_, _03275_);
  or (_19302_, _19301_, _03650_);
  nor (_19303_, _19302_, _19298_);
  nor (_19304_, _19303_, _19248_);
  or (_19306_, _19304_, _03649_);
  and (_19307_, _12019_, _05376_);
  or (_19308_, _19307_, _19242_);
  or (_19309_, _19308_, _04591_);
  and (_19310_, _19309_, _04589_);
  and (_19311_, _19310_, _19306_);
  nor (_19312_, _19311_, _19245_);
  nor (_19313_, _19312_, _03655_);
  or (_19314_, _19247_, _04596_);
  nor (_19315_, _19314_, _19259_);
  nor (_19317_, _19315_, _19313_);
  nor (_19318_, _19317_, _03773_);
  and (_19319_, _12144_, _05376_);
  or (_19320_, _19319_, _19242_);
  and (_19321_, _19320_, _03773_);
  or (_19322_, _19321_, _19318_);
  and (_19323_, _19322_, _04608_);
  nor (_19324_, _12017_, _09161_);
  nor (_19325_, _19324_, _19242_);
  nor (_19326_, _19325_, _04608_);
  or (_19328_, _19326_, _19323_);
  and (_19329_, _19328_, _04606_);
  nor (_19330_, _12015_, _09161_);
  nor (_19331_, _19330_, _19242_);
  nor (_19332_, _19331_, _04606_);
  or (_19333_, _19332_, _19329_);
  and (_19334_, _19333_, _04260_);
  nor (_19335_, _19260_, _04260_);
  or (_19336_, _19335_, _19334_);
  and (_19337_, _19336_, _03206_);
  and (_19339_, _19242_, _03205_);
  nor (_19340_, _19339_, _03816_);
  not (_19341_, _19340_);
  nor (_19342_, _19341_, _19337_);
  and (_19343_, _19260_, _03816_);
  or (_19344_, _19343_, _19342_);
  nand (_19345_, _19344_, _43227_);
  or (_19346_, _43227_, \oc8051_golden_model_1.IP [0]);
  and (_19347_, _19346_, _41991_);
  and (_43467_, _19347_, _19345_);
  not (_19349_, \oc8051_golden_model_1.IP [1]);
  nor (_19350_, _05376_, _19349_);
  and (_19351_, _06835_, _05376_);
  or (_19352_, _19351_, _19350_);
  and (_19353_, _19352_, _05969_);
  nor (_19354_, _05376_, \oc8051_golden_model_1.IP [1]);
  and (_19355_, _05376_, _03320_);
  nor (_19356_, _19355_, _19354_);
  and (_19357_, _19356_, _04499_);
  nor (_19358_, _04499_, _19349_);
  or (_19360_, _19358_, _19357_);
  and (_19361_, _19360_, _04515_);
  and (_19362_, _12234_, _05376_);
  nor (_19363_, _19362_, _19354_);
  and (_19364_, _19363_, _03599_);
  or (_19365_, _19364_, _19361_);
  and (_19366_, _19365_, _03516_);
  nor (_19367_, _05989_, _19349_);
  and (_19368_, _12238_, _05989_);
  nor (_19369_, _19368_, _19367_);
  nor (_19371_, _19369_, _03516_);
  or (_19372_, _19371_, _19366_);
  and (_19373_, _19372_, _04524_);
  and (_19374_, _05376_, _05898_);
  nor (_19375_, _19374_, _19350_);
  nor (_19376_, _19375_, _04524_);
  or (_19377_, _19376_, _19373_);
  and (_19378_, _19377_, _03611_);
  and (_19379_, _19356_, _03603_);
  or (_19380_, _19379_, _19378_);
  and (_19382_, _19380_, _03512_);
  and (_19383_, _12224_, _05989_);
  nor (_19384_, _19383_, _19367_);
  nor (_19385_, _19384_, _03512_);
  or (_19386_, _19385_, _19382_);
  and (_19387_, _19386_, _03505_);
  and (_19388_, _19368_, _12253_);
  or (_19389_, _19388_, _19367_);
  and (_19390_, _19389_, _03504_);
  or (_19391_, _19390_, _19387_);
  and (_19393_, _19391_, _03501_);
  nor (_19394_, _12270_, _09198_);
  nor (_19395_, _19367_, _19394_);
  nor (_19396_, _19395_, _03501_);
  or (_19397_, _19396_, _07441_);
  nor (_19398_, _19397_, _19393_);
  and (_19399_, _19375_, _07441_);
  or (_19400_, _19399_, _05969_);
  nor (_19401_, _19400_, _19398_);
  or (_19402_, _19401_, _19353_);
  and (_19404_, _19402_, _03275_);
  nor (_19405_, _12330_, _09161_);
  nor (_19406_, _19405_, _19350_);
  nor (_19407_, _19406_, _03275_);
  nor (_19408_, _19407_, _19404_);
  nor (_19409_, _19408_, _08861_);
  not (_19410_, _19354_);
  nor (_19411_, _12220_, _09161_);
  nor (_19412_, _19411_, _04591_);
  and (_19413_, _05376_, _04347_);
  nor (_19415_, _19413_, _04582_);
  or (_19416_, _19415_, _19412_);
  and (_19417_, _19416_, _19410_);
  nor (_19418_, _19417_, _19409_);
  nor (_19419_, _19418_, _03778_);
  nor (_19420_, _12347_, _09161_);
  nor (_19421_, _19420_, _04589_);
  and (_19422_, _19421_, _19410_);
  nor (_19423_, _19422_, _19419_);
  nor (_19424_, _19423_, _03655_);
  nor (_19426_, _12219_, _09161_);
  nor (_19427_, _19426_, _04596_);
  and (_19428_, _19427_, _19410_);
  nor (_19429_, _19428_, _19424_);
  nor (_19430_, _19429_, _03773_);
  nor (_19431_, _19350_, _05699_);
  nor (_19432_, _19431_, _04594_);
  and (_19433_, _19432_, _19356_);
  nor (_19434_, _19433_, _19430_);
  or (_19435_, _19434_, _18553_);
  and (_19437_, _19413_, _05698_);
  or (_19438_, _19354_, _04608_);
  or (_19439_, _19438_, _19437_);
  and (_19440_, _19355_, _05698_);
  or (_19441_, _19354_, _04606_);
  or (_19442_, _19441_, _19440_);
  and (_19443_, _19442_, _04260_);
  and (_19444_, _19443_, _19439_);
  and (_19445_, _19444_, _19435_);
  nor (_19446_, _19363_, _04260_);
  or (_19448_, _19446_, _03205_);
  nor (_19449_, _19448_, _19445_);
  nor (_19450_, _19384_, _03206_);
  or (_19451_, _19450_, _03816_);
  nor (_19452_, _19451_, _19449_);
  or (_19453_, _19350_, _03820_);
  nor (_19454_, _19453_, _19362_);
  nor (_19455_, _19454_, _19452_);
  or (_19456_, _19455_, _43231_);
  or (_19457_, _43227_, \oc8051_golden_model_1.IP [1]);
  and (_19459_, _19457_, _41991_);
  and (_43468_, _19459_, _19456_);
  not (_19460_, \oc8051_golden_model_1.IP [2]);
  nor (_19461_, _05376_, _19460_);
  and (_19462_, _05376_, _06414_);
  nor (_19463_, _19462_, _19461_);
  and (_19464_, _19463_, _03650_);
  nor (_19465_, _09161_, _05130_);
  nor (_19466_, _19465_, _19461_);
  and (_19467_, _19466_, _07441_);
  and (_19469_, _05376_, \oc8051_golden_model_1.ACC [2]);
  nor (_19470_, _19469_, _19461_);
  nor (_19471_, _19470_, _04500_);
  nor (_19472_, _04499_, _19460_);
  or (_19473_, _19472_, _19471_);
  and (_19474_, _19473_, _04515_);
  nor (_19475_, _12430_, _09161_);
  nor (_19476_, _19475_, _19461_);
  nor (_19477_, _19476_, _04515_);
  or (_19478_, _19477_, _19474_);
  and (_19480_, _19478_, _03516_);
  nor (_19481_, _05989_, _19460_);
  and (_19482_, _12416_, _05989_);
  nor (_19483_, _19482_, _19481_);
  nor (_19484_, _19483_, _03516_);
  or (_19485_, _19484_, _19480_);
  and (_19486_, _19485_, _04524_);
  nor (_19487_, _19466_, _04524_);
  or (_19488_, _19487_, _19486_);
  and (_19489_, _19488_, _03611_);
  nor (_19491_, _19470_, _03611_);
  or (_19492_, _19491_, _19489_);
  and (_19493_, _19492_, _03512_);
  and (_19494_, _12414_, _05989_);
  nor (_19495_, _19494_, _19481_);
  nor (_19496_, _19495_, _03512_);
  or (_19497_, _19496_, _03504_);
  or (_19498_, _19497_, _19493_);
  and (_19499_, _19482_, _12447_);
  or (_19500_, _19481_, _03505_);
  or (_19502_, _19500_, _19499_);
  and (_19503_, _19502_, _03501_);
  and (_19504_, _19503_, _19498_);
  nor (_19505_, _12465_, _09198_);
  nor (_19506_, _19505_, _19481_);
  nor (_19507_, _19506_, _03501_);
  nor (_19508_, _19507_, _07441_);
  not (_19509_, _19508_);
  nor (_19510_, _19509_, _19504_);
  nor (_19511_, _19510_, _19467_);
  nor (_19513_, _19511_, _05969_);
  and (_19514_, _06839_, _05376_);
  nor (_19515_, _19461_, _05970_);
  not (_19516_, _19515_);
  nor (_19517_, _19516_, _19514_);
  or (_19518_, _19517_, _03644_);
  nor (_19519_, _19518_, _19513_);
  nor (_19520_, _12524_, _09161_);
  nor (_19521_, _19461_, _19520_);
  nor (_19522_, _19521_, _03275_);
  or (_19524_, _19522_, _03650_);
  nor (_19525_, _19524_, _19519_);
  nor (_19526_, _19525_, _19464_);
  or (_19527_, _19526_, _03649_);
  and (_19528_, _12538_, _05376_);
  or (_19529_, _19528_, _19461_);
  or (_19530_, _19529_, _04591_);
  and (_19531_, _19530_, _04589_);
  and (_19532_, _19531_, _19527_);
  and (_19533_, _12544_, _05376_);
  nor (_19535_, _19533_, _19461_);
  nor (_19536_, _19535_, _04589_);
  nor (_19537_, _19536_, _19532_);
  nor (_19538_, _19537_, _03655_);
  nor (_19539_, _19461_, _05793_);
  not (_19540_, _19539_);
  nor (_19541_, _19463_, _04596_);
  and (_19542_, _19541_, _19540_);
  nor (_19543_, _19542_, _19538_);
  nor (_19544_, _19543_, _03773_);
  nor (_19546_, _19470_, _04594_);
  and (_19547_, _19546_, _19540_);
  nor (_19548_, _19547_, _03653_);
  not (_19549_, _19548_);
  nor (_19550_, _19549_, _19544_);
  nor (_19551_, _12537_, _09161_);
  or (_19552_, _19461_, _04608_);
  nor (_19553_, _19552_, _19551_);
  or (_19554_, _19553_, _03786_);
  nor (_19555_, _19554_, _19550_);
  nor (_19557_, _12543_, _09161_);
  nor (_19558_, _19557_, _19461_);
  nor (_19559_, _19558_, _04606_);
  or (_19560_, _19559_, _19555_);
  and (_19561_, _19560_, _04260_);
  nor (_19562_, _19476_, _04260_);
  or (_19563_, _19562_, _19561_);
  and (_19564_, _19563_, _03206_);
  nor (_19565_, _19495_, _03206_);
  or (_19566_, _19565_, _19564_);
  and (_19568_, _19566_, _03820_);
  and (_19569_, _12600_, _05376_);
  nor (_19570_, _19569_, _19461_);
  nor (_19571_, _19570_, _03820_);
  or (_19572_, _19571_, _19568_);
  or (_19573_, _19572_, _43231_);
  or (_19574_, _43227_, \oc8051_golden_model_1.IP [2]);
  and (_19575_, _19574_, _41991_);
  and (_43469_, _19575_, _19573_);
  not (_19576_, \oc8051_golden_model_1.IP [3]);
  nor (_19578_, _05376_, _19576_);
  and (_19579_, _05376_, _06347_);
  nor (_19580_, _19579_, _19578_);
  and (_19581_, _19580_, _03650_);
  nor (_19582_, _09161_, _04944_);
  nor (_19583_, _19582_, _19578_);
  and (_19584_, _19583_, _07441_);
  and (_19585_, _05376_, \oc8051_golden_model_1.ACC [3]);
  nor (_19586_, _19585_, _19578_);
  nor (_19587_, _19586_, _04500_);
  nor (_19589_, _04499_, _19576_);
  or (_19590_, _19589_, _19587_);
  and (_19591_, _19590_, _04515_);
  nor (_19592_, _12625_, _09161_);
  nor (_19593_, _19592_, _19578_);
  nor (_19594_, _19593_, _04515_);
  or (_19595_, _19594_, _19591_);
  and (_19596_, _19595_, _03516_);
  nor (_19597_, _05989_, _19576_);
  and (_19598_, _12638_, _05989_);
  nor (_19600_, _19598_, _19597_);
  nor (_19601_, _19600_, _03516_);
  or (_19602_, _19601_, _03597_);
  or (_19603_, _19602_, _19596_);
  nand (_19604_, _19583_, _03597_);
  and (_19605_, _19604_, _19603_);
  and (_19606_, _19605_, _03611_);
  nor (_19607_, _19586_, _03611_);
  or (_19608_, _19607_, _19606_);
  and (_19609_, _19608_, _03512_);
  and (_19611_, _12622_, _05989_);
  nor (_19612_, _19611_, _19597_);
  nor (_19613_, _19612_, _03512_);
  or (_19614_, _19613_, _19609_);
  and (_19615_, _19614_, _03505_);
  nor (_19616_, _19597_, _12653_);
  nor (_19617_, _19616_, _19600_);
  and (_19618_, _19617_, _03504_);
  or (_19619_, _19618_, _19615_);
  and (_19620_, _19619_, _03501_);
  nor (_19622_, _12671_, _09198_);
  nor (_19623_, _19622_, _19597_);
  nor (_19624_, _19623_, _03501_);
  nor (_19625_, _19624_, _07441_);
  not (_19626_, _19625_);
  nor (_19627_, _19626_, _19620_);
  nor (_19628_, _19627_, _19584_);
  nor (_19629_, _19628_, _05969_);
  and (_19630_, _06838_, _05376_);
  nor (_19631_, _19578_, _05970_);
  not (_19633_, _19631_);
  nor (_19634_, _19633_, _19630_);
  or (_19635_, _19634_, _03644_);
  nor (_19636_, _19635_, _19629_);
  nor (_19637_, _12731_, _09161_);
  nor (_19638_, _19578_, _19637_);
  nor (_19639_, _19638_, _03275_);
  or (_19640_, _19639_, _03650_);
  nor (_19641_, _19640_, _19636_);
  nor (_19642_, _19641_, _19581_);
  or (_19644_, _19642_, _03649_);
  and (_19645_, _12746_, _05376_);
  or (_19646_, _19645_, _19578_);
  or (_19647_, _19646_, _04591_);
  and (_19648_, _19647_, _04589_);
  and (_19649_, _19648_, _19644_);
  and (_19650_, _12619_, _05376_);
  nor (_19651_, _19650_, _19578_);
  nor (_19652_, _19651_, _04589_);
  nor (_19653_, _19652_, _19649_);
  nor (_19655_, _19653_, _03655_);
  nor (_19656_, _19578_, _05650_);
  not (_19657_, _19656_);
  nor (_19658_, _19580_, _04596_);
  and (_19659_, _19658_, _19657_);
  nor (_19660_, _19659_, _19655_);
  nor (_19661_, _19660_, _03773_);
  nor (_19662_, _19586_, _04594_);
  and (_19663_, _19662_, _19657_);
  nor (_19664_, _19663_, _03653_);
  not (_19666_, _19664_);
  nor (_19667_, _19666_, _19661_);
  nor (_19668_, _12745_, _09161_);
  or (_19669_, _19578_, _04608_);
  nor (_19670_, _19669_, _19668_);
  or (_19671_, _19670_, _03786_);
  nor (_19672_, _19671_, _19667_);
  nor (_19673_, _12618_, _09161_);
  nor (_19674_, _19673_, _19578_);
  nor (_19675_, _19674_, _04606_);
  or (_19677_, _19675_, _19672_);
  and (_19678_, _19677_, _04260_);
  nor (_19679_, _19593_, _04260_);
  or (_19680_, _19679_, _19678_);
  and (_19681_, _19680_, _03206_);
  nor (_19682_, _19612_, _03206_);
  or (_19683_, _19682_, _19681_);
  and (_19684_, _19683_, _03820_);
  and (_19685_, _12806_, _05376_);
  nor (_19686_, _19685_, _19578_);
  nor (_19688_, _19686_, _03820_);
  or (_19689_, _19688_, _19684_);
  or (_19690_, _19689_, _43231_);
  or (_19691_, _43227_, \oc8051_golden_model_1.IP [3]);
  and (_19692_, _19691_, _41991_);
  and (_43472_, _19692_, _19690_);
  not (_19693_, \oc8051_golden_model_1.IP [4]);
  nor (_19694_, _05376_, _19693_);
  nor (_19695_, _05840_, _09161_);
  nor (_19696_, _19695_, _19694_);
  and (_19698_, _19696_, _07441_);
  nor (_19699_, _05989_, _19693_);
  and (_19700_, _12853_, _05989_);
  nor (_19701_, _19700_, _19699_);
  nor (_19702_, _19701_, _03512_);
  and (_19703_, _05376_, \oc8051_golden_model_1.ACC [4]);
  nor (_19704_, _19703_, _19694_);
  nor (_19705_, _19704_, _04500_);
  nor (_19706_, _04499_, _19693_);
  or (_19707_, _19706_, _19705_);
  and (_19709_, _19707_, _04515_);
  nor (_19710_, _12820_, _09161_);
  nor (_19711_, _19710_, _19694_);
  nor (_19712_, _19711_, _04515_);
  or (_19713_, _19712_, _19709_);
  and (_19714_, _19713_, _03516_);
  and (_19715_, _12830_, _05989_);
  nor (_19716_, _19715_, _19699_);
  nor (_19717_, _19716_, _03516_);
  or (_19718_, _19717_, _03597_);
  or (_19720_, _19718_, _19714_);
  nand (_19721_, _19696_, _03597_);
  and (_19722_, _19721_, _19720_);
  and (_19723_, _19722_, _03611_);
  nor (_19724_, _19704_, _03611_);
  or (_19725_, _19724_, _19723_);
  and (_19726_, _19725_, _03512_);
  nor (_19727_, _19726_, _19702_);
  nor (_19728_, _19727_, _03504_);
  nor (_19729_, _19699_, _12860_);
  or (_19731_, _19716_, _03505_);
  nor (_19732_, _19731_, _19729_);
  nor (_19733_, _19732_, _19728_);
  nor (_19734_, _19733_, _03500_);
  nor (_19735_, _12828_, _09198_);
  nor (_19736_, _19735_, _19699_);
  nor (_19737_, _19736_, _03501_);
  nor (_19738_, _19737_, _07441_);
  not (_19739_, _19738_);
  nor (_19740_, _19739_, _19734_);
  nor (_19742_, _19740_, _19698_);
  nor (_19743_, _19742_, _05969_);
  and (_19744_, _06843_, _05376_);
  nor (_19745_, _19694_, _05970_);
  not (_19746_, _19745_);
  nor (_19747_, _19746_, _19744_);
  nor (_19748_, _19747_, _03644_);
  not (_19749_, _19748_);
  nor (_19750_, _19749_, _19743_);
  nor (_19751_, _12936_, _09161_);
  nor (_19753_, _19751_, _19694_);
  nor (_19754_, _19753_, _03275_);
  or (_19755_, _19754_, _08861_);
  or (_19756_, _19755_, _19750_);
  and (_19757_, _12951_, _05376_);
  or (_19758_, _19694_, _04591_);
  or (_19759_, _19758_, _19757_);
  and (_19760_, _06375_, _05376_);
  nor (_19761_, _19760_, _19694_);
  and (_19762_, _19761_, _03650_);
  nor (_19764_, _19762_, _03778_);
  and (_19765_, _19764_, _19759_);
  and (_19766_, _19765_, _19756_);
  and (_19767_, _12957_, _05376_);
  nor (_19768_, _19767_, _19694_);
  nor (_19769_, _19768_, _04589_);
  nor (_19770_, _19769_, _19766_);
  nor (_19771_, _19770_, _03655_);
  nor (_19772_, _19694_, _05889_);
  not (_19773_, _19772_);
  nor (_19775_, _19761_, _04596_);
  and (_19776_, _19775_, _19773_);
  nor (_19777_, _19776_, _19771_);
  nor (_19778_, _19777_, _03773_);
  nor (_19779_, _19704_, _04594_);
  and (_19780_, _19779_, _19773_);
  or (_19781_, _19780_, _19778_);
  and (_19782_, _19781_, _04608_);
  nor (_19783_, _12949_, _09161_);
  nor (_19784_, _19783_, _19694_);
  nor (_19786_, _19784_, _04608_);
  or (_19787_, _19786_, _19782_);
  and (_19788_, _19787_, _04606_);
  nor (_19789_, _12956_, _09161_);
  nor (_19790_, _19789_, _19694_);
  nor (_19791_, _19790_, _04606_);
  or (_19792_, _19791_, _19788_);
  and (_19793_, _19792_, _04260_);
  nor (_19794_, _19711_, _04260_);
  or (_19795_, _19794_, _19793_);
  and (_19797_, _19795_, _03206_);
  nor (_19798_, _19701_, _03206_);
  or (_19799_, _19798_, _19797_);
  and (_19800_, _19799_, _03820_);
  and (_19801_, _13013_, _05376_);
  nor (_19802_, _19801_, _19694_);
  nor (_19803_, _19802_, _03820_);
  or (_19804_, _19803_, _19800_);
  or (_19805_, _19804_, _43231_);
  or (_19806_, _43227_, \oc8051_golden_model_1.IP [4]);
  and (_19808_, _19806_, _41991_);
  and (_43473_, _19808_, _19805_);
  not (_19809_, \oc8051_golden_model_1.IP [5]);
  nor (_19810_, _05376_, _19809_);
  and (_19811_, _06842_, _05376_);
  or (_19812_, _19811_, _19810_);
  and (_19813_, _19812_, _05969_);
  and (_19814_, _05376_, \oc8051_golden_model_1.ACC [5]);
  nor (_19815_, _19814_, _19810_);
  nor (_19816_, _19815_, _04500_);
  nor (_19818_, _04499_, _19809_);
  or (_19819_, _19818_, _19816_);
  and (_19820_, _19819_, _04515_);
  nor (_19821_, _13035_, _09161_);
  nor (_19822_, _19821_, _19810_);
  nor (_19823_, _19822_, _04515_);
  or (_19824_, _19823_, _19820_);
  and (_19825_, _19824_, _03516_);
  nor (_19826_, _05989_, _19809_);
  and (_19827_, _13051_, _05989_);
  nor (_19829_, _19827_, _19826_);
  nor (_19830_, _19829_, _03516_);
  or (_19831_, _19830_, _03597_);
  or (_19832_, _19831_, _19825_);
  nor (_19833_, _05552_, _09161_);
  nor (_19834_, _19833_, _19810_);
  nand (_19835_, _19834_, _03597_);
  and (_19836_, _19835_, _19832_);
  and (_19837_, _19836_, _03611_);
  nor (_19838_, _19815_, _03611_);
  or (_19840_, _19838_, _19837_);
  and (_19841_, _19840_, _03512_);
  and (_19842_, _13032_, _05989_);
  nor (_19843_, _19842_, _19826_);
  nor (_19844_, _19843_, _03512_);
  or (_19845_, _19844_, _19841_);
  and (_19846_, _19845_, _03505_);
  nor (_19847_, _19826_, _13066_);
  nor (_19848_, _19847_, _19829_);
  and (_19849_, _19848_, _03504_);
  or (_19851_, _19849_, _19846_);
  and (_19852_, _19851_, _03501_);
  nor (_19853_, _13030_, _09198_);
  nor (_19854_, _19853_, _19826_);
  nor (_19855_, _19854_, _03501_);
  nor (_19856_, _19855_, _07441_);
  not (_19857_, _19856_);
  nor (_19858_, _19857_, _19852_);
  and (_19859_, _19834_, _07441_);
  or (_19860_, _19859_, _05969_);
  nor (_19862_, _19860_, _19858_);
  or (_19863_, _19862_, _19813_);
  and (_19864_, _19863_, _03275_);
  nor (_19865_, _13139_, _09161_);
  nor (_19866_, _19865_, _19810_);
  nor (_19867_, _19866_, _03275_);
  or (_19868_, _19867_, _08861_);
  or (_19869_, _19868_, _19864_);
  and (_19870_, _13154_, _05376_);
  or (_19871_, _19810_, _04591_);
  or (_19873_, _19871_, _19870_);
  and (_19874_, _06358_, _05376_);
  nor (_19875_, _19874_, _19810_);
  and (_19876_, _19875_, _03650_);
  nor (_19877_, _19876_, _03778_);
  and (_19878_, _19877_, _19873_);
  and (_19879_, _19878_, _19869_);
  and (_19880_, _13160_, _05376_);
  nor (_19881_, _19880_, _19810_);
  nor (_19882_, _19881_, _04589_);
  nor (_19884_, _19882_, _19879_);
  nor (_19885_, _19884_, _03655_);
  nor (_19886_, _19810_, _05601_);
  not (_19887_, _19886_);
  nor (_19888_, _19875_, _04596_);
  and (_19889_, _19888_, _19887_);
  nor (_19890_, _19889_, _19885_);
  nor (_19891_, _19890_, _03773_);
  nor (_19892_, _19815_, _04594_);
  and (_19893_, _19892_, _19887_);
  or (_19895_, _19893_, _19891_);
  and (_19896_, _19895_, _04608_);
  nor (_19897_, _13152_, _09161_);
  nor (_19898_, _19897_, _19810_);
  nor (_19899_, _19898_, _04608_);
  or (_19900_, _19899_, _19896_);
  and (_19901_, _19900_, _04606_);
  nor (_19902_, _13159_, _09161_);
  nor (_19903_, _19902_, _19810_);
  nor (_19904_, _19903_, _04606_);
  or (_19906_, _19904_, _19901_);
  and (_19907_, _19906_, _04260_);
  nor (_19908_, _19822_, _04260_);
  or (_19909_, _19908_, _19907_);
  and (_19910_, _19909_, _03206_);
  nor (_19911_, _19843_, _03206_);
  or (_19912_, _19911_, _19910_);
  and (_19913_, _19912_, _03820_);
  and (_19914_, _13217_, _05376_);
  nor (_19915_, _19914_, _19810_);
  nor (_19917_, _19915_, _03820_);
  or (_19918_, _19917_, _19913_);
  or (_19919_, _19918_, _43231_);
  or (_19920_, _43227_, \oc8051_golden_model_1.IP [5]);
  and (_19921_, _19920_, _41991_);
  and (_43474_, _19921_, _19919_);
  not (_19922_, \oc8051_golden_model_1.IP [6]);
  nor (_19923_, _05376_, _19922_);
  and (_19924_, _06531_, _05376_);
  or (_19925_, _19924_, _19923_);
  and (_19927_, _19925_, _05969_);
  and (_19928_, _05376_, \oc8051_golden_model_1.ACC [6]);
  nor (_19929_, _19928_, _19923_);
  nor (_19930_, _19929_, _04500_);
  nor (_19931_, _04499_, _19922_);
  or (_19932_, _19931_, _19930_);
  and (_19933_, _19932_, _04515_);
  nor (_19934_, _13235_, _09161_);
  nor (_19935_, _19934_, _19923_);
  nor (_19936_, _19935_, _04515_);
  or (_19938_, _19936_, _19933_);
  and (_19939_, _19938_, _03516_);
  nor (_19940_, _05989_, _19922_);
  and (_19941_, _13266_, _05989_);
  nor (_19942_, _19941_, _19940_);
  nor (_19943_, _19942_, _03516_);
  or (_19944_, _19943_, _03597_);
  or (_19945_, _19944_, _19939_);
  nor (_19946_, _05442_, _09161_);
  nor (_19947_, _19946_, _19923_);
  nand (_19949_, _19947_, _03597_);
  and (_19950_, _19949_, _19945_);
  and (_19951_, _19950_, _03611_);
  nor (_19952_, _19929_, _03611_);
  or (_19953_, _19952_, _19951_);
  and (_19954_, _19953_, _03512_);
  and (_19955_, _13251_, _05989_);
  nor (_19956_, _19955_, _19940_);
  nor (_19957_, _19956_, _03512_);
  or (_19958_, _19957_, _03504_);
  or (_19960_, _19958_, _19954_);
  nor (_19961_, _19940_, _13281_);
  nor (_19962_, _19961_, _19942_);
  or (_19963_, _19962_, _03505_);
  and (_19964_, _19963_, _03501_);
  and (_19965_, _19964_, _19960_);
  nor (_19966_, _13249_, _09198_);
  nor (_19967_, _19966_, _19940_);
  nor (_19968_, _19967_, _03501_);
  nor (_19969_, _19968_, _07441_);
  not (_19971_, _19969_);
  nor (_19972_, _19971_, _19965_);
  and (_19973_, _19947_, _07441_);
  or (_19974_, _19973_, _05969_);
  nor (_19975_, _19974_, _19972_);
  or (_19976_, _19975_, _19927_);
  and (_19977_, _19976_, _03275_);
  nor (_19978_, _13356_, _09161_);
  nor (_19979_, _19978_, _19923_);
  nor (_19980_, _19979_, _03275_);
  or (_19982_, _19980_, _08861_);
  or (_19983_, _19982_, _19977_);
  and (_19984_, _13245_, _05376_);
  or (_19985_, _19923_, _04591_);
  or (_19986_, _19985_, _19984_);
  and (_19987_, _13363_, _05376_);
  nor (_19988_, _19987_, _19923_);
  and (_19989_, _19988_, _03650_);
  nor (_19990_, _19989_, _03778_);
  and (_19991_, _19990_, _19986_);
  and (_19993_, _19991_, _19983_);
  and (_19994_, _13374_, _05376_);
  nor (_19995_, _19994_, _19923_);
  nor (_19996_, _19995_, _04589_);
  nor (_19997_, _19996_, _19993_);
  nor (_19998_, _19997_, _03655_);
  nor (_19999_, _19923_, _05491_);
  not (_20000_, _19999_);
  nor (_20001_, _19988_, _04596_);
  and (_20002_, _20001_, _20000_);
  nor (_20004_, _20002_, _19998_);
  nor (_20005_, _20004_, _03773_);
  nor (_20006_, _19929_, _04594_);
  and (_20007_, _20006_, _20000_);
  or (_20008_, _20007_, _20005_);
  and (_20009_, _20008_, _04608_);
  nor (_20010_, _13243_, _09161_);
  nor (_20011_, _20010_, _19923_);
  nor (_20012_, _20011_, _04608_);
  or (_20013_, _20012_, _20009_);
  and (_20015_, _20013_, _04606_);
  nor (_20016_, _13373_, _09161_);
  nor (_20017_, _20016_, _19923_);
  nor (_20018_, _20017_, _04606_);
  or (_20019_, _20018_, _20015_);
  and (_20020_, _20019_, _04260_);
  nor (_20021_, _19935_, _04260_);
  or (_20022_, _20021_, _20020_);
  and (_20023_, _20022_, _03206_);
  nor (_20024_, _19956_, _03206_);
  or (_20026_, _20024_, _20023_);
  and (_20027_, _20026_, _03820_);
  and (_20028_, _13425_, _05376_);
  nor (_20029_, _20028_, _19923_);
  nor (_20030_, _20029_, _03820_);
  or (_20031_, _20030_, _20027_);
  or (_20032_, _20031_, _43231_);
  or (_20033_, _43227_, \oc8051_golden_model_1.IP [6]);
  and (_20034_, _20033_, _41991_);
  and (_43475_, _20034_, _20032_);
  not (_20036_, \oc8051_golden_model_1.P0 [0]);
  nor (_20037_, _43227_, _20036_);
  or (_20038_, _20037_, rst);
  nor (_20039_, _05363_, _20036_);
  and (_20040_, _12145_, _05363_);
  or (_20041_, _20040_, _20039_);
  and (_20042_, _20041_, _03778_);
  and (_20043_, _05363_, _04491_);
  or (_20044_, _20043_, _20039_);
  or (_20045_, _20044_, _06889_);
  nor (_20047_, _05744_, _09268_);
  or (_20048_, _20047_, _20039_);
  and (_20049_, _20048_, _03599_);
  nor (_20050_, _04499_, _20036_);
  and (_20051_, _05363_, \oc8051_golden_model_1.ACC [0]);
  or (_20052_, _20051_, _20039_);
  and (_20053_, _20052_, _04499_);
  or (_20054_, _20053_, _20050_);
  and (_20055_, _20054_, _04515_);
  or (_20056_, _20055_, _03515_);
  or (_20058_, _20056_, _20049_);
  and (_20059_, _12035_, _05294_);
  nor (_20060_, _05294_, _20036_);
  or (_20061_, _20060_, _03516_);
  or (_20062_, _20061_, _20059_);
  and (_20063_, _20062_, _04524_);
  and (_20064_, _20063_, _20058_);
  and (_20065_, _20044_, _03597_);
  or (_20066_, _20065_, _03603_);
  or (_20067_, _20066_, _20064_);
  or (_20069_, _20052_, _03611_);
  and (_20070_, _20069_, _03512_);
  and (_20071_, _20070_, _20067_);
  and (_20072_, _20039_, _03511_);
  or (_20073_, _20072_, _03504_);
  or (_20074_, _20073_, _20071_);
  or (_20075_, _20048_, _03505_);
  and (_20076_, _20075_, _03501_);
  and (_20077_, _20076_, _20074_);
  or (_20078_, _12065_, _12023_);
  and (_20080_, _20078_, _05294_);
  or (_20081_, _20080_, _20060_);
  and (_20082_, _20081_, _03500_);
  or (_20083_, _20082_, _07441_);
  or (_20084_, _20083_, _20077_);
  and (_20085_, _20084_, _20045_);
  or (_20086_, _20085_, _05969_);
  and (_20087_, _06836_, _05363_);
  or (_20088_, _20039_, _05970_);
  or (_20089_, _20088_, _20087_);
  and (_20091_, _20089_, _03275_);
  and (_20092_, _20091_, _20086_);
  and (_20093_, _06378_, \oc8051_golden_model_1.P1 [0]);
  and (_20094_, _06356_, \oc8051_golden_model_1.P0 [0]);
  and (_20095_, _06361_, \oc8051_golden_model_1.P2 [0]);
  nor (_20096_, _20095_, _20094_);
  nand (_20097_, _20096_, _12090_);
  or (_20098_, _20097_, _20093_);
  not (_20099_, _12121_);
  and (_20100_, _12112_, _20099_);
  nand (_20102_, _20100_, _12103_);
  not (_20103_, _12119_);
  nand (_20104_, _20103_, _12115_);
  or (_20105_, _12091_, _12093_);
  and (_20106_, _06382_, \oc8051_golden_model_1.P3 [0]);
  or (_20107_, _20106_, _12117_);
  or (_20108_, _20107_, _20105_);
  or (_20109_, _20108_, _12122_);
  or (_20110_, _20109_, _20104_);
  or (_20111_, _20110_, _20102_);
  or (_20113_, _20111_, _20098_);
  or (_20114_, _20113_, _12078_);
  and (_20115_, _20114_, _05363_);
  or (_20116_, _20115_, _20039_);
  and (_20117_, _20116_, _03644_);
  or (_20118_, _20117_, _20092_);
  or (_20119_, _20118_, _08861_);
  and (_20120_, _12019_, _05363_);
  or (_20121_, _20039_, _04591_);
  or (_20122_, _20121_, _20120_);
  and (_20124_, _05363_, _06366_);
  or (_20125_, _20124_, _20039_);
  or (_20126_, _20125_, _04582_);
  and (_20127_, _20126_, _04589_);
  and (_20128_, _20127_, _20122_);
  and (_20129_, _20128_, _20119_);
  or (_20130_, _20129_, _20042_);
  and (_20131_, _20130_, _04596_);
  nand (_20132_, _20125_, _03655_);
  nor (_20133_, _20132_, _20047_);
  or (_20135_, _20133_, _20131_);
  and (_20136_, _20135_, _04594_);
  or (_20137_, _20039_, _05744_);
  and (_20138_, _20052_, _03773_);
  and (_20139_, _20138_, _20137_);
  or (_20140_, _20139_, _03653_);
  or (_20141_, _20140_, _20136_);
  nor (_20142_, _12017_, _09268_);
  or (_20143_, _20039_, _04608_);
  or (_20144_, _20143_, _20142_);
  and (_20146_, _20144_, _04606_);
  and (_20147_, _20146_, _20141_);
  nor (_20148_, _12015_, _09268_);
  or (_20149_, _20148_, _20039_);
  and (_20150_, _20149_, _03786_);
  or (_20151_, _20150_, _03809_);
  or (_20152_, _20151_, _20147_);
  or (_20153_, _20048_, _04260_);
  and (_20154_, _20153_, _03206_);
  and (_20155_, _20154_, _20152_);
  and (_20157_, _20039_, _03205_);
  or (_20158_, _20157_, _03816_);
  or (_20159_, _20158_, _20155_);
  or (_20160_, _20048_, _03820_);
  and (_20161_, _20160_, _43227_);
  and (_20162_, _20161_, _20159_);
  or (_43476_, _20162_, _20038_);
  not (_20163_, \oc8051_golden_model_1.P0 [1]);
  nor (_20164_, _05363_, _20163_);
  and (_20165_, _05363_, _05898_);
  or (_20167_, _20165_, _20164_);
  or (_20168_, _20167_, _04524_);
  or (_20169_, _05363_, \oc8051_golden_model_1.P0 [1]);
  and (_20170_, _12234_, _05363_);
  not (_20171_, _20170_);
  and (_20172_, _20171_, _20169_);
  or (_20173_, _20172_, _04515_);
  nand (_20174_, _05363_, _03320_);
  and (_20175_, _20174_, _20169_);
  and (_20176_, _20175_, _04499_);
  nor (_20178_, _04499_, _20163_);
  or (_20179_, _20178_, _03599_);
  or (_20180_, _20179_, _20176_);
  and (_20181_, _20180_, _03516_);
  and (_20182_, _20181_, _20173_);
  nor (_20183_, _05294_, _20163_);
  and (_20184_, _12238_, _05294_);
  or (_20185_, _20184_, _20183_);
  and (_20186_, _20185_, _03515_);
  or (_20187_, _20186_, _03597_);
  or (_20189_, _20187_, _20182_);
  and (_20190_, _20189_, _20168_);
  or (_20191_, _20190_, _03603_);
  or (_20192_, _20175_, _03611_);
  and (_20193_, _20192_, _03512_);
  and (_20194_, _20193_, _20191_);
  and (_20195_, _12224_, _05294_);
  or (_20196_, _20195_, _20183_);
  and (_20197_, _20196_, _03511_);
  or (_20198_, _20197_, _03504_);
  or (_20200_, _20198_, _20194_);
  and (_20201_, _20184_, _12253_);
  or (_20202_, _20183_, _03505_);
  or (_20203_, _20202_, _20201_);
  and (_20204_, _20203_, _20200_);
  and (_20205_, _20204_, _03501_);
  or (_20206_, _12269_, _12224_);
  and (_20207_, _20206_, _05294_);
  or (_20208_, _20183_, _20207_);
  and (_20209_, _20208_, _03500_);
  or (_20211_, _20209_, _07441_);
  or (_20212_, _20211_, _20205_);
  or (_20213_, _20167_, _06889_);
  and (_20214_, _20213_, _20212_);
  or (_20215_, _20214_, _05969_);
  and (_20216_, _06835_, _05363_);
  or (_20217_, _20164_, _05970_);
  or (_20218_, _20217_, _20216_);
  and (_20219_, _20218_, _03275_);
  and (_20220_, _20219_, _20215_);
  and (_20222_, _06361_, \oc8051_golden_model_1.P2 [1]);
  and (_20223_, _06356_, \oc8051_golden_model_1.P0 [1]);
  or (_20224_, _20223_, _12283_);
  or (_20225_, _20224_, _20222_);
  and (_20226_, _06378_, \oc8051_golden_model_1.P1 [1]);
  and (_20227_, _06382_, \oc8051_golden_model_1.P3 [1]);
  or (_20228_, _20227_, _20226_);
  or (_20229_, _20228_, _12291_);
  or (_20230_, _20229_, _12289_);
  nor (_20231_, _20230_, _20225_);
  and (_20233_, _20231_, _12308_);
  nand (_20234_, _20233_, _12327_);
  or (_20235_, _20234_, _12282_);
  and (_20236_, _20235_, _05363_);
  or (_20237_, _20236_, _20164_);
  and (_20238_, _20237_, _03644_);
  or (_20239_, _20238_, _20220_);
  and (_20240_, _20239_, _03651_);
  or (_20241_, _12220_, _09268_);
  and (_20242_, _20241_, _03649_);
  nand (_20244_, _05363_, _04347_);
  and (_20245_, _20244_, _03650_);
  or (_20246_, _20245_, _20242_);
  and (_20247_, _20246_, _20169_);
  or (_20248_, _20247_, _20240_);
  and (_20249_, _20248_, _04589_);
  or (_20250_, _12347_, _09268_);
  and (_20251_, _20169_, _03778_);
  and (_20252_, _20251_, _20250_);
  or (_20253_, _20252_, _20249_);
  and (_20255_, _20253_, _04596_);
  or (_20256_, _12219_, _09268_);
  and (_20257_, _20169_, _03655_);
  and (_20258_, _20257_, _20256_);
  or (_20259_, _20258_, _20255_);
  and (_20260_, _20259_, _04594_);
  or (_20261_, _20164_, _05699_);
  and (_20262_, _20175_, _03773_);
  and (_20263_, _20262_, _20261_);
  or (_20264_, _20263_, _20260_);
  and (_20266_, _20264_, _03787_);
  or (_20267_, _20244_, _05699_);
  and (_20268_, _20169_, _03653_);
  and (_20269_, _20268_, _20267_);
  or (_20270_, _20174_, _05699_);
  and (_20271_, _20169_, _03786_);
  and (_20272_, _20271_, _20270_);
  or (_20273_, _20272_, _03809_);
  or (_20274_, _20273_, _20269_);
  or (_20275_, _20274_, _20266_);
  or (_20277_, _20172_, _04260_);
  and (_20278_, _20277_, _03206_);
  and (_20279_, _20278_, _20275_);
  and (_20280_, _20196_, _03205_);
  or (_20281_, _20280_, _03816_);
  or (_20282_, _20281_, _20279_);
  or (_20283_, _20164_, _03820_);
  or (_20284_, _20283_, _20170_);
  and (_20285_, _20284_, _43227_);
  and (_20286_, _20285_, _20282_);
  nor (_20288_, _43227_, _20163_);
  or (_20289_, _20288_, rst);
  or (_43477_, _20289_, _20286_);
  not (_20290_, \oc8051_golden_model_1.P0 [2]);
  nor (_20291_, _05363_, _20290_);
  nor (_20292_, _09268_, _05130_);
  or (_20293_, _20292_, _20291_);
  or (_20294_, _20293_, _06889_);
  or (_20295_, _20293_, _04524_);
  nor (_20296_, _12430_, _09268_);
  or (_20298_, _20296_, _20291_);
  or (_20299_, _20298_, _04515_);
  and (_20300_, _05363_, \oc8051_golden_model_1.ACC [2]);
  or (_20301_, _20300_, _20291_);
  and (_20302_, _20301_, _04499_);
  nor (_20303_, _04499_, _20290_);
  or (_20304_, _20303_, _03599_);
  or (_20305_, _20304_, _20302_);
  and (_20306_, _20305_, _03516_);
  and (_20307_, _20306_, _20299_);
  nor (_20309_, _05294_, _20290_);
  and (_20310_, _12416_, _05294_);
  or (_20311_, _20310_, _20309_);
  and (_20312_, _20311_, _03515_);
  or (_20313_, _20312_, _03597_);
  or (_20314_, _20313_, _20307_);
  and (_20315_, _20314_, _20295_);
  or (_20316_, _20315_, _03603_);
  or (_20317_, _20301_, _03611_);
  and (_20318_, _20317_, _03512_);
  and (_20320_, _20318_, _20316_);
  and (_20321_, _12414_, _05294_);
  or (_20322_, _20321_, _20309_);
  and (_20323_, _20322_, _03511_);
  or (_20324_, _20323_, _03504_);
  or (_20325_, _20324_, _20320_);
  and (_20326_, _20310_, _12447_);
  or (_20327_, _20309_, _03505_);
  or (_20328_, _20327_, _20326_);
  and (_20329_, _20328_, _03501_);
  and (_20331_, _20329_, _20325_);
  or (_20332_, _12464_, _12414_);
  and (_20333_, _20332_, _05294_);
  or (_20334_, _20333_, _20309_);
  and (_20335_, _20334_, _03500_);
  or (_20336_, _20335_, _07441_);
  or (_20337_, _20336_, _20331_);
  and (_20338_, _20337_, _20294_);
  or (_20339_, _20338_, _05969_);
  and (_20340_, _06839_, _05363_);
  or (_20342_, _20291_, _05970_);
  or (_20343_, _20342_, _20340_);
  and (_20344_, _20343_, _03275_);
  and (_20345_, _20344_, _20339_);
  and (_20346_, _06378_, \oc8051_golden_model_1.P1 [2]);
  and (_20347_, _06382_, \oc8051_golden_model_1.P3 [2]);
  or (_20348_, _20347_, _20346_);
  or (_20349_, _20348_, _12481_);
  and (_20350_, _06356_, \oc8051_golden_model_1.P0 [2]);
  and (_20351_, _06361_, \oc8051_golden_model_1.P2 [2]);
  or (_20353_, _20351_, _20350_);
  or (_20354_, _20353_, _20349_);
  nor (_20355_, _20354_, _12479_);
  and (_20356_, _20355_, _12505_);
  nand (_20357_, _20356_, _12521_);
  or (_20358_, _20357_, _12478_);
  and (_20359_, _20358_, _05363_);
  or (_20360_, _20291_, _20359_);
  and (_20361_, _20360_, _03644_);
  or (_20362_, _20361_, _20345_);
  or (_20364_, _20362_, _08861_);
  and (_20365_, _12538_, _05363_);
  or (_20366_, _20291_, _04591_);
  or (_20367_, _20366_, _20365_);
  and (_20368_, _05363_, _06414_);
  or (_20369_, _20368_, _20291_);
  or (_20370_, _20369_, _04582_);
  and (_20371_, _20370_, _04589_);
  and (_20372_, _20371_, _20367_);
  and (_20373_, _20372_, _20364_);
  and (_20375_, _12544_, _05363_);
  or (_20376_, _20375_, _20291_);
  and (_20377_, _20376_, _03778_);
  or (_20378_, _20377_, _20373_);
  and (_20379_, _20378_, _04596_);
  or (_20380_, _20291_, _05793_);
  and (_20381_, _20369_, _03655_);
  and (_20382_, _20381_, _20380_);
  or (_20383_, _20382_, _20379_);
  and (_20384_, _20383_, _04594_);
  and (_20386_, _20301_, _03773_);
  and (_20387_, _20386_, _20380_);
  or (_20388_, _20387_, _03653_);
  or (_20389_, _20388_, _20384_);
  nor (_20390_, _12537_, _09268_);
  or (_20391_, _20291_, _04608_);
  or (_20392_, _20391_, _20390_);
  and (_20393_, _20392_, _04606_);
  and (_20394_, _20393_, _20389_);
  nor (_20395_, _12543_, _09268_);
  or (_20397_, _20395_, _20291_);
  and (_20398_, _20397_, _03786_);
  or (_20399_, _20398_, _03809_);
  or (_20400_, _20399_, _20394_);
  or (_20401_, _20298_, _04260_);
  and (_20402_, _20401_, _03206_);
  and (_20403_, _20402_, _20400_);
  and (_20404_, _20322_, _03205_);
  or (_20405_, _20404_, _03816_);
  or (_20406_, _20405_, _20403_);
  and (_20408_, _12600_, _05363_);
  or (_20409_, _20291_, _03820_);
  or (_20410_, _20409_, _20408_);
  and (_20411_, _20410_, _43227_);
  and (_20412_, _20411_, _20406_);
  nor (_20413_, _43227_, _20290_);
  or (_20414_, _20413_, rst);
  or (_43478_, _20414_, _20412_);
  not (_20415_, \oc8051_golden_model_1.P0 [3]);
  nor (_20416_, _43227_, _20415_);
  or (_20418_, _20416_, rst);
  nor (_20419_, _05363_, _20415_);
  nor (_20420_, _09268_, _04944_);
  or (_20421_, _20420_, _20419_);
  or (_20422_, _20421_, _06889_);
  nor (_20423_, _12625_, _09268_);
  or (_20424_, _20423_, _20419_);
  or (_20425_, _20424_, _04515_);
  and (_20426_, _05363_, \oc8051_golden_model_1.ACC [3]);
  or (_20427_, _20426_, _20419_);
  and (_20429_, _20427_, _04499_);
  nor (_20430_, _04499_, _20415_);
  or (_20431_, _20430_, _03599_);
  or (_20432_, _20431_, _20429_);
  and (_20433_, _20432_, _03516_);
  and (_20434_, _20433_, _20425_);
  nor (_20435_, _05294_, _20415_);
  and (_20436_, _12638_, _05294_);
  or (_20437_, _20436_, _20435_);
  and (_20438_, _20437_, _03515_);
  or (_20440_, _20438_, _03597_);
  or (_20441_, _20440_, _20434_);
  or (_20442_, _20421_, _04524_);
  and (_20443_, _20442_, _20441_);
  or (_20444_, _20443_, _03603_);
  or (_20445_, _20427_, _03611_);
  and (_20446_, _20445_, _03512_);
  and (_20447_, _20446_, _20444_);
  and (_20448_, _12622_, _05294_);
  or (_20449_, _20448_, _20435_);
  and (_20450_, _20449_, _03511_);
  or (_20451_, _20450_, _03504_);
  or (_20452_, _20451_, _20447_);
  or (_20453_, _20435_, _12653_);
  and (_20454_, _20453_, _20437_);
  or (_20455_, _20454_, _03505_);
  and (_20456_, _20455_, _03501_);
  and (_20457_, _20456_, _20452_);
  or (_20458_, _12622_, _12669_);
  and (_20459_, _20458_, _05294_);
  or (_20461_, _20459_, _20435_);
  and (_20462_, _20461_, _03500_);
  or (_20463_, _20462_, _07441_);
  or (_20464_, _20463_, _20457_);
  and (_20465_, _20464_, _20422_);
  or (_20466_, _20465_, _05969_);
  and (_20467_, _06838_, _05363_);
  or (_20468_, _20419_, _05970_);
  or (_20469_, _20468_, _20467_);
  and (_20470_, _20469_, _03275_);
  and (_20472_, _20470_, _20466_);
  and (_20473_, _06378_, \oc8051_golden_model_1.P1 [3]);
  and (_20474_, _06382_, \oc8051_golden_model_1.P3 [3]);
  or (_20475_, _20474_, _20473_);
  or (_20476_, _20475_, _12723_);
  and (_20477_, _06356_, \oc8051_golden_model_1.P0 [3]);
  and (_20478_, _06361_, \oc8051_golden_model_1.P2 [3]);
  or (_20479_, _20478_, _20477_);
  or (_20480_, _20479_, _20476_);
  nor (_20481_, _20480_, _12715_);
  and (_20483_, _20481_, _12714_);
  nand (_20484_, _20483_, _12706_);
  or (_20485_, _20484_, _12683_);
  and (_20486_, _20485_, _05363_);
  or (_20487_, _20419_, _20486_);
  and (_20488_, _20487_, _03644_);
  or (_20489_, _20488_, _20472_);
  or (_20490_, _20489_, _08861_);
  and (_20491_, _12746_, _05363_);
  or (_20492_, _20419_, _04591_);
  or (_20493_, _20492_, _20491_);
  and (_20494_, _05363_, _06347_);
  or (_20495_, _20494_, _20419_);
  or (_20496_, _20495_, _04582_);
  and (_20497_, _20496_, _04589_);
  and (_20498_, _20497_, _20493_);
  and (_20499_, _20498_, _20490_);
  and (_20500_, _12619_, _05363_);
  or (_20501_, _20500_, _20419_);
  and (_20502_, _20501_, _03778_);
  or (_20504_, _20502_, _20499_);
  and (_20505_, _20504_, _04596_);
  or (_20506_, _20419_, _05650_);
  and (_20507_, _20495_, _03655_);
  and (_20508_, _20507_, _20506_);
  or (_20509_, _20508_, _20505_);
  and (_20510_, _20509_, _04594_);
  and (_20511_, _20427_, _03773_);
  and (_20512_, _20511_, _20506_);
  or (_20513_, _20512_, _03653_);
  or (_20515_, _20513_, _20510_);
  nor (_20516_, _12745_, _09268_);
  or (_20517_, _20419_, _04608_);
  or (_20518_, _20517_, _20516_);
  and (_20519_, _20518_, _04606_);
  and (_20520_, _20519_, _20515_);
  nor (_20521_, _12618_, _09268_);
  or (_20522_, _20521_, _20419_);
  and (_20523_, _20522_, _03786_);
  or (_20524_, _20523_, _03809_);
  or (_20525_, _20524_, _20520_);
  or (_20526_, _20424_, _04260_);
  and (_20527_, _20526_, _03206_);
  and (_20528_, _20527_, _20525_);
  and (_20529_, _20449_, _03205_);
  or (_20530_, _20529_, _03816_);
  or (_20531_, _20530_, _20528_);
  and (_20532_, _12806_, _05363_);
  or (_20533_, _20419_, _03820_);
  or (_20534_, _20533_, _20532_);
  and (_20536_, _20534_, _43227_);
  and (_20537_, _20536_, _20531_);
  or (_43479_, _20537_, _20418_);
  and (_20538_, _09268_, \oc8051_golden_model_1.P0 [4]);
  nor (_20539_, _05840_, _09268_);
  or (_20540_, _20539_, _20538_);
  or (_20541_, _20540_, _06889_);
  not (_20542_, \oc8051_golden_model_1.P0 [4]);
  nor (_20543_, _05294_, _20542_);
  and (_20544_, _12853_, _05294_);
  or (_20546_, _20544_, _20543_);
  and (_20547_, _20546_, _03511_);
  nor (_20548_, _12820_, _09268_);
  or (_20549_, _20548_, _20538_);
  or (_20550_, _20549_, _04515_);
  and (_20551_, _05363_, \oc8051_golden_model_1.ACC [4]);
  or (_20552_, _20551_, _20538_);
  and (_20553_, _20552_, _04499_);
  nor (_20554_, _04499_, _20542_);
  or (_20555_, _20554_, _03599_);
  or (_20556_, _20555_, _20553_);
  and (_20557_, _20556_, _03516_);
  and (_20558_, _20557_, _20550_);
  and (_20559_, _12830_, _05294_);
  or (_20560_, _20559_, _20543_);
  and (_20561_, _20560_, _03515_);
  or (_20562_, _20561_, _03597_);
  or (_20563_, _20562_, _20558_);
  or (_20564_, _20540_, _04524_);
  and (_20565_, _20564_, _20563_);
  or (_20567_, _20565_, _03603_);
  or (_20568_, _20552_, _03611_);
  and (_20569_, _20568_, _03512_);
  and (_20570_, _20569_, _20567_);
  or (_20571_, _20570_, _20547_);
  and (_20572_, _20571_, _03505_);
  and (_20573_, _12861_, _05294_);
  or (_20574_, _20573_, _20543_);
  and (_20575_, _20574_, _03504_);
  or (_20576_, _20575_, _20572_);
  and (_20578_, _20576_, _03501_);
  or (_20579_, _12853_, _12827_);
  and (_20580_, _20579_, _05294_);
  or (_20581_, _20580_, _20543_);
  and (_20582_, _20581_, _03500_);
  or (_20583_, _20582_, _07441_);
  or (_20584_, _20583_, _20578_);
  and (_20585_, _20584_, _20541_);
  or (_20586_, _20585_, _05969_);
  and (_20587_, _06843_, _05363_);
  or (_20588_, _20538_, _05970_);
  or (_20589_, _20588_, _20587_);
  and (_20590_, _20589_, _03275_);
  and (_20591_, _20590_, _20586_);
  and (_20592_, _06356_, \oc8051_golden_model_1.P0 [4]);
  and (_20593_, _06361_, \oc8051_golden_model_1.P2 [4]);
  or (_20594_, _20593_, _12888_);
  or (_20595_, _20594_, _20592_);
  and (_20596_, _06378_, \oc8051_golden_model_1.P1 [4]);
  and (_20597_, _06382_, \oc8051_golden_model_1.P3 [4]);
  or (_20599_, _20597_, _20596_);
  or (_20600_, _20599_, _12896_);
  or (_20601_, _20600_, _12894_);
  nor (_20602_, _20601_, _20595_);
  and (_20603_, _20602_, _12913_);
  nand (_20604_, _20603_, _12933_);
  or (_20605_, _20604_, _12887_);
  and (_20606_, _20605_, _05363_);
  or (_20607_, _20606_, _20538_);
  and (_20608_, _20607_, _03644_);
  or (_20610_, _20608_, _08861_);
  or (_20611_, _20610_, _20591_);
  and (_20612_, _12951_, _05363_);
  or (_20613_, _20538_, _04591_);
  or (_20614_, _20613_, _20612_);
  and (_20615_, _06375_, _05363_);
  or (_20616_, _20615_, _20538_);
  or (_20617_, _20616_, _04582_);
  and (_20618_, _20617_, _04589_);
  and (_20619_, _20618_, _20614_);
  and (_20620_, _20619_, _20611_);
  and (_20621_, _12957_, _05363_);
  or (_20622_, _20621_, _20538_);
  and (_20623_, _20622_, _03778_);
  or (_20624_, _20623_, _20620_);
  and (_20625_, _20624_, _04596_);
  or (_20626_, _20538_, _05889_);
  and (_20627_, _20616_, _03655_);
  and (_20628_, _20627_, _20626_);
  or (_20629_, _20628_, _20625_);
  and (_20631_, _20629_, _04594_);
  and (_20632_, _20552_, _03773_);
  and (_20633_, _20632_, _20626_);
  or (_20634_, _20633_, _03653_);
  or (_20635_, _20634_, _20631_);
  nor (_20636_, _12949_, _09268_);
  or (_20637_, _20538_, _04608_);
  or (_20638_, _20637_, _20636_);
  and (_20639_, _20638_, _04606_);
  and (_20640_, _20639_, _20635_);
  nor (_20642_, _12956_, _09268_);
  or (_20643_, _20642_, _20538_);
  and (_20644_, _20643_, _03786_);
  or (_20645_, _20644_, _03809_);
  or (_20646_, _20645_, _20640_);
  or (_20647_, _20549_, _04260_);
  and (_20648_, _20647_, _03206_);
  and (_20649_, _20648_, _20646_);
  and (_20650_, _20546_, _03205_);
  or (_20651_, _20650_, _03816_);
  or (_20652_, _20651_, _20649_);
  and (_20653_, _13013_, _05363_);
  or (_20654_, _20538_, _03820_);
  or (_20655_, _20654_, _20653_);
  and (_20656_, _20655_, _43227_);
  and (_20657_, _20656_, _20652_);
  nor (_20658_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_20659_, _20658_, _05217_);
  or (_43480_, _20659_, _20657_);
  not (_20660_, \oc8051_golden_model_1.P0 [5]);
  nor (_20662_, _43227_, _20660_);
  or (_20663_, _20662_, rst);
  nor (_20664_, _05363_, _20660_);
  nor (_20665_, _13035_, _09268_);
  or (_20666_, _20665_, _20664_);
  or (_20667_, _20666_, _04515_);
  and (_20668_, _05363_, \oc8051_golden_model_1.ACC [5]);
  or (_20669_, _20668_, _20664_);
  and (_20670_, _20669_, _04499_);
  nor (_20671_, _04499_, _20660_);
  or (_20673_, _20671_, _03599_);
  or (_20674_, _20673_, _20670_);
  and (_20675_, _20674_, _03516_);
  and (_20676_, _20675_, _20667_);
  nor (_20677_, _05294_, _20660_);
  and (_20678_, _13051_, _05294_);
  or (_20679_, _20678_, _20677_);
  and (_20680_, _20679_, _03515_);
  or (_20681_, _20680_, _03597_);
  or (_20682_, _20681_, _20676_);
  nor (_20683_, _05552_, _09268_);
  or (_20684_, _20683_, _20664_);
  or (_20685_, _20684_, _04524_);
  and (_20686_, _20685_, _20682_);
  or (_20687_, _20686_, _03603_);
  or (_20688_, _20669_, _03611_);
  and (_20689_, _20688_, _03512_);
  and (_20690_, _20689_, _20687_);
  and (_20691_, _13032_, _05294_);
  or (_20692_, _20691_, _20677_);
  and (_20694_, _20692_, _03511_);
  or (_20695_, _20694_, _03504_);
  or (_20696_, _20695_, _20690_);
  or (_20697_, _20677_, _13066_);
  and (_20698_, _20697_, _20679_);
  or (_20699_, _20698_, _03505_);
  and (_20700_, _20699_, _03501_);
  and (_20701_, _20700_, _20696_);
  or (_20702_, _13032_, _13029_);
  and (_20703_, _20702_, _05294_);
  or (_20705_, _20703_, _20677_);
  and (_20706_, _20705_, _03500_);
  or (_20707_, _20706_, _07441_);
  or (_20708_, _20707_, _20701_);
  or (_20709_, _20684_, _06889_);
  and (_20710_, _20709_, _20708_);
  or (_20711_, _20710_, _05969_);
  and (_20712_, _06842_, _05363_);
  or (_20713_, _20664_, _05970_);
  or (_20714_, _20713_, _20712_);
  and (_20715_, _20714_, _03275_);
  and (_20716_, _20715_, _20711_);
  and (_20717_, _06378_, \oc8051_golden_model_1.P1 [5]);
  and (_20718_, _06382_, \oc8051_golden_model_1.P3 [5]);
  or (_20719_, _20718_, _20717_);
  or (_20720_, _20719_, _13096_);
  and (_20721_, _06356_, \oc8051_golden_model_1.P0 [5]);
  and (_20722_, _06361_, \oc8051_golden_model_1.P2 [5]);
  or (_20723_, _20722_, _20721_);
  or (_20724_, _20723_, _20720_);
  nor (_20726_, _20724_, _13094_);
  and (_20727_, _20726_, _13120_);
  nand (_20728_, _20727_, _13136_);
  or (_20729_, _20728_, _13093_);
  and (_20730_, _20729_, _05363_);
  or (_20731_, _20730_, _20664_);
  and (_20732_, _20731_, _03644_);
  or (_20733_, _20732_, _08861_);
  or (_20734_, _20733_, _20716_);
  and (_20735_, _13154_, _05363_);
  or (_20737_, _20664_, _04591_);
  or (_20738_, _20737_, _20735_);
  and (_20739_, _06358_, _05363_);
  or (_20740_, _20739_, _20664_);
  or (_20741_, _20740_, _04582_);
  and (_20742_, _20741_, _04589_);
  and (_20743_, _20742_, _20738_);
  and (_20744_, _20743_, _20734_);
  and (_20745_, _13160_, _05363_);
  or (_20746_, _20745_, _20664_);
  and (_20747_, _20746_, _03778_);
  or (_20748_, _20747_, _20744_);
  and (_20749_, _20748_, _04596_);
  or (_20750_, _20664_, _05601_);
  and (_20751_, _20740_, _03655_);
  and (_20752_, _20751_, _20750_);
  or (_20753_, _20752_, _20749_);
  and (_20754_, _20753_, _04594_);
  and (_20755_, _20669_, _03773_);
  and (_20756_, _20755_, _20750_);
  or (_20758_, _20756_, _03653_);
  or (_20759_, _20758_, _20754_);
  nor (_20760_, _13152_, _09268_);
  or (_20761_, _20664_, _04608_);
  or (_20762_, _20761_, _20760_);
  and (_20763_, _20762_, _04606_);
  and (_20764_, _20763_, _20759_);
  nor (_20765_, _13159_, _09268_);
  or (_20766_, _20765_, _20664_);
  and (_20767_, _20766_, _03786_);
  or (_20769_, _20767_, _03809_);
  or (_20770_, _20769_, _20764_);
  or (_20771_, _20666_, _04260_);
  and (_20772_, _20771_, _03206_);
  and (_20773_, _20772_, _20770_);
  and (_20774_, _20692_, _03205_);
  or (_20775_, _20774_, _03816_);
  or (_20776_, _20775_, _20773_);
  and (_20777_, _13217_, _05363_);
  or (_20778_, _20664_, _03820_);
  or (_20779_, _20778_, _20777_);
  and (_20780_, _20779_, _43227_);
  and (_20781_, _20780_, _20776_);
  or (_43481_, _20781_, _20663_);
  not (_20782_, \oc8051_golden_model_1.P0 [6]);
  nor (_20783_, _05363_, _20782_);
  nor (_20784_, _13235_, _09268_);
  or (_20785_, _20784_, _20783_);
  or (_20786_, _20785_, _04515_);
  and (_20787_, _05363_, \oc8051_golden_model_1.ACC [6]);
  or (_20789_, _20787_, _20783_);
  and (_20790_, _20789_, _04499_);
  nor (_20791_, _04499_, _20782_);
  or (_20792_, _20791_, _03599_);
  or (_20793_, _20792_, _20790_);
  and (_20794_, _20793_, _03516_);
  and (_20795_, _20794_, _20786_);
  nor (_20796_, _05294_, _20782_);
  and (_20797_, _13266_, _05294_);
  or (_20798_, _20797_, _20796_);
  and (_20800_, _20798_, _03515_);
  or (_20801_, _20800_, _03597_);
  or (_20802_, _20801_, _20795_);
  nor (_20803_, _05442_, _09268_);
  or (_20804_, _20803_, _20783_);
  or (_20805_, _20804_, _04524_);
  and (_20806_, _20805_, _20802_);
  or (_20807_, _20806_, _03603_);
  or (_20808_, _20789_, _03611_);
  and (_20809_, _20808_, _03512_);
  and (_20810_, _20809_, _20807_);
  and (_20811_, _13251_, _05294_);
  or (_20812_, _20811_, _20796_);
  and (_20813_, _20812_, _03511_);
  or (_20814_, _20813_, _03504_);
  or (_20815_, _20814_, _20810_);
  or (_20816_, _20796_, _13281_);
  and (_20817_, _20816_, _20798_);
  or (_20818_, _20817_, _03505_);
  and (_20819_, _20818_, _03501_);
  and (_20821_, _20819_, _20815_);
  or (_20822_, _13251_, _13248_);
  and (_20823_, _20822_, _05294_);
  or (_20824_, _20823_, _20796_);
  and (_20825_, _20824_, _03500_);
  or (_20826_, _20825_, _07441_);
  or (_20827_, _20826_, _20821_);
  or (_20828_, _20804_, _06889_);
  and (_20829_, _20828_, _20827_);
  or (_20830_, _20829_, _05969_);
  and (_20832_, _06531_, _05363_);
  or (_20833_, _20783_, _05970_);
  or (_20834_, _20833_, _20832_);
  and (_20835_, _20834_, _03275_);
  and (_20836_, _20835_, _20830_);
  and (_20837_, _06356_, \oc8051_golden_model_1.P0 [6]);
  and (_20838_, _06361_, \oc8051_golden_model_1.P2 [6]);
  or (_20839_, _20838_, _13309_);
  or (_20840_, _20839_, _20837_);
  and (_20841_, _06378_, \oc8051_golden_model_1.P1 [6]);
  and (_20842_, _06382_, \oc8051_golden_model_1.P3 [6]);
  or (_20843_, _20842_, _20841_);
  or (_20844_, _20843_, _13317_);
  or (_20845_, _20844_, _13315_);
  nor (_20846_, _20845_, _20840_);
  and (_20847_, _20846_, _13334_);
  nand (_20848_, _20847_, _13353_);
  or (_20849_, _20848_, _13308_);
  and (_20850_, _20849_, _05363_);
  or (_20851_, _20850_, _20783_);
  and (_20853_, _20851_, _03644_);
  or (_20854_, _20853_, _08861_);
  or (_20855_, _20854_, _20836_);
  and (_20856_, _13245_, _05363_);
  or (_20857_, _20783_, _04591_);
  or (_20858_, _20857_, _20856_);
  and (_20859_, _13363_, _05363_);
  or (_20860_, _20859_, _20783_);
  or (_20861_, _20860_, _04582_);
  and (_20862_, _20861_, _04589_);
  and (_20864_, _20862_, _20858_);
  and (_20865_, _20864_, _20855_);
  and (_20866_, _13374_, _05363_);
  or (_20867_, _20866_, _20783_);
  and (_20868_, _20867_, _03778_);
  or (_20869_, _20868_, _20865_);
  and (_20870_, _20869_, _04596_);
  or (_20871_, _20783_, _05491_);
  and (_20872_, _20860_, _03655_);
  and (_20873_, _20872_, _20871_);
  or (_20875_, _20873_, _20870_);
  and (_20876_, _20875_, _04594_);
  and (_20877_, _20789_, _03773_);
  and (_20878_, _20877_, _20871_);
  or (_20879_, _20878_, _03653_);
  or (_20880_, _20879_, _20876_);
  nor (_20881_, _13243_, _09268_);
  or (_20882_, _20783_, _04608_);
  or (_20883_, _20882_, _20881_);
  and (_20884_, _20883_, _04606_);
  and (_20885_, _20884_, _20880_);
  nor (_20886_, _13373_, _09268_);
  or (_20887_, _20886_, _20783_);
  and (_20888_, _20887_, _03786_);
  or (_20889_, _20888_, _03809_);
  or (_20890_, _20889_, _20885_);
  or (_20891_, _20785_, _04260_);
  and (_20892_, _20891_, _03206_);
  and (_20893_, _20892_, _20890_);
  and (_20894_, _20812_, _03205_);
  or (_20896_, _20894_, _03816_);
  or (_20897_, _20896_, _20893_);
  and (_20898_, _13425_, _05363_);
  or (_20899_, _20783_, _03820_);
  or (_20900_, _20899_, _20898_);
  and (_20901_, _20900_, _43227_);
  and (_20902_, _20901_, _20897_);
  nor (_20903_, _43227_, _20782_);
  or (_20904_, _20903_, rst);
  or (_43482_, _20904_, _20902_);
  not (_20906_, \oc8051_golden_model_1.P1 [0]);
  nor (_20907_, _43227_, _20906_);
  or (_20908_, _20907_, rst);
  nor (_20909_, _05383_, _20906_);
  and (_20910_, _12145_, _05383_);
  or (_20911_, _20910_, _20909_);
  and (_20912_, _20911_, _03778_);
  and (_20913_, _05383_, _04491_);
  or (_20914_, _20913_, _20909_);
  or (_20915_, _20914_, _06889_);
  nor (_20916_, _05744_, _09386_);
  or (_20917_, _20916_, _20909_);
  or (_20918_, _20917_, _04515_);
  and (_20919_, _05383_, \oc8051_golden_model_1.ACC [0]);
  or (_20920_, _20919_, _20909_);
  and (_20921_, _20920_, _04499_);
  nor (_20922_, _04499_, _20906_);
  or (_20923_, _20922_, _03599_);
  or (_20924_, _20923_, _20921_);
  and (_20925_, _20924_, _03516_);
  and (_20927_, _20925_, _20918_);
  nor (_20928_, _06013_, _20906_);
  and (_20929_, _12035_, _06013_);
  or (_20930_, _20929_, _20928_);
  and (_20931_, _20930_, _03515_);
  or (_20932_, _20931_, _20927_);
  and (_20933_, _20932_, _04524_);
  and (_20934_, _20914_, _03597_);
  or (_20935_, _20934_, _03603_);
  or (_20936_, _20935_, _20933_);
  or (_20938_, _20920_, _03611_);
  and (_20939_, _20938_, _03512_);
  and (_20940_, _20939_, _20936_);
  and (_20941_, _20909_, _03511_);
  or (_20942_, _20941_, _03504_);
  or (_20943_, _20942_, _20940_);
  or (_20944_, _20917_, _03505_);
  and (_20945_, _20944_, _03501_);
  and (_20946_, _20945_, _20943_);
  and (_20947_, _20078_, _06013_);
  or (_20949_, _20947_, _20928_);
  and (_20950_, _20949_, _03500_);
  or (_20951_, _20950_, _07441_);
  or (_20952_, _20951_, _20946_);
  and (_20953_, _20952_, _20915_);
  or (_20954_, _20953_, _05969_);
  and (_20955_, _06836_, _05383_);
  or (_20956_, _20909_, _05970_);
  or (_20957_, _20956_, _20955_);
  and (_20958_, _20957_, _03275_);
  and (_20959_, _20958_, _20954_);
  and (_20960_, _20114_, _05383_);
  or (_20961_, _20960_, _20909_);
  and (_20962_, _20961_, _03644_);
  or (_20963_, _20962_, _20959_);
  or (_20964_, _20963_, _08861_);
  and (_20965_, _12019_, _05383_);
  or (_20966_, _20909_, _04591_);
  or (_20967_, _20966_, _20965_);
  and (_20968_, _05383_, _06366_);
  or (_20970_, _20968_, _20909_);
  or (_20971_, _20970_, _04582_);
  and (_20972_, _20971_, _04589_);
  and (_20973_, _20972_, _20967_);
  and (_20974_, _20973_, _20964_);
  or (_20975_, _20974_, _20912_);
  and (_20976_, _20975_, _04596_);
  nand (_20977_, _20970_, _03655_);
  nor (_20978_, _20977_, _20916_);
  or (_20979_, _20978_, _20976_);
  and (_20981_, _20979_, _04594_);
  or (_20982_, _20909_, _05744_);
  and (_20983_, _20920_, _03773_);
  and (_20984_, _20983_, _20982_);
  or (_20985_, _20984_, _03653_);
  or (_20986_, _20985_, _20981_);
  nor (_20987_, _12017_, _09386_);
  or (_20988_, _20909_, _04608_);
  or (_20989_, _20988_, _20987_);
  and (_20990_, _20989_, _04606_);
  and (_20991_, _20990_, _20986_);
  nor (_20992_, _12015_, _09386_);
  or (_20993_, _20992_, _20909_);
  and (_20994_, _20993_, _03786_);
  or (_20995_, _20994_, _03809_);
  or (_20996_, _20995_, _20991_);
  or (_20997_, _20917_, _04260_);
  and (_20998_, _20997_, _03206_);
  and (_20999_, _20998_, _20996_);
  and (_21000_, _20909_, _03205_);
  or (_21002_, _21000_, _03816_);
  or (_21003_, _21002_, _20999_);
  or (_21004_, _20917_, _03820_);
  and (_21005_, _21004_, _43227_);
  and (_21006_, _21005_, _21003_);
  or (_43485_, _21006_, _20908_);
  not (_21007_, \oc8051_golden_model_1.P1 [1]);
  nor (_21008_, _05383_, _21007_);
  and (_21009_, _05383_, _05898_);
  or (_21010_, _21009_, _21008_);
  or (_21012_, _21010_, _04524_);
  or (_21013_, _05383_, \oc8051_golden_model_1.P1 [1]);
  and (_21014_, _12234_, _05383_);
  not (_21015_, _21014_);
  and (_21016_, _21015_, _21013_);
  or (_21017_, _21016_, _04515_);
  nand (_21018_, _05383_, _03320_);
  and (_21019_, _21018_, _21013_);
  and (_21020_, _21019_, _04499_);
  nor (_21021_, _04499_, _21007_);
  or (_21023_, _21021_, _03599_);
  or (_21024_, _21023_, _21020_);
  and (_21025_, _21024_, _03516_);
  and (_21026_, _21025_, _21017_);
  nor (_21027_, _06013_, _21007_);
  and (_21028_, _12238_, _06013_);
  or (_21029_, _21028_, _21027_);
  and (_21030_, _21029_, _03515_);
  or (_21031_, _21030_, _03597_);
  or (_21032_, _21031_, _21026_);
  and (_21034_, _21032_, _21012_);
  or (_21035_, _21034_, _03603_);
  or (_21036_, _21019_, _03611_);
  and (_21037_, _21036_, _03512_);
  and (_21038_, _21037_, _21035_);
  and (_21039_, _12224_, _06013_);
  or (_21040_, _21039_, _21027_);
  and (_21041_, _21040_, _03511_);
  or (_21042_, _21041_, _03504_);
  or (_21043_, _21042_, _21038_);
  and (_21045_, _21028_, _12253_);
  or (_21046_, _21027_, _03505_);
  or (_21047_, _21046_, _21045_);
  and (_21048_, _21047_, _21043_);
  and (_21049_, _21048_, _03501_);
  and (_21050_, _20206_, _06013_);
  or (_21051_, _21027_, _21050_);
  and (_21052_, _21051_, _03500_);
  or (_21053_, _21052_, _07441_);
  or (_21054_, _21053_, _21049_);
  or (_21056_, _21010_, _06889_);
  and (_21057_, _21056_, _21054_);
  or (_21058_, _21057_, _05969_);
  and (_21059_, _06835_, _05383_);
  or (_21060_, _21008_, _05970_);
  or (_21061_, _21060_, _21059_);
  and (_21062_, _21061_, _03275_);
  and (_21063_, _21062_, _21058_);
  and (_21064_, _20235_, _05383_);
  or (_21065_, _21064_, _21008_);
  and (_21067_, _21065_, _03644_);
  or (_21068_, _21067_, _21063_);
  and (_21069_, _21068_, _03651_);
  or (_21070_, _12220_, _09386_);
  and (_21071_, _21070_, _03649_);
  nand (_21072_, _05383_, _04347_);
  and (_21073_, _21072_, _03650_);
  or (_21074_, _21073_, _21071_);
  and (_21075_, _21074_, _21013_);
  or (_21076_, _21075_, _21069_);
  and (_21078_, _21076_, _04589_);
  or (_21079_, _12347_, _09386_);
  and (_21080_, _21013_, _03778_);
  and (_21081_, _21080_, _21079_);
  or (_21082_, _21081_, _21078_);
  and (_21083_, _21082_, _04596_);
  or (_21084_, _12219_, _09386_);
  and (_21085_, _21013_, _03655_);
  and (_21086_, _21085_, _21084_);
  or (_21087_, _21086_, _21083_);
  and (_21089_, _21087_, _04594_);
  or (_21090_, _21008_, _05699_);
  and (_21091_, _21019_, _03773_);
  and (_21092_, _21091_, _21090_);
  or (_21093_, _21092_, _21089_);
  and (_21094_, _21093_, _03787_);
  or (_21095_, _21072_, _05699_);
  and (_21096_, _21013_, _03653_);
  and (_21097_, _21096_, _21095_);
  or (_21098_, _21018_, _05699_);
  and (_21099_, _21013_, _03786_);
  and (_21100_, _21099_, _21098_);
  or (_21101_, _21100_, _03809_);
  or (_21102_, _21101_, _21097_);
  or (_21103_, _21102_, _21094_);
  or (_21104_, _21016_, _04260_);
  and (_21105_, _21104_, _03206_);
  and (_21106_, _21105_, _21103_);
  and (_21107_, _21040_, _03205_);
  or (_21108_, _21107_, _03816_);
  or (_21109_, _21108_, _21106_);
  or (_21110_, _21008_, _03820_);
  or (_21111_, _21110_, _21014_);
  and (_21112_, _21111_, _43227_);
  and (_21113_, _21112_, _21109_);
  nor (_21114_, _43227_, _21007_);
  or (_21115_, _21114_, rst);
  or (_43486_, _21115_, _21113_);
  not (_21116_, \oc8051_golden_model_1.P1 [2]);
  nor (_21117_, _43227_, _21116_);
  or (_21119_, _21117_, rst);
  nor (_21120_, _05383_, _21116_);
  nor (_21121_, _09386_, _05130_);
  or (_21122_, _21121_, _21120_);
  or (_21123_, _21122_, _06889_);
  or (_21124_, _21122_, _04524_);
  nor (_21125_, _12430_, _09386_);
  or (_21126_, _21125_, _21120_);
  or (_21127_, _21126_, _04515_);
  and (_21128_, _05383_, \oc8051_golden_model_1.ACC [2]);
  or (_21130_, _21128_, _21120_);
  and (_21131_, _21130_, _04499_);
  nor (_21132_, _04499_, _21116_);
  or (_21133_, _21132_, _03599_);
  or (_21134_, _21133_, _21131_);
  and (_21135_, _21134_, _03516_);
  and (_21136_, _21135_, _21127_);
  nor (_21137_, _06013_, _21116_);
  and (_21138_, _12416_, _06013_);
  or (_21139_, _21138_, _21137_);
  and (_21141_, _21139_, _03515_);
  or (_21142_, _21141_, _03597_);
  or (_21143_, _21142_, _21136_);
  and (_21144_, _21143_, _21124_);
  or (_21145_, _21144_, _03603_);
  or (_21146_, _21130_, _03611_);
  and (_21147_, _21146_, _03512_);
  and (_21148_, _21147_, _21145_);
  and (_21149_, _12414_, _06013_);
  or (_21150_, _21149_, _21137_);
  and (_21152_, _21150_, _03511_);
  or (_21153_, _21152_, _03504_);
  or (_21154_, _21153_, _21148_);
  and (_21155_, _21138_, _12447_);
  or (_21156_, _21137_, _03505_);
  or (_21157_, _21156_, _21155_);
  and (_21158_, _21157_, _03501_);
  and (_21159_, _21158_, _21154_);
  and (_21160_, _20332_, _06013_);
  or (_21161_, _21160_, _21137_);
  and (_21163_, _21161_, _03500_);
  or (_21164_, _21163_, _07441_);
  or (_21165_, _21164_, _21159_);
  and (_21166_, _21165_, _21123_);
  or (_21167_, _21166_, _05969_);
  and (_21168_, _06839_, _05383_);
  or (_21169_, _21120_, _05970_);
  or (_21170_, _21169_, _21168_);
  and (_21171_, _21170_, _03275_);
  and (_21172_, _21171_, _21167_);
  and (_21174_, _20358_, _05383_);
  or (_21175_, _21120_, _21174_);
  and (_21176_, _21175_, _03644_);
  or (_21177_, _21176_, _21172_);
  or (_21178_, _21177_, _08861_);
  and (_21179_, _12538_, _05383_);
  or (_21180_, _21120_, _04591_);
  or (_21181_, _21180_, _21179_);
  and (_21182_, _05383_, _06414_);
  or (_21183_, _21182_, _21120_);
  or (_21185_, _21183_, _04582_);
  and (_21186_, _21185_, _04589_);
  and (_21187_, _21186_, _21181_);
  and (_21188_, _21187_, _21178_);
  and (_21189_, _12544_, _05383_);
  or (_21190_, _21189_, _21120_);
  and (_21191_, _21190_, _03778_);
  or (_21192_, _21191_, _21188_);
  and (_21193_, _21192_, _04596_);
  or (_21194_, _21120_, _05793_);
  and (_21196_, _21183_, _03655_);
  and (_21197_, _21196_, _21194_);
  or (_21198_, _21197_, _21193_);
  and (_21199_, _21198_, _04594_);
  and (_21200_, _21130_, _03773_);
  and (_21201_, _21200_, _21194_);
  or (_21202_, _21201_, _03653_);
  or (_21203_, _21202_, _21199_);
  nor (_21204_, _12537_, _09386_);
  or (_21205_, _21120_, _04608_);
  or (_21207_, _21205_, _21204_);
  and (_21208_, _21207_, _04606_);
  and (_21209_, _21208_, _21203_);
  nor (_21210_, _12543_, _09386_);
  or (_21211_, _21210_, _21120_);
  and (_21212_, _21211_, _03786_);
  or (_21213_, _21212_, _03809_);
  or (_21214_, _21213_, _21209_);
  or (_21215_, _21126_, _04260_);
  and (_21216_, _21215_, _03206_);
  and (_21218_, _21216_, _21214_);
  and (_21219_, _21150_, _03205_);
  or (_21220_, _21219_, _03816_);
  or (_21221_, _21220_, _21218_);
  and (_21222_, _12600_, _05383_);
  or (_21223_, _21120_, _03820_);
  or (_21224_, _21223_, _21222_);
  and (_21225_, _21224_, _43227_);
  and (_21226_, _21225_, _21221_);
  or (_43487_, _21226_, _21119_);
  and (_21228_, _09386_, \oc8051_golden_model_1.P1 [3]);
  nor (_21229_, _09386_, _04944_);
  or (_21230_, _21229_, _21228_);
  or (_21231_, _21230_, _06889_);
  nor (_21232_, _12625_, _09386_);
  or (_21233_, _21232_, _21228_);
  or (_21234_, _21233_, _04515_);
  and (_21235_, _05383_, \oc8051_golden_model_1.ACC [3]);
  or (_21236_, _21235_, _21228_);
  and (_21237_, _21236_, _04499_);
  and (_21239_, _04500_, \oc8051_golden_model_1.P1 [3]);
  or (_21240_, _21239_, _03599_);
  or (_21241_, _21240_, _21237_);
  and (_21242_, _21241_, _03516_);
  and (_21243_, _21242_, _21234_);
  not (_21244_, _06013_);
  and (_21245_, _21244_, \oc8051_golden_model_1.P1 [3]);
  and (_21246_, _12638_, _06013_);
  or (_21247_, _21246_, _21245_);
  and (_21248_, _21247_, _03515_);
  or (_21250_, _21248_, _03597_);
  or (_21251_, _21250_, _21243_);
  or (_21252_, _21230_, _04524_);
  and (_21253_, _21252_, _21251_);
  or (_21254_, _21253_, _03603_);
  or (_21255_, _21236_, _03611_);
  and (_21256_, _21255_, _03512_);
  and (_21257_, _21256_, _21254_);
  and (_21258_, _12622_, _06013_);
  or (_21259_, _21258_, _21245_);
  and (_21261_, _21259_, _03511_);
  or (_21262_, _21261_, _03504_);
  or (_21263_, _21262_, _21257_);
  or (_21264_, _21245_, _12653_);
  and (_21265_, _21264_, _21247_);
  or (_21266_, _21265_, _03505_);
  and (_21267_, _21266_, _03501_);
  and (_21268_, _21267_, _21263_);
  and (_21269_, _20458_, _06013_);
  or (_21270_, _21269_, _21245_);
  and (_21272_, _21270_, _03500_);
  or (_21273_, _21272_, _07441_);
  or (_21274_, _21273_, _21268_);
  and (_21275_, _21274_, _21231_);
  or (_21276_, _21275_, _05969_);
  and (_21277_, _06838_, _05383_);
  or (_21278_, _21228_, _05970_);
  or (_21279_, _21278_, _21277_);
  and (_21280_, _21279_, _03275_);
  and (_21281_, _21280_, _21276_);
  and (_21283_, _20485_, _05383_);
  or (_21284_, _21228_, _21283_);
  and (_21285_, _21284_, _03644_);
  or (_21286_, _21285_, _21281_);
  or (_21287_, _21286_, _08861_);
  and (_21288_, _12746_, _05383_);
  or (_21289_, _21228_, _04591_);
  or (_21290_, _21289_, _21288_);
  and (_21291_, _05383_, _06347_);
  or (_21292_, _21291_, _21228_);
  or (_21294_, _21292_, _04582_);
  and (_21295_, _21294_, _04589_);
  and (_21296_, _21295_, _21290_);
  and (_21297_, _21296_, _21287_);
  and (_21298_, _12619_, _05383_);
  or (_21299_, _21298_, _21228_);
  and (_21300_, _21299_, _03778_);
  or (_21301_, _21300_, _21297_);
  and (_21302_, _21301_, _04596_);
  or (_21303_, _21228_, _05650_);
  and (_21305_, _21292_, _03655_);
  and (_21306_, _21305_, _21303_);
  or (_21307_, _21306_, _21302_);
  and (_21308_, _21307_, _04594_);
  and (_21309_, _21236_, _03773_);
  and (_21310_, _21309_, _21303_);
  or (_21311_, _21310_, _03653_);
  or (_21312_, _21311_, _21308_);
  nor (_21313_, _12745_, _09386_);
  or (_21314_, _21228_, _04608_);
  or (_21316_, _21314_, _21313_);
  and (_21317_, _21316_, _04606_);
  and (_21318_, _21317_, _21312_);
  nor (_21319_, _12618_, _09386_);
  or (_21320_, _21319_, _21228_);
  and (_21321_, _21320_, _03786_);
  or (_21322_, _21321_, _03809_);
  or (_21323_, _21322_, _21318_);
  or (_21324_, _21233_, _04260_);
  and (_21325_, _21324_, _03206_);
  and (_21327_, _21325_, _21323_);
  and (_21328_, _21259_, _03205_);
  or (_21329_, _21328_, _03816_);
  or (_21330_, _21329_, _21327_);
  and (_21331_, _12806_, _05383_);
  or (_21332_, _21228_, _03820_);
  or (_21333_, _21332_, _21331_);
  and (_21334_, _21333_, _43227_);
  and (_21335_, _21334_, _21330_);
  nor (_21336_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_21338_, _21336_, _05217_);
  or (_43488_, _21338_, _21335_);
  and (_21339_, _09386_, \oc8051_golden_model_1.P1 [4]);
  nor (_21340_, _05840_, _09386_);
  or (_21341_, _21340_, _21339_);
  or (_21342_, _21341_, _06889_);
  and (_21343_, _21244_, \oc8051_golden_model_1.P1 [4]);
  and (_21344_, _12853_, _06013_);
  or (_21345_, _21344_, _21343_);
  and (_21346_, _21345_, _03511_);
  nor (_21348_, _12820_, _09386_);
  or (_21349_, _21348_, _21339_);
  or (_21350_, _21349_, _04515_);
  and (_21351_, _05383_, \oc8051_golden_model_1.ACC [4]);
  or (_21352_, _21351_, _21339_);
  and (_21353_, _21352_, _04499_);
  and (_21354_, _04500_, \oc8051_golden_model_1.P1 [4]);
  or (_21355_, _21354_, _03599_);
  or (_21356_, _21355_, _21353_);
  and (_21357_, _21356_, _03516_);
  and (_21359_, _21357_, _21350_);
  and (_21360_, _12830_, _06013_);
  or (_21361_, _21360_, _21343_);
  and (_21362_, _21361_, _03515_);
  or (_21363_, _21362_, _03597_);
  or (_21364_, _21363_, _21359_);
  or (_21365_, _21341_, _04524_);
  and (_21366_, _21365_, _21364_);
  or (_21367_, _21366_, _03603_);
  or (_21368_, _21352_, _03611_);
  and (_21370_, _21368_, _03512_);
  and (_21371_, _21370_, _21367_);
  or (_21372_, _21371_, _21346_);
  and (_21373_, _21372_, _03505_);
  and (_21374_, _12861_, _06013_);
  or (_21375_, _21374_, _21343_);
  and (_21376_, _21375_, _03504_);
  or (_21377_, _21376_, _21373_);
  and (_21378_, _21377_, _03501_);
  and (_21379_, _20579_, _06013_);
  or (_21381_, _21379_, _21343_);
  and (_21382_, _21381_, _03500_);
  or (_21383_, _21382_, _07441_);
  or (_21384_, _21383_, _21378_);
  and (_21385_, _21384_, _21342_);
  or (_21386_, _21385_, _05969_);
  and (_21387_, _06843_, _05383_);
  or (_21388_, _21339_, _05970_);
  or (_21389_, _21388_, _21387_);
  and (_21390_, _21389_, _03275_);
  and (_21392_, _21390_, _21386_);
  and (_21393_, _20605_, _05383_);
  or (_21394_, _21393_, _21339_);
  and (_21395_, _21394_, _03644_);
  or (_21396_, _21395_, _08861_);
  or (_21397_, _21396_, _21392_);
  and (_21398_, _12951_, _05383_);
  or (_21399_, _21339_, _04591_);
  or (_21400_, _21399_, _21398_);
  and (_21401_, _06375_, _05383_);
  or (_21403_, _21401_, _21339_);
  or (_21404_, _21403_, _04582_);
  and (_21405_, _21404_, _04589_);
  and (_21406_, _21405_, _21400_);
  and (_21407_, _21406_, _21397_);
  and (_21408_, _12957_, _05383_);
  or (_21409_, _21408_, _21339_);
  and (_21410_, _21409_, _03778_);
  or (_21411_, _21410_, _21407_);
  and (_21412_, _21411_, _04596_);
  or (_21414_, _21339_, _05889_);
  and (_21415_, _21403_, _03655_);
  and (_21416_, _21415_, _21414_);
  or (_21417_, _21416_, _21412_);
  and (_21418_, _21417_, _04594_);
  and (_21419_, _21352_, _03773_);
  and (_21420_, _21419_, _21414_);
  or (_21421_, _21420_, _03653_);
  or (_21422_, _21421_, _21418_);
  nor (_21423_, _12949_, _09386_);
  or (_21425_, _21339_, _04608_);
  or (_21426_, _21425_, _21423_);
  and (_21427_, _21426_, _04606_);
  and (_21428_, _21427_, _21422_);
  nor (_21429_, _12956_, _09386_);
  or (_21430_, _21429_, _21339_);
  and (_21431_, _21430_, _03786_);
  or (_21432_, _21431_, _03809_);
  or (_21433_, _21432_, _21428_);
  or (_21434_, _21349_, _04260_);
  and (_21436_, _21434_, _03206_);
  and (_21437_, _21436_, _21433_);
  and (_21438_, _21345_, _03205_);
  or (_21439_, _21438_, _03816_);
  or (_21440_, _21439_, _21437_);
  and (_21441_, _13013_, _05383_);
  or (_21442_, _21339_, _03820_);
  or (_21443_, _21442_, _21441_);
  and (_21444_, _21443_, _43227_);
  and (_21445_, _21444_, _21440_);
  nor (_21447_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_21448_, _21447_, _05217_);
  or (_43489_, _21448_, _21445_);
  nor (_21449_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_21450_, _21449_, _05217_);
  and (_21451_, _09386_, \oc8051_golden_model_1.P1 [5]);
  nor (_21452_, _13035_, _09386_);
  or (_21453_, _21452_, _21451_);
  or (_21454_, _21453_, _04515_);
  and (_21455_, _05383_, \oc8051_golden_model_1.ACC [5]);
  or (_21457_, _21455_, _21451_);
  and (_21458_, _21457_, _04499_);
  and (_21459_, _04500_, \oc8051_golden_model_1.P1 [5]);
  or (_21460_, _21459_, _03599_);
  or (_21461_, _21460_, _21458_);
  and (_21462_, _21461_, _03516_);
  and (_21463_, _21462_, _21454_);
  and (_21464_, _21244_, \oc8051_golden_model_1.P1 [5]);
  and (_21465_, _13051_, _06013_);
  or (_21466_, _21465_, _21464_);
  and (_21468_, _21466_, _03515_);
  or (_21469_, _21468_, _03597_);
  or (_21470_, _21469_, _21463_);
  nor (_21471_, _05552_, _09386_);
  or (_21472_, _21471_, _21451_);
  or (_21473_, _21472_, _04524_);
  and (_21474_, _21473_, _21470_);
  or (_21475_, _21474_, _03603_);
  or (_21476_, _21457_, _03611_);
  and (_21477_, _21476_, _03512_);
  and (_21480_, _21477_, _21475_);
  and (_21481_, _13032_, _06013_);
  or (_21482_, _21481_, _21464_);
  and (_21483_, _21482_, _03511_);
  or (_21484_, _21483_, _03504_);
  or (_21485_, _21484_, _21480_);
  or (_21486_, _21464_, _13066_);
  and (_21487_, _21486_, _21466_);
  or (_21488_, _21487_, _03505_);
  and (_21489_, _21488_, _03501_);
  and (_21492_, _21489_, _21485_);
  and (_21493_, _20702_, _06013_);
  or (_21494_, _21493_, _21464_);
  and (_21495_, _21494_, _03500_);
  or (_21496_, _21495_, _07441_);
  or (_21497_, _21496_, _21492_);
  or (_21498_, _21472_, _06889_);
  and (_21499_, _21498_, _21497_);
  or (_21500_, _21499_, _05969_);
  and (_21501_, _06842_, _05383_);
  or (_21504_, _21451_, _05970_);
  or (_21505_, _21504_, _21501_);
  and (_21506_, _21505_, _03275_);
  and (_21507_, _21506_, _21500_);
  and (_21508_, _20729_, _05383_);
  or (_21509_, _21508_, _21451_);
  and (_21510_, _21509_, _03644_);
  or (_21511_, _21510_, _08861_);
  or (_21512_, _21511_, _21507_);
  and (_21513_, _13154_, _05383_);
  or (_21516_, _21451_, _04591_);
  or (_21517_, _21516_, _21513_);
  and (_21518_, _06358_, _05383_);
  or (_21519_, _21518_, _21451_);
  or (_21520_, _21519_, _04582_);
  and (_21521_, _21520_, _04589_);
  and (_21522_, _21521_, _21517_);
  and (_21523_, _21522_, _21512_);
  and (_21524_, _13160_, _05383_);
  or (_21525_, _21524_, _21451_);
  and (_21528_, _21525_, _03778_);
  or (_21529_, _21528_, _21523_);
  and (_21530_, _21529_, _04596_);
  or (_21531_, _21451_, _05601_);
  and (_21532_, _21519_, _03655_);
  and (_21533_, _21532_, _21531_);
  or (_21534_, _21533_, _21530_);
  and (_21535_, _21534_, _04594_);
  and (_21536_, _21457_, _03773_);
  and (_21537_, _21536_, _21531_);
  or (_21540_, _21537_, _03653_);
  or (_21541_, _21540_, _21535_);
  nor (_21542_, _13152_, _09386_);
  or (_21543_, _21451_, _04608_);
  or (_21544_, _21543_, _21542_);
  and (_21545_, _21544_, _04606_);
  and (_21546_, _21545_, _21541_);
  nor (_21547_, _13159_, _09386_);
  or (_21548_, _21547_, _21451_);
  and (_21549_, _21548_, _03786_);
  or (_21551_, _21549_, _03809_);
  or (_21552_, _21551_, _21546_);
  or (_21553_, _21453_, _04260_);
  and (_21554_, _21553_, _03206_);
  and (_21555_, _21554_, _21552_);
  and (_21556_, _21482_, _03205_);
  or (_21557_, _21556_, _03816_);
  or (_21558_, _21557_, _21555_);
  and (_21559_, _13217_, _05383_);
  or (_21560_, _21451_, _03820_);
  or (_21562_, _21560_, _21559_);
  and (_21563_, _21562_, _43227_);
  and (_21564_, _21563_, _21558_);
  or (_43492_, _21564_, _21450_);
  not (_21565_, \oc8051_golden_model_1.P1 [6]);
  nor (_21566_, _05383_, _21565_);
  nor (_21567_, _13235_, _09386_);
  or (_21568_, _21567_, _21566_);
  or (_21569_, _21568_, _04515_);
  and (_21570_, _05383_, \oc8051_golden_model_1.ACC [6]);
  or (_21572_, _21570_, _21566_);
  and (_21573_, _21572_, _04499_);
  nor (_21574_, _04499_, _21565_);
  or (_21575_, _21574_, _03599_);
  or (_21576_, _21575_, _21573_);
  and (_21577_, _21576_, _03516_);
  and (_21578_, _21577_, _21569_);
  nor (_21579_, _06013_, _21565_);
  and (_21580_, _13266_, _06013_);
  or (_21581_, _21580_, _21579_);
  and (_21583_, _21581_, _03515_);
  or (_21584_, _21583_, _03597_);
  or (_21585_, _21584_, _21578_);
  nor (_21586_, _05442_, _09386_);
  or (_21587_, _21586_, _21566_);
  or (_21588_, _21587_, _04524_);
  and (_21589_, _21588_, _21585_);
  or (_21590_, _21589_, _03603_);
  or (_21591_, _21572_, _03611_);
  and (_21592_, _21591_, _03512_);
  and (_21594_, _21592_, _21590_);
  and (_21595_, _13251_, _06013_);
  or (_21596_, _21595_, _21579_);
  and (_21597_, _21596_, _03511_);
  or (_21598_, _21597_, _03504_);
  or (_21599_, _21598_, _21594_);
  or (_21600_, _21579_, _13281_);
  and (_21601_, _21600_, _21581_);
  or (_21602_, _21601_, _03505_);
  and (_21603_, _21602_, _03501_);
  and (_21605_, _21603_, _21599_);
  and (_21606_, _20822_, _06013_);
  or (_21607_, _21606_, _21579_);
  and (_21608_, _21607_, _03500_);
  or (_21609_, _21608_, _07441_);
  or (_21610_, _21609_, _21605_);
  or (_21611_, _21587_, _06889_);
  and (_21612_, _21611_, _21610_);
  or (_21613_, _21612_, _05969_);
  and (_21614_, _06531_, _05383_);
  or (_21616_, _21566_, _05970_);
  or (_21617_, _21616_, _21614_);
  and (_21618_, _21617_, _03275_);
  and (_21619_, _21618_, _21613_);
  and (_21620_, _20849_, _05383_);
  or (_21621_, _21620_, _21566_);
  and (_21622_, _21621_, _03644_);
  or (_21623_, _21622_, _08861_);
  or (_21624_, _21623_, _21619_);
  and (_21625_, _13245_, _05383_);
  or (_21627_, _21566_, _04591_);
  or (_21628_, _21627_, _21625_);
  and (_21629_, _13363_, _05383_);
  or (_21630_, _21629_, _21566_);
  or (_21631_, _21630_, _04582_);
  and (_21632_, _21631_, _04589_);
  and (_21633_, _21632_, _21628_);
  and (_21634_, _21633_, _21624_);
  and (_21635_, _13374_, _05383_);
  or (_21636_, _21635_, _21566_);
  and (_21638_, _21636_, _03778_);
  or (_21639_, _21638_, _21634_);
  and (_21640_, _21639_, _04596_);
  or (_21641_, _21566_, _05491_);
  and (_21642_, _21630_, _03655_);
  and (_21643_, _21642_, _21641_);
  or (_21644_, _21643_, _21640_);
  and (_21645_, _21644_, _04594_);
  and (_21646_, _21572_, _03773_);
  and (_21647_, _21646_, _21641_);
  or (_21649_, _21647_, _03653_);
  or (_21650_, _21649_, _21645_);
  nor (_21651_, _13243_, _09386_);
  or (_21652_, _21566_, _04608_);
  or (_21653_, _21652_, _21651_);
  and (_21654_, _21653_, _04606_);
  and (_21655_, _21654_, _21650_);
  nor (_21656_, _13373_, _09386_);
  or (_21657_, _21656_, _21566_);
  and (_21658_, _21657_, _03786_);
  or (_21660_, _21658_, _03809_);
  or (_21661_, _21660_, _21655_);
  or (_21662_, _21568_, _04260_);
  and (_21663_, _21662_, _03206_);
  and (_21664_, _21663_, _21661_);
  and (_21665_, _21596_, _03205_);
  or (_21666_, _21665_, _03816_);
  or (_21667_, _21666_, _21664_);
  and (_21668_, _13425_, _05383_);
  or (_21669_, _21566_, _03820_);
  or (_21671_, _21669_, _21668_);
  and (_21672_, _21671_, _43227_);
  and (_21673_, _21672_, _21667_);
  nor (_21674_, _43227_, _21565_);
  or (_21675_, _21674_, rst);
  or (_43493_, _21675_, _21673_);
  not (_21676_, \oc8051_golden_model_1.P2 [0]);
  nor (_21677_, _43227_, _21676_);
  or (_21678_, _21677_, rst);
  nor (_21679_, _05386_, _21676_);
  and (_21681_, _12145_, _05386_);
  or (_21682_, _21681_, _21679_);
  and (_21683_, _21682_, _03778_);
  and (_21684_, _05386_, _04491_);
  or (_21685_, _21684_, _21679_);
  or (_21686_, _21685_, _06889_);
  nor (_21687_, _05744_, _09486_);
  or (_21688_, _21687_, _21679_);
  or (_21689_, _21688_, _04515_);
  and (_21690_, _05386_, \oc8051_golden_model_1.ACC [0]);
  or (_21692_, _21690_, _21679_);
  and (_21693_, _21692_, _04499_);
  nor (_21694_, _04499_, _21676_);
  or (_21695_, _21694_, _03599_);
  or (_21696_, _21695_, _21693_);
  and (_21697_, _21696_, _03516_);
  and (_21698_, _21697_, _21689_);
  nor (_21699_, _06009_, _21676_);
  and (_21700_, _12035_, _06009_);
  or (_21701_, _21700_, _21699_);
  and (_21703_, _21701_, _03515_);
  or (_21704_, _21703_, _21698_);
  and (_21705_, _21704_, _04524_);
  and (_21706_, _21685_, _03597_);
  or (_21707_, _21706_, _03603_);
  or (_21708_, _21707_, _21705_);
  or (_21709_, _21692_, _03611_);
  and (_21710_, _21709_, _03512_);
  and (_21711_, _21710_, _21708_);
  and (_21712_, _21679_, _03511_);
  or (_21714_, _21712_, _03504_);
  or (_21715_, _21714_, _21711_);
  or (_21716_, _21688_, _03505_);
  and (_21717_, _21716_, _03501_);
  and (_21718_, _21717_, _21715_);
  and (_21719_, _20078_, _06009_);
  or (_21720_, _21719_, _21699_);
  and (_21721_, _21720_, _03500_);
  or (_21722_, _21721_, _07441_);
  or (_21723_, _21722_, _21718_);
  and (_21725_, _21723_, _21686_);
  or (_21726_, _21725_, _05969_);
  and (_21727_, _06836_, _05386_);
  or (_21728_, _21679_, _05970_);
  or (_21729_, _21728_, _21727_);
  and (_21730_, _21729_, _03275_);
  and (_21731_, _21730_, _21726_);
  and (_21732_, _20114_, _05386_);
  or (_21733_, _21732_, _21679_);
  and (_21734_, _21733_, _03644_);
  or (_21736_, _21734_, _21731_);
  or (_21737_, _21736_, _08861_);
  and (_21738_, _12019_, _05386_);
  or (_21739_, _21679_, _04591_);
  or (_21740_, _21739_, _21738_);
  and (_21741_, _05386_, _06366_);
  or (_21742_, _21741_, _21679_);
  or (_21743_, _21742_, _04582_);
  and (_21744_, _21743_, _04589_);
  and (_21745_, _21744_, _21740_);
  and (_21747_, _21745_, _21737_);
  or (_21748_, _21747_, _21683_);
  and (_21749_, _21748_, _04596_);
  nand (_21750_, _21742_, _03655_);
  nor (_21751_, _21750_, _21687_);
  or (_21752_, _21751_, _21749_);
  and (_21753_, _21752_, _04594_);
  or (_21754_, _21679_, _05744_);
  and (_21755_, _21692_, _03773_);
  and (_21756_, _21755_, _21754_);
  or (_21758_, _21756_, _03653_);
  or (_21759_, _21758_, _21753_);
  nor (_21760_, _12017_, _09486_);
  or (_21761_, _21679_, _04608_);
  or (_21762_, _21761_, _21760_);
  and (_21763_, _21762_, _04606_);
  and (_21764_, _21763_, _21759_);
  nor (_21765_, _12015_, _09486_);
  or (_21766_, _21765_, _21679_);
  and (_21767_, _21766_, _03786_);
  or (_21769_, _21767_, _03809_);
  or (_21770_, _21769_, _21764_);
  or (_21771_, _21688_, _04260_);
  and (_21772_, _21771_, _03206_);
  and (_21773_, _21772_, _21770_);
  and (_21774_, _21679_, _03205_);
  or (_21775_, _21774_, _03816_);
  or (_21776_, _21775_, _21773_);
  or (_21777_, _21688_, _03820_);
  and (_21778_, _21777_, _43227_);
  and (_21780_, _21778_, _21776_);
  or (_43494_, _21780_, _21678_);
  not (_21781_, \oc8051_golden_model_1.P2 [1]);
  nor (_21782_, _05386_, _21781_);
  and (_21783_, _05386_, _05898_);
  or (_21784_, _21783_, _21782_);
  or (_21785_, _21784_, _04524_);
  or (_21786_, _05386_, \oc8051_golden_model_1.P2 [1]);
  and (_21787_, _12234_, _05386_);
  not (_21788_, _21787_);
  and (_21790_, _21788_, _21786_);
  or (_21791_, _21790_, _04515_);
  nand (_21792_, _05386_, _03320_);
  and (_21793_, _21792_, _21786_);
  and (_21794_, _21793_, _04499_);
  nor (_21795_, _04499_, _21781_);
  or (_21796_, _21795_, _03599_);
  or (_21797_, _21796_, _21794_);
  and (_21798_, _21797_, _03516_);
  and (_21799_, _21798_, _21791_);
  nor (_21801_, _06009_, _21781_);
  and (_21802_, _12238_, _06009_);
  or (_21803_, _21802_, _21801_);
  and (_21804_, _21803_, _03515_);
  or (_21805_, _21804_, _03597_);
  or (_21806_, _21805_, _21799_);
  and (_21807_, _21806_, _21785_);
  or (_21808_, _21807_, _03603_);
  or (_21809_, _21793_, _03611_);
  and (_21810_, _21809_, _03512_);
  and (_21812_, _21810_, _21808_);
  and (_21813_, _12224_, _06009_);
  or (_21814_, _21813_, _21801_);
  and (_21815_, _21814_, _03511_);
  or (_21816_, _21815_, _03504_);
  or (_21817_, _21816_, _21812_);
  and (_21818_, _21802_, _12253_);
  or (_21819_, _21801_, _03505_);
  or (_21820_, _21819_, _21818_);
  and (_21821_, _21820_, _21817_);
  and (_21823_, _21821_, _03501_);
  and (_21824_, _20206_, _06009_);
  or (_21825_, _21801_, _21824_);
  and (_21826_, _21825_, _03500_);
  or (_21827_, _21826_, _07441_);
  or (_21828_, _21827_, _21823_);
  or (_21829_, _21784_, _06889_);
  and (_21830_, _21829_, _21828_);
  or (_21831_, _21830_, _05969_);
  and (_21832_, _06835_, _05386_);
  or (_21834_, _21782_, _05970_);
  or (_21835_, _21834_, _21832_);
  and (_21836_, _21835_, _03275_);
  and (_21837_, _21836_, _21831_);
  and (_21838_, _20235_, _05386_);
  or (_21839_, _21838_, _21782_);
  and (_21840_, _21839_, _03644_);
  or (_21841_, _21840_, _21837_);
  and (_21842_, _21841_, _03651_);
  or (_21843_, _12220_, _09486_);
  and (_21845_, _21843_, _03649_);
  nand (_21846_, _05386_, _04347_);
  and (_21847_, _21846_, _03650_);
  or (_21848_, _21847_, _21845_);
  and (_21849_, _21848_, _21786_);
  or (_21850_, _21849_, _21842_);
  and (_21851_, _21850_, _04589_);
  or (_21852_, _12347_, _09486_);
  and (_21853_, _21786_, _03778_);
  and (_21854_, _21853_, _21852_);
  or (_21856_, _21854_, _21851_);
  and (_21857_, _21856_, _04596_);
  or (_21858_, _12219_, _09486_);
  and (_21859_, _21786_, _03655_);
  and (_21860_, _21859_, _21858_);
  or (_21861_, _21860_, _21857_);
  and (_21862_, _21861_, _04594_);
  or (_21863_, _21782_, _05699_);
  and (_21864_, _21793_, _03773_);
  and (_21865_, _21864_, _21863_);
  or (_21867_, _21865_, _21862_);
  and (_21868_, _21867_, _03787_);
  or (_21869_, _21846_, _05699_);
  and (_21870_, _21786_, _03653_);
  and (_21871_, _21870_, _21869_);
  or (_21872_, _21792_, _05699_);
  and (_21873_, _21786_, _03786_);
  and (_21874_, _21873_, _21872_);
  or (_21875_, _21874_, _03809_);
  or (_21876_, _21875_, _21871_);
  or (_21878_, _21876_, _21868_);
  or (_21879_, _21790_, _04260_);
  and (_21880_, _21879_, _03206_);
  and (_21881_, _21880_, _21878_);
  and (_21882_, _21814_, _03205_);
  or (_21883_, _21882_, _03816_);
  or (_21884_, _21883_, _21881_);
  or (_21885_, _21782_, _03820_);
  or (_21886_, _21885_, _21787_);
  and (_21887_, _21886_, _43227_);
  and (_21889_, _21887_, _21884_);
  nor (_21890_, _43227_, _21781_);
  or (_21891_, _21890_, rst);
  or (_43495_, _21891_, _21889_);
  not (_21892_, \oc8051_golden_model_1.P2 [2]);
  nor (_21893_, _43227_, _21892_);
  or (_21894_, _21893_, rst);
  nor (_21895_, _05386_, _21892_);
  nor (_21896_, _09486_, _05130_);
  or (_21897_, _21896_, _21895_);
  or (_21899_, _21897_, _06889_);
  or (_21900_, _21897_, _04524_);
  nor (_21901_, _12430_, _09486_);
  or (_21902_, _21901_, _21895_);
  or (_21903_, _21902_, _04515_);
  and (_21904_, _05386_, \oc8051_golden_model_1.ACC [2]);
  or (_21905_, _21904_, _21895_);
  and (_21906_, _21905_, _04499_);
  nor (_21907_, _04499_, _21892_);
  or (_21908_, _21907_, _03599_);
  or (_21910_, _21908_, _21906_);
  and (_21911_, _21910_, _03516_);
  and (_21912_, _21911_, _21903_);
  nor (_21913_, _06009_, _21892_);
  and (_21914_, _12416_, _06009_);
  or (_21915_, _21914_, _21913_);
  and (_21916_, _21915_, _03515_);
  or (_21917_, _21916_, _03597_);
  or (_21918_, _21917_, _21912_);
  and (_21919_, _21918_, _21900_);
  or (_21921_, _21919_, _03603_);
  or (_21922_, _21905_, _03611_);
  and (_21923_, _21922_, _03512_);
  and (_21924_, _21923_, _21921_);
  and (_21925_, _12414_, _06009_);
  or (_21926_, _21925_, _21913_);
  and (_21927_, _21926_, _03511_);
  or (_21928_, _21927_, _03504_);
  or (_21929_, _21928_, _21924_);
  and (_21930_, _21914_, _12447_);
  or (_21932_, _21913_, _03505_);
  or (_21933_, _21932_, _21930_);
  and (_21934_, _21933_, _03501_);
  and (_21935_, _21934_, _21929_);
  and (_21936_, _20332_, _06009_);
  or (_21937_, _21936_, _21913_);
  and (_21938_, _21937_, _03500_);
  or (_21939_, _21938_, _07441_);
  or (_21940_, _21939_, _21935_);
  and (_21941_, _21940_, _21899_);
  or (_21943_, _21941_, _05969_);
  and (_21944_, _06839_, _05386_);
  or (_21945_, _21895_, _05970_);
  or (_21946_, _21945_, _21944_);
  and (_21947_, _21946_, _03275_);
  and (_21948_, _21947_, _21943_);
  and (_21949_, _20358_, _05386_);
  or (_21950_, _21895_, _21949_);
  and (_21951_, _21950_, _03644_);
  or (_21952_, _21951_, _21948_);
  or (_21954_, _21952_, _08861_);
  and (_21955_, _12538_, _05386_);
  or (_21956_, _21895_, _04591_);
  or (_21957_, _21956_, _21955_);
  and (_21958_, _05386_, _06414_);
  or (_21959_, _21958_, _21895_);
  or (_21960_, _21959_, _04582_);
  and (_21961_, _21960_, _04589_);
  and (_21962_, _21961_, _21957_);
  and (_21963_, _21962_, _21954_);
  and (_21965_, _12544_, _05386_);
  or (_21966_, _21965_, _21895_);
  and (_21967_, _21966_, _03778_);
  or (_21968_, _21967_, _21963_);
  and (_21969_, _21968_, _04596_);
  or (_21970_, _21895_, _05793_);
  and (_21971_, _21959_, _03655_);
  and (_21972_, _21971_, _21970_);
  or (_21973_, _21972_, _21969_);
  and (_21974_, _21973_, _04594_);
  and (_21976_, _21905_, _03773_);
  and (_21977_, _21976_, _21970_);
  or (_21978_, _21977_, _03653_);
  or (_21979_, _21978_, _21974_);
  nor (_21980_, _12537_, _09486_);
  or (_21981_, _21895_, _04608_);
  or (_21982_, _21981_, _21980_);
  and (_21983_, _21982_, _04606_);
  and (_21984_, _21983_, _21979_);
  nor (_21985_, _12543_, _09486_);
  or (_21987_, _21985_, _21895_);
  and (_21988_, _21987_, _03786_);
  or (_21989_, _21988_, _03809_);
  or (_21990_, _21989_, _21984_);
  or (_21991_, _21902_, _04260_);
  and (_21992_, _21991_, _03206_);
  and (_21993_, _21992_, _21990_);
  and (_21994_, _21926_, _03205_);
  or (_21995_, _21994_, _03816_);
  or (_21996_, _21995_, _21993_);
  and (_21998_, _12600_, _05386_);
  or (_21999_, _21895_, _03820_);
  or (_22000_, _21999_, _21998_);
  and (_22001_, _22000_, _43227_);
  and (_22002_, _22001_, _21996_);
  or (_43496_, _22002_, _21894_);
  and (_22003_, _09486_, \oc8051_golden_model_1.P2 [3]);
  nor (_22004_, _09486_, _04944_);
  or (_22005_, _22004_, _22003_);
  or (_22006_, _22005_, _06889_);
  nor (_22008_, _12625_, _09486_);
  or (_22009_, _22008_, _22003_);
  or (_22010_, _22009_, _04515_);
  and (_22011_, _05386_, \oc8051_golden_model_1.ACC [3]);
  or (_22012_, _22011_, _22003_);
  and (_22013_, _22012_, _04499_);
  and (_22014_, _04500_, \oc8051_golden_model_1.P2 [3]);
  or (_22015_, _22014_, _03599_);
  or (_22016_, _22015_, _22013_);
  and (_22017_, _22016_, _03516_);
  and (_22019_, _22017_, _22010_);
  not (_22020_, _06009_);
  and (_22021_, _22020_, \oc8051_golden_model_1.P2 [3]);
  and (_22022_, _12638_, _06009_);
  or (_22023_, _22022_, _22021_);
  and (_22024_, _22023_, _03515_);
  or (_22025_, _22024_, _03597_);
  or (_22026_, _22025_, _22019_);
  or (_22027_, _22005_, _04524_);
  and (_22028_, _22027_, _22026_);
  or (_22030_, _22028_, _03603_);
  or (_22031_, _22012_, _03611_);
  and (_22032_, _22031_, _03512_);
  and (_22033_, _22032_, _22030_);
  and (_22034_, _12622_, _06009_);
  or (_22035_, _22034_, _22021_);
  and (_22036_, _22035_, _03511_);
  or (_22037_, _22036_, _03504_);
  or (_22038_, _22037_, _22033_);
  or (_22039_, _22021_, _12653_);
  and (_22040_, _22039_, _22023_);
  or (_22041_, _22040_, _03505_);
  and (_22042_, _22041_, _03501_);
  and (_22043_, _22042_, _22038_);
  and (_22044_, _20458_, _06009_);
  or (_22045_, _22044_, _22021_);
  and (_22046_, _22045_, _03500_);
  or (_22047_, _22046_, _07441_);
  or (_22048_, _22047_, _22043_);
  and (_22049_, _22048_, _22006_);
  or (_22052_, _22049_, _05969_);
  and (_22053_, _06838_, _05386_);
  or (_22054_, _22003_, _05970_);
  or (_22055_, _22054_, _22053_);
  and (_22056_, _22055_, _03275_);
  and (_22057_, _22056_, _22052_);
  and (_22058_, _20485_, _05386_);
  or (_22059_, _22003_, _22058_);
  and (_22060_, _22059_, _03644_);
  or (_22061_, _22060_, _22057_);
  or (_22063_, _22061_, _08861_);
  and (_22064_, _12746_, _05386_);
  or (_22065_, _22003_, _04591_);
  or (_22066_, _22065_, _22064_);
  and (_22067_, _05386_, _06347_);
  or (_22068_, _22067_, _22003_);
  or (_22069_, _22068_, _04582_);
  and (_22070_, _22069_, _04589_);
  and (_22071_, _22070_, _22066_);
  and (_22072_, _22071_, _22063_);
  and (_22074_, _12619_, _05386_);
  or (_22075_, _22074_, _22003_);
  and (_22076_, _22075_, _03778_);
  or (_22077_, _22076_, _22072_);
  and (_22078_, _22077_, _04596_);
  or (_22079_, _22003_, _05650_);
  and (_22080_, _22068_, _03655_);
  and (_22081_, _22080_, _22079_);
  or (_22082_, _22081_, _22078_);
  and (_22083_, _22082_, _04594_);
  and (_22085_, _22012_, _03773_);
  and (_22086_, _22085_, _22079_);
  or (_22087_, _22086_, _03653_);
  or (_22088_, _22087_, _22083_);
  nor (_22089_, _12745_, _09486_);
  or (_22090_, _22003_, _04608_);
  or (_22091_, _22090_, _22089_);
  and (_22092_, _22091_, _04606_);
  and (_22093_, _22092_, _22088_);
  nor (_22094_, _12618_, _09486_);
  or (_22096_, _22094_, _22003_);
  and (_22097_, _22096_, _03786_);
  or (_22098_, _22097_, _03809_);
  or (_22099_, _22098_, _22093_);
  or (_22100_, _22009_, _04260_);
  and (_22101_, _22100_, _03206_);
  and (_22102_, _22101_, _22099_);
  and (_22103_, _22035_, _03205_);
  or (_22104_, _22103_, _03816_);
  or (_22105_, _22104_, _22102_);
  and (_22107_, _12806_, _05386_);
  or (_22108_, _22003_, _03820_);
  or (_22109_, _22108_, _22107_);
  and (_22110_, _22109_, _43227_);
  and (_22111_, _22110_, _22105_);
  nor (_22112_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_22113_, _22112_, _05217_);
  or (_43497_, _22113_, _22111_);
  and (_22114_, _09486_, \oc8051_golden_model_1.P2 [4]);
  nor (_22115_, _05840_, _09486_);
  or (_22117_, _22115_, _22114_);
  or (_22118_, _22117_, _06889_);
  and (_22119_, _22020_, \oc8051_golden_model_1.P2 [4]);
  and (_22120_, _12853_, _06009_);
  or (_22121_, _22120_, _22119_);
  and (_22122_, _22121_, _03511_);
  nor (_22123_, _12820_, _09486_);
  or (_22124_, _22123_, _22114_);
  or (_22125_, _22124_, _04515_);
  and (_22126_, _05386_, \oc8051_golden_model_1.ACC [4]);
  or (_22128_, _22126_, _22114_);
  and (_22129_, _22128_, _04499_);
  and (_22130_, _04500_, \oc8051_golden_model_1.P2 [4]);
  or (_22131_, _22130_, _03599_);
  or (_22132_, _22131_, _22129_);
  and (_22133_, _22132_, _03516_);
  and (_22134_, _22133_, _22125_);
  and (_22135_, _12830_, _06009_);
  or (_22136_, _22135_, _22119_);
  and (_22137_, _22136_, _03515_);
  or (_22139_, _22137_, _03597_);
  or (_22140_, _22139_, _22134_);
  or (_22141_, _22117_, _04524_);
  and (_22142_, _22141_, _22140_);
  or (_22143_, _22142_, _03603_);
  or (_22144_, _22128_, _03611_);
  and (_22145_, _22144_, _03512_);
  and (_22146_, _22145_, _22143_);
  or (_22147_, _22146_, _22122_);
  and (_22148_, _22147_, _03505_);
  and (_22150_, _12861_, _06009_);
  or (_22151_, _22150_, _22119_);
  and (_22152_, _22151_, _03504_);
  or (_22153_, _22152_, _22148_);
  and (_22154_, _22153_, _03501_);
  and (_22155_, _20579_, _06009_);
  or (_22156_, _22155_, _22119_);
  and (_22157_, _22156_, _03500_);
  or (_22158_, _22157_, _07441_);
  or (_22159_, _22158_, _22154_);
  and (_22161_, _22159_, _22118_);
  or (_22162_, _22161_, _05969_);
  and (_22163_, _06843_, _05386_);
  or (_22164_, _22114_, _05970_);
  or (_22165_, _22164_, _22163_);
  and (_22166_, _22165_, _03275_);
  and (_22167_, _22166_, _22162_);
  and (_22168_, _20605_, _05386_);
  or (_22169_, _22168_, _22114_);
  and (_22170_, _22169_, _03644_);
  or (_22172_, _22170_, _08861_);
  or (_22173_, _22172_, _22167_);
  and (_22174_, _12951_, _05386_);
  or (_22175_, _22114_, _04591_);
  or (_22176_, _22175_, _22174_);
  and (_22177_, _06375_, _05386_);
  or (_22178_, _22177_, _22114_);
  or (_22179_, _22178_, _04582_);
  and (_22180_, _22179_, _04589_);
  and (_22181_, _22180_, _22176_);
  and (_22183_, _22181_, _22173_);
  and (_22184_, _12957_, _05386_);
  or (_22185_, _22184_, _22114_);
  and (_22186_, _22185_, _03778_);
  or (_22187_, _22186_, _22183_);
  and (_22188_, _22187_, _04596_);
  or (_22189_, _22114_, _05889_);
  and (_22190_, _22178_, _03655_);
  and (_22191_, _22190_, _22189_);
  or (_22192_, _22191_, _22188_);
  and (_22194_, _22192_, _04594_);
  and (_22195_, _22128_, _03773_);
  and (_22196_, _22195_, _22189_);
  or (_22197_, _22196_, _03653_);
  or (_22198_, _22197_, _22194_);
  nor (_22199_, _12949_, _09486_);
  or (_22200_, _22114_, _04608_);
  or (_22201_, _22200_, _22199_);
  and (_22202_, _22201_, _04606_);
  and (_22203_, _22202_, _22198_);
  nor (_22205_, _12956_, _09486_);
  or (_22206_, _22205_, _22114_);
  and (_22207_, _22206_, _03786_);
  or (_22208_, _22207_, _03809_);
  or (_22209_, _22208_, _22203_);
  or (_22210_, _22124_, _04260_);
  and (_22211_, _22210_, _03206_);
  and (_22212_, _22211_, _22209_);
  and (_22213_, _22121_, _03205_);
  or (_22214_, _22213_, _03816_);
  or (_22216_, _22214_, _22212_);
  and (_22217_, _13013_, _05386_);
  or (_22218_, _22114_, _03820_);
  or (_22219_, _22218_, _22217_);
  and (_22220_, _22219_, _43227_);
  and (_22221_, _22220_, _22216_);
  nor (_22222_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_22223_, _22222_, _05217_);
  or (_43498_, _22223_, _22221_);
  and (_22224_, _09486_, \oc8051_golden_model_1.P2 [5]);
  nor (_22226_, _13035_, _09486_);
  or (_22227_, _22226_, _22224_);
  or (_22228_, _22227_, _04515_);
  and (_22229_, _05386_, \oc8051_golden_model_1.ACC [5]);
  or (_22230_, _22229_, _22224_);
  and (_22231_, _22230_, _04499_);
  and (_22232_, _04500_, \oc8051_golden_model_1.P2 [5]);
  or (_22233_, _22232_, _03599_);
  or (_22234_, _22233_, _22231_);
  and (_22235_, _22234_, _03516_);
  and (_22237_, _22235_, _22228_);
  and (_22238_, _22020_, \oc8051_golden_model_1.P2 [5]);
  and (_22239_, _13051_, _06009_);
  or (_22240_, _22239_, _22238_);
  and (_22241_, _22240_, _03515_);
  or (_22242_, _22241_, _03597_);
  or (_22243_, _22242_, _22237_);
  nor (_22244_, _05552_, _09486_);
  or (_22245_, _22244_, _22224_);
  or (_22246_, _22245_, _04524_);
  and (_22248_, _22246_, _22243_);
  or (_22249_, _22248_, _03603_);
  or (_22250_, _22230_, _03611_);
  and (_22251_, _22250_, _03512_);
  and (_22252_, _22251_, _22249_);
  and (_22253_, _13032_, _06009_);
  or (_22254_, _22253_, _22238_);
  and (_22255_, _22254_, _03511_);
  or (_22256_, _22255_, _03504_);
  or (_22257_, _22256_, _22252_);
  or (_22259_, _22238_, _13066_);
  and (_22260_, _22259_, _22240_);
  or (_22261_, _22260_, _03505_);
  and (_22262_, _22261_, _03501_);
  and (_22263_, _22262_, _22257_);
  and (_22264_, _20702_, _06009_);
  or (_22265_, _22264_, _22238_);
  and (_22266_, _22265_, _03500_);
  or (_22267_, _22266_, _07441_);
  or (_22268_, _22267_, _22263_);
  or (_22270_, _22245_, _06889_);
  and (_22271_, _22270_, _22268_);
  or (_22272_, _22271_, _05969_);
  and (_22273_, _06842_, _05386_);
  or (_22274_, _22224_, _05970_);
  or (_22275_, _22274_, _22273_);
  and (_22276_, _22275_, _03275_);
  and (_22277_, _22276_, _22272_);
  and (_22278_, _20729_, _05386_);
  or (_22279_, _22278_, _22224_);
  and (_22281_, _22279_, _03644_);
  or (_22282_, _22281_, _08861_);
  or (_22283_, _22282_, _22277_);
  and (_22284_, _13154_, _05386_);
  or (_22285_, _22224_, _04591_);
  or (_22286_, _22285_, _22284_);
  and (_22287_, _06358_, _05386_);
  or (_22288_, _22287_, _22224_);
  or (_22289_, _22288_, _04582_);
  and (_22290_, _22289_, _04589_);
  and (_22292_, _22290_, _22286_);
  and (_22293_, _22292_, _22283_);
  and (_22294_, _13160_, _05386_);
  or (_22295_, _22294_, _22224_);
  and (_22296_, _22295_, _03778_);
  or (_22297_, _22296_, _22293_);
  and (_22298_, _22297_, _04596_);
  or (_22299_, _22224_, _05601_);
  and (_22300_, _22288_, _03655_);
  and (_22301_, _22300_, _22299_);
  or (_22303_, _22301_, _22298_);
  and (_22304_, _22303_, _04594_);
  and (_22305_, _22230_, _03773_);
  and (_22306_, _22305_, _22299_);
  or (_22307_, _22306_, _03653_);
  or (_22308_, _22307_, _22304_);
  nor (_22309_, _13152_, _09486_);
  or (_22310_, _22224_, _04608_);
  or (_22311_, _22310_, _22309_);
  and (_22312_, _22311_, _04606_);
  and (_22315_, _22312_, _22308_);
  nor (_22316_, _13159_, _09486_);
  or (_22317_, _22316_, _22224_);
  and (_22318_, _22317_, _03786_);
  or (_22319_, _22318_, _03809_);
  or (_22320_, _22319_, _22315_);
  or (_22321_, _22227_, _04260_);
  and (_22322_, _22321_, _03206_);
  and (_22323_, _22322_, _22320_);
  and (_22324_, _22254_, _03205_);
  or (_22326_, _22324_, _03816_);
  or (_22327_, _22326_, _22323_);
  and (_22328_, _13217_, _05386_);
  or (_22329_, _22224_, _03820_);
  or (_22330_, _22329_, _22328_);
  and (_22331_, _22330_, _43227_);
  and (_22332_, _22331_, _22327_);
  nor (_22333_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_22334_, _22333_, _05217_);
  or (_43499_, _22334_, _22332_);
  not (_22336_, \oc8051_golden_model_1.P2 [6]);
  nor (_22337_, _43227_, _22336_);
  or (_22338_, _22337_, rst);
  nor (_22339_, _05386_, _22336_);
  nor (_22340_, _13235_, _09486_);
  or (_22341_, _22340_, _22339_);
  or (_22342_, _22341_, _04515_);
  and (_22343_, _05386_, \oc8051_golden_model_1.ACC [6]);
  or (_22344_, _22343_, _22339_);
  and (_22345_, _22344_, _04499_);
  nor (_22347_, _04499_, _22336_);
  or (_22348_, _22347_, _03599_);
  or (_22349_, _22348_, _22345_);
  and (_22350_, _22349_, _03516_);
  and (_22351_, _22350_, _22342_);
  nor (_22352_, _06009_, _22336_);
  and (_22353_, _13266_, _06009_);
  or (_22354_, _22353_, _22352_);
  and (_22355_, _22354_, _03515_);
  or (_22356_, _22355_, _03597_);
  or (_22358_, _22356_, _22351_);
  nor (_22359_, _05442_, _09486_);
  or (_22360_, _22359_, _22339_);
  or (_22361_, _22360_, _04524_);
  and (_22362_, _22361_, _22358_);
  or (_22363_, _22362_, _03603_);
  or (_22364_, _22344_, _03611_);
  and (_22365_, _22364_, _03512_);
  and (_22366_, _22365_, _22363_);
  and (_22367_, _13251_, _06009_);
  or (_22369_, _22367_, _22352_);
  and (_22370_, _22369_, _03511_);
  or (_22371_, _22370_, _03504_);
  or (_22372_, _22371_, _22366_);
  or (_22373_, _22352_, _13281_);
  and (_22374_, _22373_, _22354_);
  or (_22375_, _22374_, _03505_);
  and (_22376_, _22375_, _03501_);
  and (_22377_, _22376_, _22372_);
  and (_22378_, _20822_, _06009_);
  or (_22380_, _22378_, _22352_);
  and (_22381_, _22380_, _03500_);
  or (_22382_, _22381_, _07441_);
  or (_22383_, _22382_, _22377_);
  or (_22384_, _22360_, _06889_);
  and (_22385_, _22384_, _22383_);
  or (_22386_, _22385_, _05969_);
  and (_22387_, _06531_, _05386_);
  or (_22388_, _22339_, _05970_);
  or (_22389_, _22388_, _22387_);
  and (_22391_, _22389_, _03275_);
  and (_22392_, _22391_, _22386_);
  and (_22393_, _20849_, _05386_);
  or (_22394_, _22393_, _22339_);
  and (_22395_, _22394_, _03644_);
  or (_22396_, _22395_, _08861_);
  or (_22397_, _22396_, _22392_);
  and (_22398_, _13245_, _05386_);
  or (_22399_, _22339_, _04591_);
  or (_22400_, _22399_, _22398_);
  and (_22402_, _13363_, _05386_);
  or (_22403_, _22402_, _22339_);
  or (_22404_, _22403_, _04582_);
  and (_22405_, _22404_, _04589_);
  and (_22406_, _22405_, _22400_);
  and (_22407_, _22406_, _22397_);
  and (_22408_, _13374_, _05386_);
  or (_22409_, _22408_, _22339_);
  and (_22410_, _22409_, _03778_);
  or (_22411_, _22410_, _22407_);
  and (_22413_, _22411_, _04596_);
  or (_22414_, _22339_, _05491_);
  and (_22415_, _22403_, _03655_);
  and (_22416_, _22415_, _22414_);
  or (_22417_, _22416_, _22413_);
  and (_22418_, _22417_, _04594_);
  and (_22419_, _22344_, _03773_);
  and (_22420_, _22419_, _22414_);
  or (_22421_, _22420_, _03653_);
  or (_22422_, _22421_, _22418_);
  nor (_22425_, _13243_, _09486_);
  or (_22426_, _22339_, _04608_);
  or (_22427_, _22426_, _22425_);
  and (_22428_, _22427_, _04606_);
  and (_22429_, _22428_, _22422_);
  nor (_22430_, _13373_, _09486_);
  or (_22431_, _22430_, _22339_);
  and (_22432_, _22431_, _03786_);
  or (_22433_, _22432_, _03809_);
  or (_22434_, _22433_, _22429_);
  or (_22436_, _22341_, _04260_);
  and (_22437_, _22436_, _03206_);
  and (_22438_, _22437_, _22434_);
  and (_22439_, _22369_, _03205_);
  or (_22440_, _22439_, _03816_);
  or (_22441_, _22440_, _22438_);
  and (_22442_, _13425_, _05386_);
  or (_22443_, _22339_, _03820_);
  or (_22444_, _22443_, _22442_);
  and (_22445_, _22444_, _43227_);
  and (_22447_, _22445_, _22441_);
  or (_43500_, _22447_, _22338_);
  not (_22448_, \oc8051_golden_model_1.P3 [0]);
  nor (_22449_, _05388_, _22448_);
  and (_22450_, _12145_, _05388_);
  or (_22451_, _22450_, _22449_);
  and (_22452_, _22451_, _03778_);
  and (_22453_, _05388_, _04491_);
  or (_22454_, _22453_, _22449_);
  or (_22455_, _22454_, _06889_);
  nor (_22457_, _05744_, _09592_);
  or (_22458_, _22457_, _22449_);
  and (_22459_, _22458_, _03599_);
  nor (_22460_, _04499_, _22448_);
  and (_22461_, _05388_, \oc8051_golden_model_1.ACC [0]);
  or (_22462_, _22461_, _22449_);
  and (_22463_, _22462_, _04499_);
  or (_22464_, _22463_, _22460_);
  and (_22465_, _22464_, _04515_);
  or (_22466_, _22465_, _03515_);
  or (_22468_, _22466_, _22459_);
  and (_22469_, _12035_, _06016_);
  nor (_22470_, _06016_, _22448_);
  or (_22471_, _22470_, _03516_);
  or (_22472_, _22471_, _22469_);
  and (_22473_, _22472_, _04524_);
  and (_22474_, _22473_, _22468_);
  and (_22475_, _22454_, _03597_);
  or (_22476_, _22475_, _03603_);
  or (_22477_, _22476_, _22474_);
  or (_22479_, _22462_, _03611_);
  and (_22480_, _22479_, _03512_);
  and (_22481_, _22480_, _22477_);
  and (_22482_, _22449_, _03511_);
  or (_22483_, _22482_, _03504_);
  or (_22484_, _22483_, _22481_);
  or (_22485_, _22458_, _03505_);
  and (_22486_, _22485_, _03501_);
  and (_22487_, _22486_, _22484_);
  and (_22488_, _20078_, _06016_);
  or (_22490_, _22488_, _22470_);
  and (_22491_, _22490_, _03500_);
  or (_22492_, _22491_, _07441_);
  or (_22493_, _22492_, _22487_);
  and (_22494_, _22493_, _22455_);
  or (_22495_, _22494_, _05969_);
  and (_22496_, _06836_, _05388_);
  or (_22497_, _22449_, _05970_);
  or (_22498_, _22497_, _22496_);
  and (_22499_, _22498_, _03275_);
  and (_22501_, _22499_, _22495_);
  and (_22502_, _20114_, _05388_);
  or (_22503_, _22502_, _22449_);
  and (_22504_, _22503_, _03644_);
  or (_22505_, _22504_, _22501_);
  or (_22506_, _22505_, _08861_);
  and (_22507_, _12019_, _05388_);
  or (_22508_, _22449_, _04591_);
  or (_22509_, _22508_, _22507_);
  and (_22510_, _05388_, _06366_);
  or (_22512_, _22510_, _22449_);
  or (_22513_, _22512_, _04582_);
  and (_22514_, _22513_, _04589_);
  and (_22515_, _22514_, _22509_);
  and (_22516_, _22515_, _22506_);
  or (_22517_, _22516_, _22452_);
  and (_22518_, _22517_, _04596_);
  nand (_22519_, _22512_, _03655_);
  nor (_22520_, _22519_, _22457_);
  or (_22521_, _22520_, _22518_);
  and (_22523_, _22521_, _04594_);
  or (_22524_, _22449_, _05744_);
  and (_22525_, _22462_, _03773_);
  and (_22526_, _22525_, _22524_);
  or (_22527_, _22526_, _03653_);
  or (_22528_, _22527_, _22523_);
  nor (_22529_, _12017_, _09592_);
  or (_22530_, _22449_, _04608_);
  or (_22531_, _22530_, _22529_);
  and (_22532_, _22531_, _04606_);
  and (_22534_, _22532_, _22528_);
  nor (_22535_, _12015_, _09592_);
  or (_22536_, _22535_, _22449_);
  and (_22537_, _22536_, _03786_);
  or (_22538_, _22537_, _03809_);
  or (_22539_, _22538_, _22534_);
  or (_22540_, _22458_, _04260_);
  and (_22541_, _22540_, _03206_);
  and (_22542_, _22541_, _22539_);
  and (_22543_, _22449_, _03205_);
  or (_22545_, _22543_, _03816_);
  or (_22546_, _22545_, _22542_);
  or (_22547_, _22458_, _03820_);
  and (_22548_, _22547_, _43227_);
  and (_22549_, _22548_, _22546_);
  nor (_22550_, _43227_, _22448_);
  or (_22551_, _22550_, rst);
  or (_43503_, _22551_, _22549_);
  not (_22552_, \oc8051_golden_model_1.P3 [1]);
  nor (_22553_, _05388_, _22552_);
  and (_22555_, _05388_, _05898_);
  or (_22556_, _22555_, _22553_);
  or (_22557_, _22556_, _04524_);
  or (_22558_, _05388_, \oc8051_golden_model_1.P3 [1]);
  and (_22559_, _12234_, _05388_);
  not (_22560_, _22559_);
  and (_22561_, _22560_, _22558_);
  or (_22562_, _22561_, _04515_);
  nand (_22563_, _05388_, _03320_);
  and (_22564_, _22563_, _22558_);
  and (_22566_, _22564_, _04499_);
  nor (_22567_, _04499_, _22552_);
  or (_22568_, _22567_, _03599_);
  or (_22569_, _22568_, _22566_);
  and (_22570_, _22569_, _03516_);
  and (_22571_, _22570_, _22562_);
  nor (_22572_, _06016_, _22552_);
  and (_22573_, _12238_, _06016_);
  or (_22574_, _22573_, _22572_);
  and (_22575_, _22574_, _03515_);
  or (_22577_, _22575_, _03597_);
  or (_22578_, _22577_, _22571_);
  and (_22579_, _22578_, _22557_);
  or (_22580_, _22579_, _03603_);
  or (_22581_, _22564_, _03611_);
  and (_22582_, _22581_, _03512_);
  and (_22583_, _22582_, _22580_);
  and (_22584_, _12224_, _06016_);
  or (_22585_, _22584_, _22572_);
  and (_22586_, _22585_, _03511_);
  or (_22588_, _22586_, _03504_);
  or (_22589_, _22588_, _22583_);
  and (_22590_, _22573_, _12253_);
  or (_22591_, _22572_, _03505_);
  or (_22592_, _22591_, _22590_);
  and (_22593_, _22592_, _22589_);
  and (_22594_, _22593_, _03501_);
  and (_22595_, _20206_, _06016_);
  or (_22596_, _22572_, _22595_);
  and (_22597_, _22596_, _03500_);
  or (_22599_, _22597_, _07441_);
  or (_22600_, _22599_, _22594_);
  or (_22601_, _22556_, _06889_);
  and (_22602_, _22601_, _22600_);
  or (_22603_, _22602_, _05969_);
  and (_22604_, _06835_, _05388_);
  or (_22605_, _22553_, _05970_);
  or (_22606_, _22605_, _22604_);
  and (_22607_, _22606_, _03275_);
  and (_22608_, _22607_, _22603_);
  and (_22610_, _20235_, _05388_);
  or (_22611_, _22610_, _22553_);
  and (_22612_, _22611_, _03644_);
  or (_22613_, _22612_, _22608_);
  and (_22614_, _22613_, _03651_);
  or (_22615_, _12220_, _09592_);
  and (_22616_, _22615_, _03649_);
  nand (_22617_, _05388_, _04347_);
  and (_22618_, _22617_, _03650_);
  or (_22619_, _22618_, _22616_);
  and (_22621_, _22619_, _22558_);
  or (_22622_, _22621_, _22614_);
  and (_22623_, _22622_, _04589_);
  or (_22624_, _12347_, _09592_);
  and (_22625_, _22558_, _03778_);
  and (_22626_, _22625_, _22624_);
  or (_22627_, _22626_, _22623_);
  and (_22628_, _22627_, _04596_);
  or (_22629_, _12219_, _09592_);
  and (_22630_, _22558_, _03655_);
  and (_22632_, _22630_, _22629_);
  or (_22633_, _22632_, _22628_);
  and (_22634_, _22633_, _04594_);
  or (_22635_, _22553_, _05699_);
  and (_22636_, _22564_, _03773_);
  and (_22637_, _22636_, _22635_);
  or (_22638_, _22637_, _22634_);
  and (_22639_, _22638_, _03787_);
  or (_22640_, _22617_, _05699_);
  and (_22641_, _22558_, _03653_);
  and (_22643_, _22641_, _22640_);
  or (_22644_, _22563_, _05699_);
  and (_22645_, _22558_, _03786_);
  and (_22646_, _22645_, _22644_);
  or (_22647_, _22646_, _03809_);
  or (_22648_, _22647_, _22643_);
  or (_22649_, _22648_, _22639_);
  or (_22650_, _22561_, _04260_);
  and (_22651_, _22650_, _03206_);
  and (_22652_, _22651_, _22649_);
  and (_22654_, _22585_, _03205_);
  or (_22655_, _22654_, _03816_);
  or (_22656_, _22655_, _22652_);
  or (_22657_, _22553_, _03820_);
  or (_22658_, _22657_, _22559_);
  and (_22659_, _22658_, _43227_);
  and (_22660_, _22659_, _22656_);
  nor (_22661_, _43227_, _22552_);
  or (_22662_, _22661_, rst);
  or (_43504_, _22662_, _22660_);
  not (_22664_, \oc8051_golden_model_1.P3 [2]);
  nor (_22665_, _05388_, _22664_);
  nor (_22666_, _09592_, _05130_);
  or (_22667_, _22666_, _22665_);
  or (_22668_, _22667_, _06889_);
  and (_22669_, _22667_, _03597_);
  nor (_22670_, _06016_, _22664_);
  and (_22671_, _12416_, _06016_);
  or (_22672_, _22671_, _22670_);
  or (_22673_, _22672_, _03516_);
  nor (_22675_, _12430_, _09592_);
  or (_22676_, _22675_, _22665_);
  and (_22677_, _22676_, _03599_);
  nor (_22678_, _04499_, _22664_);
  and (_22679_, _05388_, \oc8051_golden_model_1.ACC [2]);
  or (_22680_, _22679_, _22665_);
  and (_22681_, _22680_, _04499_);
  or (_22682_, _22681_, _22678_);
  and (_22683_, _22682_, _04515_);
  or (_22684_, _22683_, _03515_);
  or (_22686_, _22684_, _22677_);
  and (_22687_, _22686_, _22673_);
  and (_22688_, _22687_, _04524_);
  or (_22689_, _22688_, _22669_);
  or (_22690_, _22689_, _03603_);
  or (_22691_, _22680_, _03611_);
  and (_22692_, _22691_, _03512_);
  and (_22693_, _22692_, _22690_);
  and (_22694_, _12414_, _06016_);
  or (_22695_, _22694_, _22670_);
  and (_22697_, _22695_, _03511_);
  or (_22698_, _22697_, _03504_);
  or (_22699_, _22698_, _22693_);
  or (_22700_, _22670_, _12447_);
  and (_22701_, _22700_, _22672_);
  or (_22702_, _22701_, _03505_);
  and (_22703_, _22702_, _03501_);
  and (_22704_, _22703_, _22699_);
  and (_22705_, _20332_, _06016_);
  or (_22706_, _22705_, _22670_);
  and (_22708_, _22706_, _03500_);
  or (_22709_, _22708_, _07441_);
  or (_22710_, _22709_, _22704_);
  and (_22711_, _22710_, _22668_);
  or (_22712_, _22711_, _05969_);
  and (_22713_, _06839_, _05388_);
  or (_22714_, _22665_, _05970_);
  or (_22715_, _22714_, _22713_);
  and (_22716_, _22715_, _03275_);
  and (_22717_, _22716_, _22712_);
  and (_22719_, _20358_, _05388_);
  or (_22720_, _22665_, _22719_);
  and (_22721_, _22720_, _03644_);
  or (_22722_, _22721_, _22717_);
  or (_22723_, _22722_, _08861_);
  and (_22724_, _12538_, _05388_);
  or (_22725_, _22665_, _04591_);
  or (_22726_, _22725_, _22724_);
  and (_22727_, _05388_, _06414_);
  or (_22728_, _22727_, _22665_);
  or (_22730_, _22728_, _04582_);
  and (_22731_, _22730_, _04589_);
  and (_22732_, _22731_, _22726_);
  and (_22733_, _22732_, _22723_);
  and (_22734_, _12544_, _05388_);
  or (_22735_, _22734_, _22665_);
  and (_22736_, _22735_, _03778_);
  or (_22737_, _22736_, _22733_);
  and (_22738_, _22737_, _04596_);
  or (_22739_, _22665_, _05793_);
  and (_22741_, _22728_, _03655_);
  and (_22742_, _22741_, _22739_);
  or (_22743_, _22742_, _22738_);
  and (_22744_, _22743_, _04594_);
  and (_22745_, _22680_, _03773_);
  and (_22746_, _22745_, _22739_);
  or (_22747_, _22746_, _03653_);
  or (_22748_, _22747_, _22744_);
  nor (_22749_, _12537_, _09592_);
  or (_22750_, _22665_, _04608_);
  or (_22752_, _22750_, _22749_);
  and (_22753_, _22752_, _04606_);
  and (_22754_, _22753_, _22748_);
  nor (_22755_, _12543_, _09592_);
  or (_22756_, _22755_, _22665_);
  and (_22757_, _22756_, _03786_);
  or (_22758_, _22757_, _03809_);
  or (_22759_, _22758_, _22754_);
  or (_22760_, _22676_, _04260_);
  and (_22761_, _22760_, _03206_);
  and (_22763_, _22761_, _22759_);
  and (_22764_, _22695_, _03205_);
  or (_22765_, _22764_, _03816_);
  or (_22766_, _22765_, _22763_);
  and (_22767_, _12600_, _05388_);
  or (_22768_, _22665_, _03820_);
  or (_22769_, _22768_, _22767_);
  and (_22770_, _22769_, _43227_);
  and (_22771_, _22770_, _22766_);
  nor (_22772_, _43227_, _22664_);
  or (_22774_, _22772_, rst);
  or (_43505_, _22774_, _22771_);
  and (_22775_, _09592_, \oc8051_golden_model_1.P3 [3]);
  nor (_22776_, _09592_, _04944_);
  or (_22777_, _22776_, _22775_);
  or (_22778_, _22777_, _06889_);
  nor (_22779_, _12625_, _09592_);
  or (_22780_, _22779_, _22775_);
  or (_22781_, _22780_, _04515_);
  and (_22782_, _05388_, \oc8051_golden_model_1.ACC [3]);
  or (_22784_, _22782_, _22775_);
  and (_22785_, _22784_, _04499_);
  and (_22786_, _04500_, \oc8051_golden_model_1.P3 [3]);
  or (_22787_, _22786_, _03599_);
  or (_22788_, _22787_, _22785_);
  and (_22789_, _22788_, _03516_);
  and (_22790_, _22789_, _22781_);
  not (_22791_, _06016_);
  and (_22792_, _22791_, \oc8051_golden_model_1.P3 [3]);
  and (_22793_, _12638_, _06016_);
  or (_22795_, _22793_, _22792_);
  and (_22796_, _22795_, _03515_);
  or (_22797_, _22796_, _03597_);
  or (_22798_, _22797_, _22790_);
  or (_22799_, _22777_, _04524_);
  and (_22800_, _22799_, _22798_);
  or (_22801_, _22800_, _03603_);
  or (_22802_, _22784_, _03611_);
  and (_22803_, _22802_, _03512_);
  and (_22804_, _22803_, _22801_);
  and (_22806_, _12622_, _06016_);
  or (_22807_, _22806_, _22792_);
  and (_22808_, _22807_, _03511_);
  or (_22809_, _22808_, _03504_);
  or (_22810_, _22809_, _22804_);
  or (_22811_, _22792_, _12653_);
  and (_22812_, _22811_, _22795_);
  or (_22813_, _22812_, _03505_);
  and (_22814_, _22813_, _03501_);
  and (_22815_, _22814_, _22810_);
  and (_22817_, _20458_, _06016_);
  or (_22818_, _22817_, _22792_);
  and (_22819_, _22818_, _03500_);
  or (_22820_, _22819_, _07441_);
  or (_22821_, _22820_, _22815_);
  and (_22822_, _22821_, _22778_);
  or (_22823_, _22822_, _05969_);
  and (_22824_, _06838_, _05388_);
  or (_22825_, _22775_, _05970_);
  or (_22826_, _22825_, _22824_);
  and (_22828_, _22826_, _03275_);
  and (_22829_, _22828_, _22823_);
  and (_22830_, _20485_, _05388_);
  or (_22831_, _22775_, _22830_);
  and (_22832_, _22831_, _03644_);
  or (_22833_, _22832_, _22829_);
  or (_22834_, _22833_, _08861_);
  and (_22835_, _12746_, _05388_);
  or (_22836_, _22775_, _04591_);
  or (_22837_, _22836_, _22835_);
  and (_22839_, _05388_, _06347_);
  or (_22840_, _22839_, _22775_);
  or (_22841_, _22840_, _04582_);
  and (_22842_, _22841_, _04589_);
  and (_22843_, _22842_, _22837_);
  and (_22844_, _22843_, _22834_);
  and (_22845_, _12619_, _05388_);
  or (_22846_, _22845_, _22775_);
  and (_22847_, _22846_, _03778_);
  or (_22848_, _22847_, _22844_);
  and (_22850_, _22848_, _04596_);
  or (_22851_, _22775_, _05650_);
  and (_22852_, _22840_, _03655_);
  and (_22853_, _22852_, _22851_);
  or (_22854_, _22853_, _22850_);
  and (_22855_, _22854_, _04594_);
  and (_22856_, _22784_, _03773_);
  and (_22857_, _22856_, _22851_);
  or (_22858_, _22857_, _03653_);
  or (_22859_, _22858_, _22855_);
  nor (_22861_, _12745_, _09592_);
  or (_22862_, _22775_, _04608_);
  or (_22863_, _22862_, _22861_);
  and (_22864_, _22863_, _04606_);
  and (_22865_, _22864_, _22859_);
  nor (_22866_, _12618_, _09592_);
  or (_22867_, _22866_, _22775_);
  and (_22868_, _22867_, _03786_);
  or (_22869_, _22868_, _03809_);
  or (_22870_, _22869_, _22865_);
  or (_22872_, _22780_, _04260_);
  and (_22873_, _22872_, _03206_);
  and (_22874_, _22873_, _22870_);
  and (_22875_, _22807_, _03205_);
  or (_22876_, _22875_, _03816_);
  or (_22877_, _22876_, _22874_);
  and (_22878_, _12806_, _05388_);
  or (_22879_, _22775_, _03820_);
  or (_22880_, _22879_, _22878_);
  and (_22881_, _22880_, _43227_);
  and (_22883_, _22881_, _22877_);
  nor (_22884_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_22885_, _22884_, _05217_);
  or (_43506_, _22885_, _22883_);
  and (_22886_, _09592_, \oc8051_golden_model_1.P3 [4]);
  nor (_22887_, _05840_, _09592_);
  or (_22888_, _22887_, _22886_);
  or (_22889_, _22888_, _06889_);
  and (_22890_, _22791_, \oc8051_golden_model_1.P3 [4]);
  and (_22891_, _12853_, _06016_);
  or (_22893_, _22891_, _22890_);
  and (_22894_, _22893_, _03511_);
  nor (_22895_, _12820_, _09592_);
  or (_22896_, _22895_, _22886_);
  or (_22897_, _22896_, _04515_);
  and (_22898_, _05388_, \oc8051_golden_model_1.ACC [4]);
  or (_22899_, _22898_, _22886_);
  and (_22900_, _22899_, _04499_);
  and (_22901_, _04500_, \oc8051_golden_model_1.P3 [4]);
  or (_22902_, _22901_, _03599_);
  or (_22904_, _22902_, _22900_);
  and (_22905_, _22904_, _03516_);
  and (_22906_, _22905_, _22897_);
  and (_22907_, _12830_, _06016_);
  or (_22908_, _22907_, _22890_);
  and (_22909_, _22908_, _03515_);
  or (_22910_, _22909_, _03597_);
  or (_22911_, _22910_, _22906_);
  or (_22912_, _22888_, _04524_);
  and (_22913_, _22912_, _22911_);
  or (_22915_, _22913_, _03603_);
  or (_22916_, _22899_, _03611_);
  and (_22917_, _22916_, _03512_);
  and (_22918_, _22917_, _22915_);
  or (_22919_, _22918_, _22894_);
  and (_22920_, _22919_, _03505_);
  or (_22921_, _22890_, _12860_);
  and (_22922_, _22921_, _03504_);
  and (_22923_, _22922_, _22908_);
  or (_22924_, _22923_, _22920_);
  and (_22926_, _22924_, _03501_);
  and (_22927_, _20579_, _06016_);
  or (_22928_, _22927_, _22890_);
  and (_22929_, _22928_, _03500_);
  or (_22930_, _22929_, _07441_);
  or (_22931_, _22930_, _22926_);
  and (_22932_, _22931_, _22889_);
  or (_22933_, _22932_, _05969_);
  and (_22934_, _06843_, _05388_);
  or (_22935_, _22886_, _05970_);
  or (_22937_, _22935_, _22934_);
  and (_22938_, _22937_, _03275_);
  and (_22939_, _22938_, _22933_);
  and (_22940_, _20605_, _05388_);
  or (_22941_, _22940_, _22886_);
  and (_22942_, _22941_, _03644_);
  or (_22943_, _22942_, _08861_);
  or (_22944_, _22943_, _22939_);
  and (_22945_, _12951_, _05388_);
  or (_22946_, _22886_, _04591_);
  or (_22948_, _22946_, _22945_);
  and (_22949_, _06375_, _05388_);
  or (_22950_, _22949_, _22886_);
  or (_22951_, _22950_, _04582_);
  and (_22952_, _22951_, _04589_);
  and (_22953_, _22952_, _22948_);
  and (_22954_, _22953_, _22944_);
  and (_22955_, _12957_, _05388_);
  or (_22956_, _22955_, _22886_);
  and (_22957_, _22956_, _03778_);
  or (_22959_, _22957_, _22954_);
  and (_22960_, _22959_, _04596_);
  or (_22961_, _22886_, _05889_);
  and (_22962_, _22950_, _03655_);
  and (_22963_, _22962_, _22961_);
  or (_22964_, _22963_, _22960_);
  and (_22965_, _22964_, _04594_);
  and (_22966_, _22899_, _03773_);
  and (_22967_, _22966_, _22961_);
  or (_22968_, _22967_, _03653_);
  or (_22970_, _22968_, _22965_);
  nor (_22971_, _12949_, _09592_);
  or (_22972_, _22886_, _04608_);
  or (_22973_, _22972_, _22971_);
  and (_22974_, _22973_, _04606_);
  and (_22975_, _22974_, _22970_);
  nor (_22976_, _12956_, _09592_);
  or (_22977_, _22976_, _22886_);
  and (_22978_, _22977_, _03786_);
  or (_22979_, _22978_, _03809_);
  or (_22980_, _22979_, _22975_);
  or (_22981_, _22896_, _04260_);
  and (_22982_, _22981_, _03206_);
  and (_22983_, _22982_, _22980_);
  and (_22984_, _22893_, _03205_);
  or (_22985_, _22984_, _03816_);
  or (_22986_, _22985_, _22983_);
  and (_22987_, _13013_, _05388_);
  or (_22988_, _22886_, _03820_);
  or (_22989_, _22988_, _22987_);
  and (_22992_, _22989_, _43227_);
  and (_22993_, _22992_, _22986_);
  nor (_22994_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_22995_, _22994_, _05217_);
  or (_43507_, _22995_, _22993_);
  nor (_22996_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_22997_, _22996_, _05217_);
  and (_22998_, _09592_, \oc8051_golden_model_1.P3 [5]);
  nor (_22999_, _13035_, _09592_);
  or (_23000_, _22999_, _22998_);
  or (_23002_, _23000_, _04515_);
  and (_23003_, _05388_, \oc8051_golden_model_1.ACC [5]);
  or (_23004_, _23003_, _22998_);
  and (_23005_, _23004_, _04499_);
  and (_23006_, _04500_, \oc8051_golden_model_1.P3 [5]);
  or (_23007_, _23006_, _03599_);
  or (_23008_, _23007_, _23005_);
  and (_23009_, _23008_, _03516_);
  and (_23010_, _23009_, _23002_);
  and (_23011_, _22791_, \oc8051_golden_model_1.P3 [5]);
  and (_23012_, _13051_, _06016_);
  or (_23013_, _23012_, _23011_);
  and (_23014_, _23013_, _03515_);
  or (_23015_, _23014_, _03597_);
  or (_23016_, _23015_, _23010_);
  nor (_23017_, _05552_, _09592_);
  or (_23018_, _23017_, _22998_);
  or (_23019_, _23018_, _04524_);
  and (_23020_, _23019_, _23016_);
  or (_23021_, _23020_, _03603_);
  or (_23024_, _23004_, _03611_);
  and (_23025_, _23024_, _03512_);
  and (_23026_, _23025_, _23021_);
  and (_23027_, _13032_, _06016_);
  or (_23028_, _23027_, _23011_);
  and (_23029_, _23028_, _03511_);
  or (_23030_, _23029_, _03504_);
  or (_23031_, _23030_, _23026_);
  or (_23032_, _23011_, _13066_);
  and (_23033_, _23032_, _23013_);
  or (_23035_, _23033_, _03505_);
  and (_23036_, _23035_, _03501_);
  and (_23037_, _23036_, _23031_);
  and (_23038_, _20702_, _06016_);
  or (_23039_, _23038_, _23011_);
  and (_23040_, _23039_, _03500_);
  or (_23041_, _23040_, _07441_);
  or (_23042_, _23041_, _23037_);
  or (_23043_, _23018_, _06889_);
  and (_23044_, _23043_, _23042_);
  or (_23045_, _23044_, _05969_);
  and (_23046_, _06842_, _05388_);
  or (_23047_, _22998_, _05970_);
  or (_23048_, _23047_, _23046_);
  and (_23049_, _23048_, _03275_);
  and (_23050_, _23049_, _23045_);
  and (_23051_, _20729_, _05388_);
  or (_23052_, _23051_, _22998_);
  and (_23053_, _23052_, _03644_);
  or (_23054_, _23053_, _08861_);
  or (_23057_, _23054_, _23050_);
  and (_23058_, _13154_, _05388_);
  or (_23059_, _22998_, _04591_);
  or (_23060_, _23059_, _23058_);
  and (_23061_, _06358_, _05388_);
  or (_23062_, _23061_, _22998_);
  or (_23063_, _23062_, _04582_);
  and (_23064_, _23063_, _04589_);
  and (_23065_, _23064_, _23060_);
  and (_23066_, _23065_, _23057_);
  and (_23068_, _13160_, _05388_);
  or (_23069_, _23068_, _22998_);
  and (_23070_, _23069_, _03778_);
  or (_23071_, _23070_, _23066_);
  and (_23072_, _23071_, _04596_);
  or (_23073_, _22998_, _05601_);
  and (_23074_, _23062_, _03655_);
  and (_23075_, _23074_, _23073_);
  or (_23076_, _23075_, _23072_);
  and (_23077_, _23076_, _04594_);
  and (_23078_, _23004_, _03773_);
  and (_23079_, _23078_, _23073_);
  or (_23080_, _23079_, _03653_);
  or (_23081_, _23080_, _23077_);
  nor (_23082_, _13152_, _09592_);
  or (_23083_, _22998_, _04608_);
  or (_23084_, _23083_, _23082_);
  and (_23085_, _23084_, _04606_);
  and (_23086_, _23085_, _23081_);
  nor (_23087_, _13159_, _09592_);
  or (_23090_, _23087_, _22998_);
  and (_23091_, _23090_, _03786_);
  or (_23092_, _23091_, _03809_);
  or (_23093_, _23092_, _23086_);
  or (_23094_, _23000_, _04260_);
  and (_23095_, _23094_, _03206_);
  and (_23096_, _23095_, _23093_);
  and (_23097_, _23028_, _03205_);
  or (_23098_, _23097_, _03816_);
  or (_23099_, _23098_, _23096_);
  and (_23101_, _13217_, _05388_);
  or (_23102_, _22998_, _03820_);
  or (_23103_, _23102_, _23101_);
  and (_23104_, _23103_, _43227_);
  and (_23105_, _23104_, _23099_);
  or (_43508_, _23105_, _22997_);
  not (_23106_, \oc8051_golden_model_1.P3 [6]);
  nor (_23107_, _05388_, _23106_);
  nor (_23108_, _13235_, _09592_);
  or (_23109_, _23108_, _23107_);
  or (_23110_, _23109_, _04515_);
  and (_23111_, _05388_, \oc8051_golden_model_1.ACC [6]);
  or (_23112_, _23111_, _23107_);
  and (_23113_, _23112_, _04499_);
  nor (_23114_, _04499_, _23106_);
  or (_23115_, _23114_, _03599_);
  or (_23116_, _23115_, _23113_);
  and (_23117_, _23116_, _03516_);
  and (_23118_, _23117_, _23110_);
  nor (_23119_, _06016_, _23106_);
  and (_23122_, _13266_, _06016_);
  or (_23123_, _23122_, _23119_);
  and (_23124_, _23123_, _03515_);
  or (_23125_, _23124_, _03597_);
  or (_23126_, _23125_, _23118_);
  nor (_23127_, _05442_, _09592_);
  or (_23128_, _23127_, _23107_);
  or (_23129_, _23128_, _04524_);
  and (_23130_, _23129_, _23126_);
  or (_23131_, _23130_, _03603_);
  or (_23133_, _23112_, _03611_);
  and (_23134_, _23133_, _03512_);
  and (_23135_, _23134_, _23131_);
  and (_23136_, _13251_, _06016_);
  or (_23137_, _23136_, _23119_);
  and (_23138_, _23137_, _03511_);
  or (_23139_, _23138_, _03504_);
  or (_23140_, _23139_, _23135_);
  or (_23141_, _23119_, _13281_);
  and (_23142_, _23141_, _23123_);
  or (_23143_, _23142_, _03505_);
  and (_23144_, _23143_, _03501_);
  and (_23145_, _23144_, _23140_);
  and (_23146_, _20822_, _06016_);
  or (_23147_, _23146_, _23119_);
  and (_23148_, _23147_, _03500_);
  or (_23149_, _23148_, _07441_);
  or (_23150_, _23149_, _23145_);
  or (_23151_, _23128_, _06889_);
  and (_23152_, _23151_, _23150_);
  or (_23155_, _23152_, _05969_);
  and (_23156_, _06531_, _05388_);
  or (_23157_, _23107_, _05970_);
  or (_23158_, _23157_, _23156_);
  and (_23159_, _23158_, _03275_);
  and (_23160_, _23159_, _23155_);
  and (_23161_, _20849_, _05388_);
  or (_23162_, _23161_, _23107_);
  and (_23163_, _23162_, _03644_);
  or (_23164_, _23163_, _08861_);
  or (_23166_, _23164_, _23160_);
  and (_23167_, _13245_, _05388_);
  or (_23168_, _23107_, _04591_);
  or (_23169_, _23168_, _23167_);
  and (_23170_, _13363_, _05388_);
  or (_23171_, _23170_, _23107_);
  or (_23172_, _23171_, _04582_);
  and (_23173_, _23172_, _04589_);
  and (_23174_, _23173_, _23169_);
  and (_23175_, _23174_, _23166_);
  and (_23176_, _13374_, _05388_);
  or (_23177_, _23176_, _23107_);
  and (_23178_, _23177_, _03778_);
  or (_23179_, _23178_, _23175_);
  and (_23180_, _23179_, _04596_);
  or (_23181_, _23107_, _05491_);
  and (_23182_, _23171_, _03655_);
  and (_23183_, _23182_, _23181_);
  or (_23184_, _23183_, _23180_);
  and (_23185_, _23184_, _04594_);
  and (_23188_, _23112_, _03773_);
  and (_23189_, _23188_, _23181_);
  or (_23190_, _23189_, _03653_);
  or (_23191_, _23190_, _23185_);
  nor (_23192_, _13243_, _09592_);
  or (_23193_, _23107_, _04608_);
  or (_23194_, _23193_, _23192_);
  and (_23195_, _23194_, _04606_);
  and (_23196_, _23195_, _23191_);
  nor (_23197_, _13373_, _09592_);
  or (_23199_, _23197_, _23107_);
  and (_23200_, _23199_, _03786_);
  or (_23201_, _23200_, _03809_);
  or (_23202_, _23201_, _23196_);
  or (_23203_, _23109_, _04260_);
  and (_23204_, _23203_, _03206_);
  and (_23205_, _23204_, _23202_);
  and (_23206_, _23137_, _03205_);
  or (_23207_, _23206_, _03816_);
  or (_23208_, _23207_, _23205_);
  and (_23210_, _13425_, _05388_);
  or (_23211_, _23107_, _03820_);
  or (_23212_, _23211_, _23210_);
  and (_23213_, _23212_, _43227_);
  and (_23214_, _23213_, _23208_);
  nor (_23215_, _43227_, _23106_);
  or (_23216_, _23215_, rst);
  or (_43509_, _23216_, _23214_);
  not (_23217_, \oc8051_golden_model_1.PSW [0]);
  nor (_23218_, _43227_, _23217_);
  nor (_23220_, _07578_, _07577_);
  nor (_23221_, _23220_, _07484_);
  and (_23222_, _23220_, _07484_);
  nor (_23223_, _23222_, _23221_);
  nor (_23224_, _07501_, _07500_);
  nor (_23225_, _23224_, _15488_);
  and (_23226_, _23224_, _15488_);
  nor (_23227_, _23226_, _23225_);
  and (_23228_, _23227_, _23223_);
  nor (_23229_, _23227_, _23223_);
  nor (_23231_, _23229_, _23228_);
  or (_23232_, _23231_, _06061_);
  nand (_23233_, _23231_, _06061_);
  and (_23234_, _23233_, _23232_);
  or (_23235_, _23234_, _05913_);
  nor (_23236_, _15122_, _08659_);
  and (_23237_, _15122_, _08659_);
  nor (_23238_, _23237_, _23236_);
  and (_23239_, _23238_, _15777_);
  nor (_23240_, _23238_, _15777_);
  nor (_23242_, _23240_, _23239_);
  and (_23243_, _23242_, _15837_);
  nor (_23244_, _23242_, _15837_);
  nor (_23245_, _23244_, _23243_);
  and (_23246_, _23245_, _16430_);
  nor (_23247_, _23245_, _16430_);
  nor (_23248_, _23247_, _23246_);
  nor (_23249_, _23248_, _16748_);
  and (_23250_, _23248_, _16748_);
  nor (_23251_, _23250_, _23249_);
  and (_23253_, _23251_, _17089_);
  nor (_23254_, _23251_, _17089_);
  or (_23255_, _23254_, _23253_);
  nor (_23256_, _23255_, _08675_);
  and (_23257_, _23255_, _08675_);
  or (_23258_, _23257_, _23256_);
  or (_23259_, _23258_, _08639_);
  or (_23260_, _08660_, _08657_);
  nand (_23261_, _08660_, _08657_);
  and (_23262_, _23261_, _23260_);
  nor (_23264_, _08652_, _08653_);
  and (_23265_, _08652_, _08653_);
  nor (_23266_, _23265_, _23264_);
  and (_23267_, _23266_, _23262_);
  nor (_23268_, _23266_, _23262_);
  nor (_23269_, _23268_, _23267_);
  not (_23270_, _08644_);
  nor (_23271_, _08646_, _08641_);
  and (_23272_, _08646_, _08641_);
  nor (_23273_, _23272_, _23271_);
  nor (_23275_, _23273_, _23270_);
  and (_23276_, _23273_, _23270_);
  nor (_23277_, _23276_, _23275_);
  and (_23278_, _23277_, _23269_);
  nor (_23279_, _23277_, _23269_);
  or (_23280_, _23279_, _23278_);
  and (_23281_, _23280_, _07946_);
  nor (_23282_, _23280_, _07946_);
  or (_23283_, _23282_, _23281_);
  or (_23284_, _23283_, _07945_);
  and (_23286_, _11374_, _11373_);
  not (_23287_, _23286_);
  nor (_23288_, _23287_, _05965_);
  or (_23289_, _23288_, _23234_);
  and (_23290_, _03582_, _03503_);
  not (_23291_, _23290_);
  and (_23292_, _11697_, _23291_);
  and (_23293_, _23292_, _03672_);
  or (_23294_, _23293_, _23234_);
  or (_23295_, _06840_, _06715_);
  nand (_23297_, _23295_, _12393_);
  or (_23298_, _23295_, _12393_);
  and (_23299_, _23298_, _23297_);
  or (_23300_, _06844_, _06807_);
  nand (_23301_, _23300_, _06531_);
  or (_23302_, _23300_, _06531_);
  and (_23303_, _23302_, _23301_);
  and (_23304_, _23303_, _23299_);
  nor (_23305_, _23303_, _23299_);
  or (_23306_, _23305_, _23304_);
  nor (_23308_, _23306_, _06171_);
  and (_23309_, _23306_, _06171_);
  or (_23310_, _23309_, _23308_);
  or (_23311_, _23310_, _08052_);
  and (_23312_, _06054_, _03262_);
  nor (_23313_, _06046_, _05900_);
  nor (_23314_, _06044_, _05902_);
  not (_23315_, _23314_);
  and (_23316_, _23315_, _23313_);
  nor (_23317_, _23315_, _23313_);
  nor (_23318_, _23317_, _23316_);
  nor (_23319_, _12214_, _05907_);
  and (_23320_, _12214_, _05907_);
  nor (_23321_, _23320_, _23319_);
  nor (_23322_, _23321_, _23318_);
  and (_23323_, _23321_, _23318_);
  or (_23324_, _23323_, _23322_);
  or (_23325_, _23324_, _08048_);
  and (_23326_, _11531_, _03948_);
  nand (_23327_, _23326_, _23217_);
  or (_23329_, _23326_, _23234_);
  and (_23330_, _23329_, _23327_);
  or (_23331_, _23330_, _08049_);
  and (_23332_, _23331_, _23325_);
  or (_23333_, _23332_, _08051_);
  and (_23334_, _23333_, _23312_);
  and (_23335_, _23334_, _23311_);
  and (_23336_, _23234_, _12226_);
  or (_23337_, _23336_, _04509_);
  or (_23338_, _23337_, _23335_);
  nor (_23340_, _23224_, \oc8051_golden_model_1.ACC [6]);
  and (_23341_, _23224_, \oc8051_golden_model_1.ACC [6]);
  nor (_23342_, _23341_, _23340_);
  nor (_23343_, _23342_, \oc8051_golden_model_1.ACC [7]);
  and (_23344_, _23342_, \oc8051_golden_model_1.ACC [7]);
  nor (_23345_, _23344_, _23343_);
  nor (_23346_, _23345_, _23299_);
  and (_23347_, _23345_, _23299_);
  or (_23348_, _23347_, _23346_);
  or (_23349_, _23348_, _06068_);
  and (_23350_, _23349_, _04515_);
  and (_23351_, _23350_, _23338_);
  not (_23352_, _16857_);
  not (_23353_, _15044_);
  nor (_23354_, _15273_, _23353_);
  and (_23355_, _15273_, _23353_);
  nor (_23356_, _23355_, _23354_);
  and (_23357_, _23356_, _15539_);
  nor (_23358_, _23356_, _15539_);
  nor (_23359_, _23358_, _23357_);
  and (_23360_, _23359_, _16542_);
  nor (_23361_, _23359_, _16542_);
  or (_23362_, _23361_, _23360_);
  nor (_23363_, _16217_, _15888_);
  and (_23364_, _16217_, _15888_);
  nor (_23365_, _23364_, _23363_);
  and (_23366_, _23365_, _23362_);
  nor (_23367_, _23365_, _23362_);
  nor (_23368_, _23367_, _23366_);
  nor (_23369_, _23368_, _23352_);
  and (_23370_, _23368_, _23352_);
  or (_23371_, _23370_, _23369_);
  and (_23372_, _23371_, _08065_);
  nor (_23373_, _23371_, _08065_);
  or (_23374_, _23373_, _23372_);
  and (_23375_, _23374_, _03599_);
  or (_23376_, _23375_, _08063_);
  or (_23377_, _23376_, _23351_);
  and (_23378_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_23379_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_23380_, _23379_, _23378_);
  and (_23381_, _23380_, _15279_);
  nor (_23382_, _23380_, _15279_);
  nor (_23383_, _23382_, _23381_);
  nor (_23384_, _15894_, _07536_);
  and (_23385_, _15894_, _07536_);
  nor (_23386_, _23385_, _23384_);
  and (_23387_, _23386_, _23383_);
  nor (_23388_, _23386_, _23383_);
  nor (_23389_, _23388_, _23387_);
  nor (_23390_, _23389_, _16550_);
  and (_23391_, _23389_, _16550_);
  nor (_23392_, _23391_, _23390_);
  not (_23393_, _23392_);
  nor (_23394_, _16876_, _08088_);
  and (_23395_, _16876_, _08088_);
  nor (_23396_, _23395_, _23394_);
  nor (_23397_, _23396_, _23393_);
  and (_23398_, _23396_, _23393_);
  or (_23399_, _23398_, _23397_);
  or (_23401_, _23399_, _09952_);
  and (_23402_, _23401_, _23377_);
  or (_23403_, _23402_, _09965_);
  or (_23404_, _23234_, _09966_);
  and (_23405_, _23404_, _03516_);
  and (_23406_, _23405_, _23403_);
  not (_23407_, _08094_);
  and (_23408_, _15286_, _15050_);
  nor (_23409_, _15286_, _15050_);
  or (_23410_, _23409_, _23408_);
  nor (_23412_, _16882_, _16229_);
  and (_23413_, _16882_, _16229_);
  nor (_23414_, _23413_, _23412_);
  nor (_23415_, _23414_, _23410_);
  and (_23416_, _23414_, _23410_);
  or (_23417_, _23416_, _23415_);
  not (_23418_, _16554_);
  nor (_23419_, _15900_, _15553_);
  and (_23420_, _15900_, _15553_);
  nor (_23421_, _23420_, _23419_);
  nor (_23422_, _23421_, _23418_);
  and (_23423_, _23421_, _23418_);
  nor (_23424_, _23423_, _23422_);
  and (_23425_, _23424_, _23417_);
  nor (_23426_, _23424_, _23417_);
  nor (_23427_, _23426_, _23425_);
  nand (_23428_, _23427_, _23407_);
  or (_23429_, _23427_, _23407_);
  and (_23430_, _23429_, _03515_);
  and (_23431_, _23430_, _23428_);
  or (_23433_, _23431_, _04857_);
  or (_23434_, _23433_, _23406_);
  or (_23435_, _23234_, _03257_);
  and (_23436_, _23435_, _23434_);
  or (_23437_, _23436_, _03597_);
  not (_23438_, _16826_);
  and (_23439_, _23438_, _07959_);
  nor (_23440_, _23438_, _07959_);
  nor (_23441_, _23440_, _23439_);
  and (_23442_, _15249_, _15026_);
  nor (_23444_, _15249_, _15026_);
  nor (_23445_, _23444_, _23442_);
  not (_23446_, _15851_);
  and (_23447_, _23446_, _15523_);
  nor (_23448_, _23446_, _15523_);
  nor (_23449_, _23448_, _23447_);
  nor (_23450_, _23449_, _23445_);
  and (_23451_, _23449_, _23445_);
  or (_23452_, _23451_, _23450_);
  not (_23453_, _16503_);
  and (_23455_, _23453_, _16173_);
  nor (_23456_, _23453_, _16173_);
  nor (_23457_, _23456_, _23455_);
  and (_23458_, _23457_, _23452_);
  nor (_23459_, _23457_, _23452_);
  nor (_23460_, _23459_, _23458_);
  or (_23461_, _23460_, _23441_);
  nand (_23462_, _23460_, _23441_);
  and (_23463_, _23462_, _23461_);
  or (_23464_, _23463_, _04524_);
  and (_23466_, _23464_, _08040_);
  and (_23467_, _23466_, _23437_);
  not (_23468_, _08040_);
  and (_23469_, _23324_, _23468_);
  or (_23470_, _23469_, _23467_);
  and (_23471_, _23470_, _08039_);
  and (_23472_, _23324_, _04848_);
  or (_23473_, _23472_, _04529_);
  or (_23474_, _23473_, _23471_);
  or (_23475_, _23310_, _08102_);
  and (_23476_, _23475_, _03611_);
  and (_23477_, _23476_, _23474_);
  not (_23478_, _08238_);
  nor (_23479_, _08223_, _08208_);
  and (_23480_, _08223_, _08208_);
  nor (_23481_, _23480_, _23479_);
  nor (_23482_, _23481_, _23478_);
  and (_23483_, _23481_, _23478_);
  nor (_23484_, _23483_, _23482_);
  and (_23485_, _08269_, _08255_);
  nor (_23487_, _23485_, _08270_);
  and (_23488_, _08191_, _08173_);
  nor (_23489_, _08191_, _08173_);
  or (_23490_, _23489_, _23488_);
  and (_23491_, _23490_, _23487_);
  nor (_23492_, _23490_, _23487_);
  nor (_23493_, _23492_, _23491_);
  nor (_23494_, _23493_, _23484_);
  and (_23495_, _23493_, _23484_);
  nor (_23496_, _23495_, _23494_);
  or (_23498_, _23496_, _06211_);
  nand (_23499_, _23496_, _06211_);
  and (_23500_, _23499_, _03603_);
  and (_23501_, _23500_, _23498_);
  or (_23502_, _23501_, _11694_);
  or (_23503_, _23502_, _23477_);
  or (_23504_, _23234_, _11692_);
  and (_23505_, _23504_, _03512_);
  and (_23506_, _23505_, _23503_);
  nor (_23507_, _15305_, _15011_);
  and (_23509_, _15305_, _15011_);
  nor (_23510_, _23509_, _23507_);
  nor (_23511_, _16903_, _08114_);
  and (_23512_, _16903_, _08114_);
  nor (_23513_, _23512_, _23511_);
  nor (_23514_, _23513_, _23510_);
  and (_23515_, _23513_, _23510_);
  nor (_23516_, _23515_, _23514_);
  not (_23517_, _15921_);
  and (_23518_, _23517_, _15571_);
  nor (_23520_, _23517_, _15571_);
  nor (_23521_, _23520_, _23518_);
  nor (_23522_, _16574_, _16249_);
  and (_23523_, _16574_, _16249_);
  nor (_23524_, _23523_, _23522_);
  nor (_23525_, _23524_, _23521_);
  and (_23526_, _23524_, _23521_);
  or (_23527_, _23526_, _23525_);
  nor (_23528_, _23527_, _23516_);
  and (_23529_, _23527_, _23516_);
  or (_23531_, _23529_, _23528_);
  nand (_23532_, _23531_, _03511_);
  nand (_23533_, _23532_, _23293_);
  or (_23534_, _23533_, _23506_);
  nand (_23535_, _23534_, _23294_);
  and (_23536_, _11389_, _03683_);
  nand (_23537_, _23536_, _23535_);
  or (_23538_, _23536_, _23234_);
  and (_23539_, _23538_, _03505_);
  and (_23540_, _23539_, _23537_);
  not (_23541_, _16909_);
  and (_23542_, _23541_, _08119_);
  nor (_23543_, _23541_, _08119_);
  nor (_23544_, _23543_, _23542_);
  nor (_23545_, _15870_, _23353_);
  and (_23546_, _15870_, _23353_);
  nor (_23547_, _23546_, _23545_);
  nor (_23548_, _23547_, _16254_);
  and (_23549_, _23547_, _16254_);
  nor (_23550_, _23549_, _23548_);
  not (_23552_, _16527_);
  nor (_23553_, _15576_, _15310_);
  and (_23554_, _15576_, _15310_);
  nor (_23555_, _23554_, _23553_);
  nor (_23556_, _23555_, _23552_);
  and (_23557_, _23555_, _23552_);
  nor (_23558_, _23557_, _23556_);
  not (_23559_, _23558_);
  and (_23560_, _23559_, _23550_);
  nor (_23561_, _23559_, _23550_);
  nor (_23563_, _23561_, _23560_);
  nand (_23564_, _23563_, _23544_);
  or (_23565_, _23563_, _23544_);
  and (_23566_, _23565_, _03504_);
  and (_23567_, _23566_, _23564_);
  or (_23568_, _23567_, _23540_);
  nor (_23569_, _03583_, _03621_);
  and (_23570_, _23569_, _03253_);
  and (_23571_, _23570_, _23568_);
  nor (_23572_, _04846_, _04551_);
  nor (_23574_, _11383_, _04741_);
  and (_23575_, _23574_, _23572_);
  and (_23576_, _23575_, _04837_);
  not (_23577_, _23570_);
  nand (_23578_, _23577_, _23234_);
  nand (_23579_, _23578_, _23576_);
  or (_23580_, _23579_, _23571_);
  or (_23581_, _23576_, _23234_);
  and (_23582_, _23581_, _06925_);
  and (_23583_, _23582_, _23580_);
  nor (_23585_, _15315_, _07379_);
  nor (_23586_, _15316_, _15074_);
  nor (_23587_, _23586_, _23585_);
  nor (_23588_, _23587_, _15581_);
  and (_23589_, _23587_, _15581_);
  nor (_23590_, _23589_, _23588_);
  nor (_23591_, _23590_, _15928_);
  and (_23592_, _23590_, _15928_);
  or (_23593_, _23592_, _23591_);
  not (_23594_, _23593_);
  nor (_23596_, _23594_, _16260_);
  and (_23597_, _23594_, _16260_);
  nor (_23598_, _23597_, _23596_);
  nor (_23599_, _23598_, _16521_);
  and (_23600_, _23598_, _16521_);
  or (_23601_, _23600_, _23599_);
  not (_23602_, _23601_);
  nor (_23603_, _23602_, _16914_);
  and (_23604_, _23602_, _16914_);
  nor (_23605_, _23604_, _23603_);
  and (_23606_, _23605_, _08124_);
  nor (_23607_, _23605_, _08124_);
  or (_23608_, _23607_, _23606_);
  and (_23609_, _23608_, _06919_);
  or (_23610_, _23609_, _23583_);
  and (_23611_, _11741_, _08881_);
  and (_23612_, _23611_, _23610_);
  not (_23613_, _23611_);
  and (_23614_, _23613_, _23234_);
  or (_23615_, _23614_, _10245_);
  or (_23617_, _23615_, _23612_);
  and (_23618_, _15324_, _15081_);
  or (_23619_, _23618_, _08145_);
  nor (_23620_, _23619_, _15599_);
  and (_23621_, _23619_, _15599_);
  nor (_23622_, _23621_, _23620_);
  nand (_23623_, _23622_, _15944_);
  or (_23624_, _23622_, _15944_);
  and (_23625_, _23624_, _23623_);
  or (_23626_, _23625_, _16278_);
  nand (_23628_, _23625_, _16278_);
  and (_23629_, _23628_, _23626_);
  nor (_23630_, _23629_, _16597_);
  and (_23631_, _23629_, _16597_);
  or (_23632_, _23631_, _23630_);
  nor (_23633_, _23632_, _16931_);
  and (_23634_, _23632_, _16931_);
  or (_23635_, _23634_, _23633_);
  nor (_23636_, _23635_, _08154_);
  and (_23637_, _23635_, _08154_);
  or (_23639_, _23637_, _23636_);
  or (_23640_, _23639_, _10244_);
  and (_23641_, _23640_, _10251_);
  and (_23642_, _23641_, _23617_);
  and (_23643_, _23639_, _10250_);
  or (_23644_, _23643_, _08032_);
  or (_23645_, _23644_, _23642_);
  not (_23646_, _16201_);
  nor (_23647_, _15256_, _08021_);
  and (_23648_, _15256_, _08021_);
  nor (_23650_, _23648_, _23647_);
  not (_23651_, _23650_);
  and (_23652_, _23651_, _15618_);
  nor (_23653_, _23651_, _15618_);
  nor (_23654_, _23653_, _23652_);
  and (_23655_, _23654_, _15960_);
  nor (_23656_, _23654_, _15960_);
  or (_23657_, _23656_, _23655_);
  and (_23658_, _23657_, _23646_);
  nor (_23659_, _23657_, _23646_);
  nor (_23661_, _23659_, _23658_);
  nor (_23662_, _23661_, _16518_);
  and (_23663_, _23661_, _16518_);
  nor (_23664_, _23663_, _23662_);
  nor (_23665_, _23664_, _16853_);
  and (_23666_, _23664_, _16853_);
  nor (_23667_, _23666_, _23665_);
  nor (_23668_, _23667_, _08031_);
  and (_23669_, _23667_, _08031_);
  or (_23670_, _23669_, _08128_);
  or (_23671_, _23670_, _23668_);
  and (_23672_, _23671_, _03640_);
  and (_23673_, _23672_, _23645_);
  and (_23674_, _15334_, _15088_);
  nor (_23675_, _15334_, _15088_);
  nor (_23676_, _23675_, _23674_);
  nor (_23677_, _23676_, _15632_);
  and (_23678_, _23676_, _15632_);
  nor (_23679_, _23678_, _23677_);
  nor (_23680_, _23679_, _15972_);
  and (_23682_, _23679_, _15972_);
  or (_23683_, _23682_, _23680_);
  nor (_23684_, _23683_, _16184_);
  and (_23685_, _23683_, _16184_);
  or (_23686_, _23685_, _23684_);
  and (_23687_, _23686_, _16612_);
  nor (_23688_, _23686_, _16612_);
  or (_23689_, _23688_, _23687_);
  nor (_23690_, _23689_, _16837_);
  and (_23691_, _23689_, _16837_);
  or (_23693_, _23691_, _23690_);
  nor (_23694_, _23693_, _08331_);
  and (_23695_, _23693_, _08331_);
  or (_23696_, _23695_, _23694_);
  and (_23697_, _23696_, _03635_);
  or (_23698_, _23697_, _08160_);
  or (_23699_, _23698_, _23673_);
  not (_23700_, _16298_);
  or (_23701_, _08390_, _08380_);
  and (_23702_, _23701_, _08391_);
  and (_23704_, _23702_, _15650_);
  nor (_23705_, _23702_, _15650_);
  or (_23706_, _23705_, _23704_);
  and (_23707_, _23706_, _15865_);
  nor (_23708_, _23706_, _15865_);
  or (_23709_, _23708_, _23707_);
  and (_23710_, _23709_, _23700_);
  nor (_23711_, _23709_, _23700_);
  nor (_23712_, _23711_, _23710_);
  or (_23713_, _23712_, _16629_);
  nand (_23715_, _23712_, _16629_);
  and (_23716_, _23715_, _23713_);
  nor (_23717_, _23716_, _16948_);
  and (_23718_, _23716_, _16948_);
  nor (_23719_, _23718_, _23717_);
  nor (_23720_, _23719_, _08414_);
  and (_23721_, _23719_, _08414_);
  or (_23722_, _23721_, _23720_);
  or (_23723_, _23722_, _08161_);
  and (_23724_, _23723_, _23699_);
  or (_23726_, _23724_, _03371_);
  nor (_23727_, _05301_, _05295_);
  nor (_23728_, _05291_, _03557_);
  and (_23729_, _23728_, _23727_);
  nor (_23730_, _23728_, _23727_);
  nor (_23731_, _23730_, _23729_);
  nor (_23732_, _05302_, _05361_);
  not (_23733_, _23732_);
  nor (_23734_, _05335_, _05328_);
  and (_23735_, _23734_, _23733_);
  nor (_23736_, _23734_, _23733_);
  nor (_23737_, _23736_, _23735_);
  nor (_23738_, _23737_, _23731_);
  and (_23739_, _23737_, _23731_);
  or (_23740_, _23739_, _23738_);
  or (_23741_, _23740_, _03285_);
  and (_23742_, _23741_, _03501_);
  and (_23743_, _23742_, _23726_);
  and (_23744_, _15345_, _15099_);
  nor (_23745_, _15345_, _15099_);
  or (_23747_, _23745_, _23744_);
  not (_23748_, _15983_);
  and (_23749_, _23748_, _15659_);
  nor (_23750_, _23748_, _15659_);
  nor (_23751_, _23750_, _23749_);
  and (_23752_, _23751_, _23747_);
  nor (_23753_, _23751_, _23747_);
  or (_23754_, _23753_, _23752_);
  nor (_23755_, _16638_, _16307_);
  and (_23756_, _16638_, _16307_);
  nor (_23758_, _23756_, _23755_);
  and (_23759_, _23758_, _16957_);
  nor (_23760_, _23758_, _16957_);
  nor (_23761_, _23760_, _23759_);
  nor (_23762_, _23761_, _23754_);
  and (_23763_, _23761_, _23754_);
  nor (_23764_, _23763_, _23762_);
  and (_23765_, _23764_, _08423_);
  nor (_23766_, _23764_, _08423_);
  or (_23767_, _23766_, _23765_);
  and (_23769_, _23767_, _03500_);
  nor (_23770_, _03656_, _03497_);
  not (_23771_, _23770_);
  or (_23772_, _23771_, _23769_);
  or (_23773_, _23772_, _23743_);
  or (_23774_, _23770_, _23234_);
  and (_23775_, _23774_, _06889_);
  and (_23776_, _23775_, _23773_);
  and (_23777_, _23463_, _07441_);
  or (_23778_, _23777_, _05969_);
  or (_23780_, _23778_, _23776_);
  and (_23781_, _15352_, _15106_);
  nor (_23782_, _15352_, _15106_);
  nor (_23783_, _23782_, _23781_);
  and (_23784_, _23783_, _15666_);
  nor (_23785_, _23783_, _15666_);
  or (_23786_, _23785_, _23784_);
  and (_23787_, _23786_, _15991_);
  nor (_23788_, _23786_, _15991_);
  or (_23789_, _23788_, _23787_);
  not (_23791_, _16646_);
  and (_23792_, _23791_, _16315_);
  nor (_23793_, _23791_, _16315_);
  nor (_23794_, _23793_, _23792_);
  nand (_23795_, _23794_, _16965_);
  or (_23796_, _23794_, _16965_);
  and (_23797_, _23796_, _23795_);
  or (_23798_, _23797_, _23789_);
  nand (_23799_, _23797_, _23789_);
  and (_23800_, _23799_, _23798_);
  nor (_23802_, _23800_, _08430_);
  and (_23803_, _23800_, _08430_);
  or (_23804_, _23803_, _05970_);
  or (_23805_, _23804_, _23802_);
  and (_23806_, _23805_, _03275_);
  and (_23807_, _23806_, _23780_);
  not (_23808_, _16970_);
  and (_23809_, _23808_, _08435_);
  nor (_23810_, _23808_, _08435_);
  nor (_23811_, _23810_, _23809_);
  and (_23813_, _15357_, _15023_);
  nor (_23814_, _15357_, _15023_);
  nor (_23815_, _23814_, _23813_);
  not (_23816_, _15997_);
  and (_23817_, _23816_, _15672_);
  nor (_23818_, _23816_, _15672_);
  nor (_23819_, _23818_, _23817_);
  nor (_23820_, _23819_, _23815_);
  and (_23821_, _23819_, _23815_);
  or (_23822_, _23821_, _23820_);
  not (_23823_, _16651_);
  and (_23824_, _23823_, _16320_);
  nor (_23825_, _23823_, _16320_);
  nor (_23826_, _23825_, _23824_);
  and (_23827_, _23826_, _23822_);
  nor (_23828_, _23826_, _23822_);
  nor (_23829_, _23828_, _23827_);
  or (_23830_, _23829_, _23811_);
  nand (_23831_, _23829_, _23811_);
  and (_23832_, _23831_, _03644_);
  and (_23834_, _23832_, _23830_);
  or (_23835_, _23834_, _23807_);
  and (_23836_, _23835_, _07805_);
  and (_23837_, _07515_, _16976_);
  nor (_23838_, _07515_, _16976_);
  nor (_23839_, _23838_, _23837_);
  nor (_23840_, _07648_, _07595_);
  and (_23841_, _07648_, _07595_);
  nor (_23842_, _23841_, _23840_);
  nor (_23843_, _23842_, _07545_);
  and (_23845_, _23842_, _07545_);
  nor (_23846_, _23845_, _23843_);
  nor (_23847_, _23846_, _23839_);
  and (_23848_, _23846_, _23839_);
  or (_23849_, _23848_, _23847_);
  nor (_23850_, _23849_, _07473_);
  and (_23851_, _23849_, _07473_);
  or (_23852_, _23851_, _23850_);
  and (_23853_, _23852_, _07724_);
  nor (_23854_, _23852_, _07724_);
  nor (_23856_, _23854_, _23853_);
  nor (_23857_, _23856_, _07803_);
  and (_23858_, _23856_, _07803_);
  or (_23859_, _23858_, _23857_);
  and (_23860_, _23859_, _07455_);
  or (_23861_, _23860_, _23836_);
  and (_23862_, _23861_, _03314_);
  nand (_23863_, _23740_, _03313_);
  nand (_23864_, _23863_, _23288_);
  or (_23865_, _23864_, _23862_);
  and (_23867_, _23865_, _23289_);
  or (_23868_, _23867_, _04816_);
  or (_23869_, _23234_, _04815_);
  and (_23870_, _23869_, _04582_);
  and (_23871_, _23870_, _23868_);
  nor (_23872_, _15367_, _15013_);
  and (_23873_, _15367_, _15013_);
  or (_23874_, _23873_, _23872_);
  nor (_23875_, _15845_, _15683_);
  and (_23876_, _15845_, _15683_);
  nor (_23878_, _23876_, _23875_);
  nor (_23879_, _23878_, _23874_);
  and (_23880_, _23878_, _23874_);
  or (_23881_, _23880_, _23879_);
  nor (_23882_, _16662_, _16331_);
  and (_23883_, _16662_, _16331_);
  nor (_23884_, _23883_, _23882_);
  and (_23885_, _23884_, _16983_);
  nor (_23886_, _23884_, _16983_);
  nor (_23887_, _23886_, _23885_);
  nor (_23888_, _23887_, _23881_);
  and (_23889_, _23887_, _23881_);
  nor (_23890_, _23889_, _23888_);
  and (_23891_, _23890_, _07939_);
  nor (_23892_, _23890_, _07939_);
  or (_23893_, _23892_, _23891_);
  and (_23894_, _23893_, _03650_);
  or (_23895_, _23894_, _23871_);
  and (_23896_, _23895_, _08446_);
  nand (_23897_, _23740_, _08445_);
  and (_23899_, _11822_, _11785_);
  and (_23900_, _23899_, _11827_);
  nand (_23901_, _23900_, _23897_);
  or (_23902_, _23901_, _23896_);
  or (_23903_, _23900_, _23234_);
  and (_23904_, _23903_, _16011_);
  and (_23905_, _23904_, _23902_);
  and (_23906_, _15123_, _08659_);
  nor (_23907_, _23906_, _15592_);
  nor (_23908_, _15834_, _08655_);
  and (_23910_, _15834_, _08655_);
  nor (_23911_, _23910_, _23908_);
  nor (_23912_, _23911_, _23907_);
  and (_23913_, _23911_, _23907_);
  nor (_23914_, _23913_, _23912_);
  nor (_23915_, _16498_, _08648_);
  and (_23916_, _16498_, _08648_);
  nor (_23917_, _23916_, _23915_);
  not (_23918_, _23917_);
  nor (_23919_, _08643_, _08466_);
  and (_23921_, _08643_, _08466_);
  nor (_23922_, _23921_, _23919_);
  and (_23923_, _23922_, _23918_);
  nor (_23924_, _23922_, _23918_);
  nor (_23925_, _23924_, _23923_);
  nand (_23926_, _23925_, _23914_);
  or (_23927_, _23925_, _23914_);
  and (_23928_, _23927_, _16012_);
  and (_23929_, _23928_, _23926_);
  or (_23930_, _23929_, _07952_);
  or (_23932_, _23930_, _23905_);
  not (_23933_, _08688_);
  nor (_23934_, _23933_, _08691_);
  and (_23935_, _23933_, _08691_);
  nor (_23936_, _23935_, _23934_);
  and (_23937_, _15006_, _08700_);
  nor (_23938_, _23937_, _15610_);
  nor (_23939_, _15950_, _08696_);
  and (_23940_, _15950_, _08696_);
  nor (_23941_, _23940_, _23939_);
  nor (_23943_, _23941_, _23938_);
  and (_23944_, _23941_, _23938_);
  nor (_23945_, _23944_, _23943_);
  nor (_23946_, _23945_, _23936_);
  and (_23947_, _23945_, _23936_);
  nor (_23948_, _23947_, _23946_);
  nor (_23949_, _23948_, _08685_);
  and (_23950_, _23948_, _08685_);
  or (_23951_, _23950_, _23949_);
  nor (_23952_, _23951_, _07955_);
  and (_23954_, _23951_, _07955_);
  or (_23955_, _23954_, _23952_);
  or (_23956_, _23955_, _07953_);
  and (_23957_, _23956_, _03777_);
  and (_23958_, _23957_, _23932_);
  and (_23959_, _12347_, _12145_);
  nor (_23960_, _12347_, _12145_);
  or (_23961_, _23960_, _23959_);
  nor (_23962_, _12619_, _12544_);
  and (_23963_, _12619_, _12544_);
  nor (_23965_, _23963_, _23962_);
  nor (_23966_, _23965_, _23961_);
  and (_23967_, _23965_, _23961_);
  nor (_23968_, _23967_, _23966_);
  or (_23969_, _23968_, _12957_);
  nand (_23970_, _23968_, _12957_);
  and (_23971_, _23970_, _23969_);
  or (_23972_, _23971_, _13160_);
  nand (_23973_, _23971_, _13160_);
  and (_23974_, _23973_, _23972_);
  or (_23976_, _23974_, _13374_);
  nand (_23977_, _23974_, _13374_);
  and (_23978_, _23977_, _23976_);
  nor (_23979_, _23978_, _06458_);
  and (_23980_, _23978_, _06458_);
  or (_23981_, _23980_, _23979_);
  or (_23982_, _23981_, _08472_);
  and (_23983_, _23982_, _11844_);
  or (_23984_, _23983_, _23958_);
  and (_23985_, _10130_, _08383_);
  nor (_23987_, _23985_, _10131_);
  and (_23988_, _10097_, _08785_);
  nor (_23989_, _23988_, _10098_);
  not (_23990_, _23989_);
  and (_23991_, _23990_, _23987_);
  nor (_23992_, _23990_, _23987_);
  nor (_23993_, _23992_, _23991_);
  and (_23994_, _10112_, _08780_);
  nor (_23995_, _23994_, _10113_);
  and (_23996_, _08775_, _08479_);
  nor (_23998_, _10114_, _23996_);
  and (_23999_, _23998_, _23995_);
  nor (_24000_, _23998_, _23995_);
  or (_24001_, _24000_, _23999_);
  not (_24002_, _24001_);
  nor (_24003_, _24002_, _23993_);
  and (_24004_, _24002_, _23993_);
  or (_24005_, _24004_, _24003_);
  or (_24006_, _24005_, _08473_);
  and (_24007_, _24006_, _04591_);
  and (_24009_, _24007_, _23984_);
  nor (_24010_, _15245_, _15017_);
  and (_24011_, _15245_, _15017_);
  nor (_24012_, _24011_, _24010_);
  and (_24013_, _24012_, _15517_);
  nor (_24014_, _24012_, _15517_);
  or (_24015_, _24014_, _24013_);
  nand (_24016_, _24015_, _16030_);
  or (_24017_, _24015_, _16030_);
  and (_24018_, _24017_, _24016_);
  nor (_24020_, _17012_, _16496_);
  and (_24021_, _17012_, _16496_);
  nor (_24022_, _24021_, _24020_);
  not (_24023_, _16168_);
  and (_24024_, _24023_, _07950_);
  nor (_24025_, _24023_, _07950_);
  nor (_24026_, _24025_, _24024_);
  nor (_24027_, _24026_, _24022_);
  and (_24028_, _24026_, _24022_);
  nor (_24029_, _24028_, _24027_);
  nand (_24031_, _24029_, _24018_);
  or (_24032_, _24029_, _24018_);
  and (_24033_, _24032_, _03649_);
  and (_24034_, _24033_, _24031_);
  or (_24035_, _24034_, _24009_);
  and (_24036_, _24035_, _04589_);
  nand (_24037_, _23234_, _03778_);
  or (_24038_, _24037_, _05371_);
  nor (_24039_, _11856_, _03231_);
  nand (_24040_, _24039_, _24038_);
  or (_24042_, _24040_, _24036_);
  or (_24043_, _24039_, _23234_);
  and (_24044_, _24043_, _08487_);
  and (_24045_, _24044_, _24042_);
  and (_24046_, _23283_, _08490_);
  or (_24047_, _24046_, _04200_);
  or (_24048_, _24047_, _24045_);
  and (_24049_, _24048_, _23284_);
  or (_24050_, _24049_, _04198_);
  or (_24051_, _08701_, _08698_);
  nand (_24053_, _08701_, _08698_);
  and (_24054_, _24053_, _24051_);
  not (_24055_, _08692_);
  and (_24056_, _24055_, _08694_);
  nor (_24057_, _24055_, _08694_);
  nor (_24058_, _24057_, _24056_);
  not (_24059_, _24058_);
  and (_24060_, _24059_, _24054_);
  nor (_24061_, _24059_, _24054_);
  nor (_24062_, _24061_, _24060_);
  nor (_24064_, _08686_, _08689_);
  and (_24065_, _08686_, _08689_);
  nor (_24066_, _24065_, _24064_);
  nor (_24067_, _24066_, _08683_);
  and (_24068_, _24066_, _08683_);
  nor (_24069_, _24068_, _24067_);
  not (_24070_, _24069_);
  and (_24071_, _24070_, _24062_);
  nor (_24072_, _24070_, _24062_);
  or (_24073_, _24072_, _24071_);
  nand (_24075_, _24073_, _07954_);
  or (_24076_, _24073_, _07954_);
  and (_24077_, _24076_, _24075_);
  or (_24078_, _24077_, _07944_);
  and (_24079_, _24078_, _03772_);
  and (_24080_, _24079_, _24050_);
  nor (_24081_, _12345_, _12144_);
  and (_24082_, _12345_, _12144_);
  nor (_24083_, _24082_, _24081_);
  not (_24084_, _12617_);
  and (_24086_, _24084_, _12542_);
  nor (_24087_, _24084_, _12542_);
  nor (_24088_, _24087_, _24086_);
  and (_24089_, _24088_, _24083_);
  nor (_24090_, _24088_, _24083_);
  nor (_24091_, _24090_, _24089_);
  not (_24092_, _13372_);
  nor (_24093_, _13158_, _12955_);
  and (_24094_, _13158_, _12955_);
  nor (_24095_, _24094_, _24093_);
  nor (_24097_, _24095_, _24092_);
  and (_24098_, _24095_, _24092_);
  nor (_24099_, _24098_, _24097_);
  and (_24100_, _24099_, _24091_);
  nor (_24101_, _24099_, _24091_);
  or (_24102_, _24101_, _24100_);
  nor (_24103_, _24102_, _06456_);
  and (_24104_, _24102_, _06456_);
  or (_24105_, _24104_, _07942_);
  or (_24106_, _24105_, _24103_);
  and (_24108_, _24106_, _11368_);
  or (_24109_, _24108_, _24080_);
  not (_24110_, _08778_);
  or (_24111_, _08787_, _08381_);
  nand (_24112_, _08787_, _08381_);
  and (_24113_, _24112_, _24111_);
  not (_24114_, _08781_);
  and (_24115_, _24114_, _08783_);
  nor (_24116_, _24114_, _08783_);
  nor (_24117_, _24116_, _24115_);
  not (_24119_, _24117_);
  and (_24120_, _24119_, _24113_);
  nor (_24121_, _24119_, _24113_);
  nor (_24122_, _24121_, _24120_);
  nand (_24123_, _24122_, _24110_);
  or (_24124_, _24122_, _24110_);
  and (_24125_, _24124_, _24123_);
  or (_24126_, _24125_, _08776_);
  nand (_24127_, _24125_, _08776_);
  and (_24128_, _24127_, _24126_);
  or (_24130_, _24128_, _08772_);
  nand (_24131_, _24128_, _08772_);
  and (_24132_, _24131_, _24130_);
  and (_24133_, _24132_, _08477_);
  nor (_24134_, _24132_, _08477_);
  or (_24135_, _24134_, _24133_);
  or (_24136_, _24135_, _08500_);
  and (_24137_, _24136_, _04596_);
  and (_24138_, _24137_, _24109_);
  and (_24139_, _11364_, _10776_);
  nor (_24141_, _15724_, _15014_);
  and (_24142_, _15724_, _15014_);
  nor (_24143_, _24142_, _24141_);
  nor (_24144_, _17034_, _16381_);
  and (_24145_, _17034_, _16381_);
  nor (_24146_, _24145_, _24144_);
  and (_24147_, _24146_, _24143_);
  nor (_24148_, _24146_, _24143_);
  nor (_24149_, _24148_, _24147_);
  nor (_24150_, _16703_, _15846_);
  and (_24152_, _16703_, _15846_);
  nor (_24153_, _24152_, _24150_);
  nor (_24154_, _15242_, _07940_);
  and (_24155_, _15242_, _07940_);
  nor (_24156_, _24155_, _24154_);
  and (_24157_, _24156_, _24153_);
  nor (_24158_, _24156_, _24153_);
  nor (_24159_, _24158_, _24157_);
  not (_24160_, _24159_);
  nand (_24161_, _24160_, _24149_);
  or (_24163_, _24160_, _24149_);
  and (_24164_, _24163_, _03655_);
  nand (_24165_, _24164_, _24161_);
  nand (_24166_, _24165_, _24139_);
  or (_24167_, _24166_, _24138_);
  or (_24168_, _23234_, _24139_);
  and (_24169_, _24168_, _16383_);
  and (_24170_, _24169_, _24167_);
  nor (_24171_, _15122_, _08658_);
  and (_24172_, _15122_, _08658_);
  nor (_24175_, _24172_, _24171_);
  not (_24176_, _24175_);
  nor (_24177_, _08650_, _08654_);
  and (_24178_, _08650_, _08654_);
  nor (_24179_, _24178_, _24177_);
  nor (_24180_, _24179_, _24176_);
  and (_24181_, _24179_, _24176_);
  nor (_24182_, _24181_, _24180_);
  not (_24183_, _08645_);
  nor (_24184_, _08647_, _08642_);
  and (_24187_, _08647_, _08642_);
  nor (_24188_, _24187_, _24184_);
  nor (_24189_, _24188_, _24183_);
  and (_24190_, _24188_, _24183_);
  nor (_24191_, _24190_, _24189_);
  not (_24192_, _24191_);
  nor (_24193_, _24192_, _24182_);
  and (_24194_, _24192_, _24182_);
  or (_24195_, _24194_, _24193_);
  and (_24196_, _24195_, _08459_);
  nor (_24199_, _24195_, _08459_);
  or (_24200_, _24199_, _24196_);
  and (_24201_, _24200_, _16384_);
  or (_24202_, _24201_, _04207_);
  or (_24203_, _24202_, _24170_);
  nor (_24204_, _15005_, _08699_);
  and (_24205_, _15005_, _08699_);
  nor (_24206_, _24205_, _24204_);
  not (_24207_, _24206_);
  not (_24208_, _08693_);
  and (_24211_, _24208_, _08695_);
  nor (_24212_, _24208_, _08695_);
  nor (_24213_, _24212_, _24211_);
  nor (_24214_, _24213_, _24207_);
  and (_24215_, _24213_, _24207_);
  nor (_24216_, _24215_, _24214_);
  not (_24217_, _08687_);
  nor (_24218_, _08690_, _08684_);
  and (_24219_, _08690_, _08684_);
  nor (_24220_, _24219_, _24218_);
  nor (_24223_, _24220_, _24217_);
  and (_24224_, _24220_, _24217_);
  nor (_24225_, _24224_, _24223_);
  nor (_24226_, _24225_, _24216_);
  and (_24227_, _24225_, _24216_);
  nor (_24228_, _24227_, _24226_);
  nor (_24229_, _24228_, _07935_);
  and (_24230_, _24228_, _07935_);
  nor (_24231_, _24230_, _24229_);
  nand (_24232_, _24231_, _04207_);
  and (_24235_, _24232_, _03785_);
  and (_24236_, _24235_, _24203_);
  nor (_24237_, _12346_, _12015_);
  and (_24238_, _12346_, _12015_);
  nor (_24239_, _24238_, _24237_);
  and (_24240_, _24239_, _12543_);
  nor (_24241_, _24239_, _12543_);
  or (_24242_, _24241_, _24240_);
  nand (_24243_, _24242_, _12618_);
  or (_24244_, _24242_, _12618_);
  and (_24247_, _24244_, _24243_);
  nor (_24248_, _13159_, _12956_);
  and (_24249_, _13159_, _12956_);
  nor (_24250_, _24249_, _24248_);
  nor (_24251_, _24250_, _13373_);
  and (_24252_, _24250_, _13373_);
  nor (_24253_, _24252_, _24251_);
  not (_24254_, _24253_);
  nor (_24255_, _24254_, _24247_);
  and (_24256_, _24254_, _24247_);
  nor (_24258_, _24256_, _24255_);
  or (_24259_, _24258_, _06457_);
  nand (_24260_, _24258_, _06457_);
  and (_24261_, _24260_, _03784_);
  and (_24262_, _24261_, _24259_);
  or (_24263_, _24262_, _08524_);
  or (_24264_, _24263_, _24236_);
  nor (_24265_, _10129_, _08382_);
  and (_24266_, _10129_, _08382_);
  nor (_24267_, _24266_, _24265_);
  not (_24269_, _24267_);
  not (_24270_, _08782_);
  and (_24271_, _24270_, _08784_);
  nor (_24272_, _24270_, _08784_);
  nor (_24273_, _24272_, _24271_);
  and (_24274_, _24273_, _24269_);
  nor (_24275_, _24273_, _24269_);
  nor (_24276_, _24275_, _24274_);
  nor (_24277_, _08777_, _08773_);
  and (_24278_, _08777_, _08773_);
  nor (_24280_, _24278_, _24277_);
  and (_24281_, _24280_, _08779_);
  nor (_24282_, _24280_, _08779_);
  nor (_24283_, _24282_, _24281_);
  nor (_24284_, _24283_, _24276_);
  and (_24285_, _24283_, _24276_);
  or (_24286_, _24285_, _24284_);
  and (_24287_, _24286_, _08478_);
  nor (_24288_, _24286_, _08478_);
  or (_24289_, _24288_, _24287_);
  or (_24291_, _24289_, _08525_);
  and (_24292_, _24291_, _04608_);
  and (_24293_, _24292_, _24264_);
  and (_24294_, _11894_, _11890_);
  nor (_24295_, _15437_, _15184_);
  and (_24296_, _15437_, _15184_);
  or (_24297_, _24296_, _24295_);
  nor (_24298_, _16079_, _15748_);
  and (_24299_, _16079_, _15748_);
  nor (_24300_, _24299_, _24298_);
  nor (_24302_, _24300_, _24297_);
  and (_24303_, _24300_, _24297_);
  nor (_24304_, _24303_, _24302_);
  nor (_24305_, _16813_, _16491_);
  and (_24306_, _16813_, _16491_);
  nor (_24307_, _24306_, _24305_);
  not (_24308_, _16400_);
  and (_24309_, _24308_, _08534_);
  nor (_24310_, _24308_, _08534_);
  nor (_24311_, _24310_, _24309_);
  nor (_24313_, _24311_, _24307_);
  and (_24314_, _24311_, _24307_);
  nor (_24315_, _24314_, _24313_);
  not (_24316_, _24315_);
  nand (_24317_, _24316_, _24304_);
  or (_24318_, _24316_, _24304_);
  and (_24319_, _24318_, _03653_);
  nand (_24320_, _24319_, _24317_);
  nand (_24321_, _24320_, _24294_);
  or (_24322_, _24321_, _24293_);
  or (_24324_, _23234_, _24294_);
  and (_24325_, _24324_, _24322_);
  and (_24326_, _03589_, _03247_);
  or (_24327_, _24326_, _07932_);
  or (_24328_, _24327_, _24325_);
  not (_24329_, _04219_);
  not (_24330_, _15840_);
  nor (_24331_, _08144_, _07910_);
  nor (_24332_, _15442_, _15081_);
  nor (_24333_, _24332_, _24331_);
  nor (_24335_, _24333_, _15753_);
  and (_24336_, _24333_, _15753_);
  nor (_24337_, _24336_, _24335_);
  and (_24338_, _24337_, _24330_);
  nor (_24339_, _24337_, _24330_);
  nor (_24340_, _24339_, _24338_);
  and (_24341_, _24340_, _16406_);
  nor (_24342_, _24340_, _16406_);
  nor (_24343_, _24342_, _24341_);
  nor (_24344_, _24343_, _16723_);
  and (_24346_, _24343_, _16723_);
  or (_24347_, _24346_, _24344_);
  nor (_24348_, _24347_, _17059_);
  and (_24349_, _24347_, _17059_);
  or (_24350_, _24349_, _24348_);
  and (_24351_, _24350_, _07930_);
  nor (_24352_, _24350_, _07930_);
  or (_24353_, _24352_, _24351_);
  and (_24354_, _24353_, _24329_);
  or (_24355_, _24354_, _07933_);
  and (_24357_, _24355_, _24328_);
  and (_24358_, _24353_, _04219_);
  or (_24359_, _24358_, _08539_);
  or (_24360_, _24359_, _24357_);
  not (_24361_, _16087_);
  nor (_24362_, _15447_, _08021_);
  and (_24363_, _15447_, _08021_);
  or (_24364_, _24363_, _24362_);
  nor (_24365_, _24364_, _15759_);
  and (_24366_, _24364_, _15759_);
  nor (_24368_, _24366_, _24365_);
  and (_24369_, _24368_, _24361_);
  nor (_24370_, _24368_, _24361_);
  nor (_24371_, _24370_, _24369_);
  and (_24372_, _24371_, _16411_);
  nor (_24373_, _24371_, _16411_);
  nor (_24374_, _24373_, _24372_);
  nor (_24375_, _24374_, _16728_);
  and (_24376_, _24374_, _16728_);
  or (_24377_, _24376_, _24375_);
  and (_24379_, _24377_, _17065_);
  nor (_24380_, _24377_, _17065_);
  or (_24381_, _24380_, _24379_);
  nor (_24382_, _24381_, _08565_);
  and (_24383_, _24381_, _08565_);
  or (_24384_, _24383_, _08541_);
  or (_24385_, _24384_, _24382_);
  and (_24386_, _24385_, _03783_);
  and (_24387_, _24386_, _24360_);
  not (_24388_, _16092_);
  nor (_24390_, _15452_, _15088_);
  and (_24391_, _15452_, _15088_);
  or (_24392_, _24391_, _24390_);
  nor (_24393_, _24392_, _15764_);
  and (_24394_, _24392_, _15764_);
  nor (_24395_, _24394_, _24393_);
  and (_24396_, _24395_, _24388_);
  nor (_24397_, _24395_, _24388_);
  nor (_24398_, _24397_, _24396_);
  nor (_24399_, _24398_, _16417_);
  and (_24401_, _24398_, _16417_);
  or (_24402_, _24401_, _24399_);
  and (_24403_, _24402_, _16734_);
  nor (_24404_, _24402_, _16734_);
  nor (_24405_, _24404_, _24403_);
  and (_24406_, _24405_, _17070_);
  nor (_24407_, _24405_, _17070_);
  or (_24408_, _24407_, _24406_);
  nor (_24409_, _24408_, _08596_);
  and (_24410_, _24408_, _08596_);
  or (_24412_, _24410_, _24409_);
  and (_24413_, _24412_, _03782_);
  or (_24414_, _24413_, _08569_);
  or (_24415_, _24414_, _24387_);
  and (_24416_, _15457_, _08380_);
  nor (_24417_, _15457_, _08380_);
  nor (_24418_, _24417_, _24416_);
  nor (_24419_, _24418_, _15770_);
  and (_24420_, _24418_, _15770_);
  nor (_24421_, _24420_, _24419_);
  and (_24423_, _24421_, _16098_);
  nor (_24424_, _24421_, _16098_);
  nor (_24425_, _24424_, _24423_);
  nor (_24426_, _24425_, _16422_);
  and (_24427_, _24425_, _16422_);
  or (_24428_, _24427_, _24426_);
  nor (_24429_, _24428_, _16739_);
  and (_24430_, _24428_, _16739_);
  or (_24431_, _24430_, _24429_);
  nor (_24432_, _24431_, _17076_);
  and (_24434_, _24431_, _17076_);
  or (_24435_, _24434_, _24432_);
  nand (_24436_, _24435_, _08627_);
  or (_24437_, _24435_, _08627_);
  and (_24438_, _24437_, _24436_);
  or (_24439_, _24438_, _08602_);
  and (_24440_, _24439_, _08601_);
  and (_24441_, _24440_, _24415_);
  nor (_24442_, _08385_, _08384_);
  nor (_24443_, _15545_, \oc8051_golden_model_1.ACC [3]);
  and (_24445_, _15545_, \oc8051_golden_model_1.ACC [3]);
  nor (_24446_, _24445_, _24443_);
  and (_24447_, _24446_, _23342_);
  nor (_24448_, _24446_, _23342_);
  nor (_24449_, _24448_, _24447_);
  not (_24450_, _24449_);
  nand (_24451_, _24450_, _24442_);
  or (_24452_, _24450_, _24442_);
  and (_24453_, _24452_, _24451_);
  nand (_24454_, _24453_, _08600_);
  and (_24456_, _10796_, _03796_);
  nand (_24457_, _24456_, _24454_);
  or (_24458_, _24457_, _24441_);
  nor (_24459_, _24456_, _23234_);
  nor (_24460_, _24459_, _08632_);
  and (_24461_, _24460_, _24458_);
  and (_24462_, _23258_, _08632_);
  nor (_24463_, _24462_, _24461_);
  nor (_24464_, _24463_, _08634_);
  and (_24465_, _23258_, _08634_);
  or (_24467_, _24465_, _08638_);
  or (_24468_, _24467_, _24464_);
  and (_24469_, _24468_, _23259_);
  or (_24470_, _24469_, _08679_);
  nor (_24471_, _15005_, _08700_);
  and (_24472_, _15005_, _08700_);
  nor (_24473_, _24472_, _24471_);
  and (_24474_, _24473_, _15783_);
  nor (_24475_, _24473_, _15783_);
  nor (_24476_, _24475_, _24474_);
  and (_24478_, _24476_, _16110_);
  nor (_24479_, _24476_, _16110_);
  nor (_24480_, _24479_, _24478_);
  and (_24481_, _24480_, _16436_);
  nor (_24482_, _24480_, _16436_);
  nor (_24483_, _24482_, _24481_);
  nor (_24484_, _24483_, _16753_);
  and (_24485_, _24483_, _16753_);
  or (_24486_, _24485_, _24484_);
  nor (_24487_, _24486_, _17099_);
  and (_24489_, _24486_, _17099_);
  nor (_24490_, _24489_, _24487_);
  nand (_24491_, _24490_, _08716_);
  or (_24492_, _24490_, _08716_);
  and (_24493_, _24492_, _24491_);
  or (_24494_, _24493_, _10369_);
  and (_24495_, _24494_, _03525_);
  and (_24496_, _24495_, _24470_);
  nor (_24497_, _15474_, _09943_);
  and (_24498_, _15474_, _09943_);
  or (_24500_, _24498_, _24497_);
  and (_24501_, _24500_, _15788_);
  nor (_24502_, _24500_, _15788_);
  nor (_24503_, _24502_, _24501_);
  and (_24504_, _24503_, _16116_);
  nor (_24505_, _24503_, _16116_);
  or (_24506_, _24505_, _24504_);
  nor (_24507_, _24506_, _16441_);
  and (_24508_, _24506_, _16441_);
  or (_24509_, _24508_, _24507_);
  nor (_24511_, _24509_, _16759_);
  and (_24512_, _24509_, _16759_);
  or (_24513_, _24512_, _24511_);
  nor (_24514_, _24513_, _16807_);
  and (_24515_, _24513_, _16807_);
  or (_24516_, _24515_, _24514_);
  or (_24517_, _24516_, _08765_);
  nand (_24518_, _24516_, _08765_);
  and (_24519_, _24518_, _03524_);
  and (_24520_, _24519_, _24517_);
  or (_24522_, _24520_, _08720_);
  or (_24523_, _24522_, _24496_);
  nor (_24524_, _03975_, _03953_);
  nor (_24525_, _24524_, _03170_);
  not (_24526_, _24525_);
  not (_24527_, _13180_);
  nor (_24528_, _08769_, _03521_);
  and (_24529_, _24528_, _24527_);
  nor (_24530_, _03519_, _03246_);
  not (_24531_, _24530_);
  nor (_24533_, _03668_, _04050_);
  nor (_24534_, _24533_, _04253_);
  nor (_24535_, _24534_, _24531_);
  and (_24536_, _24535_, _24529_);
  and (_24537_, _24536_, _24526_);
  not (_24538_, _10129_);
  and (_24539_, _24538_, _08383_);
  nor (_24540_, _24538_, _08383_);
  nor (_24541_, _24540_, _24539_);
  and (_24542_, _24541_, _15793_);
  nor (_24544_, _24541_, _15793_);
  nor (_24545_, _24544_, _24542_);
  and (_24546_, _24545_, _16123_);
  nor (_24547_, _24545_, _16123_);
  nor (_24548_, _24547_, _24546_);
  and (_24549_, _24548_, _16447_);
  nor (_24550_, _24548_, _16447_);
  nor (_24551_, _24550_, _24549_);
  nor (_24552_, _24551_, _16766_);
  and (_24553_, _24551_, _16766_);
  or (_24555_, _24553_, _24552_);
  and (_24556_, _24555_, _17106_);
  nor (_24557_, _24555_, _17106_);
  or (_24558_, _24557_, _24556_);
  nor (_24559_, _24558_, _08802_);
  and (_24560_, _24558_, _08802_);
  or (_24561_, _24560_, _08771_);
  or (_24562_, _24561_, _24559_);
  and (_24563_, _24562_, _24537_);
  and (_24564_, _24563_, _24523_);
  nor (_24566_, _04618_, _04250_);
  not (_24567_, _24537_);
  nand (_24568_, _24567_, _23234_);
  nand (_24569_, _24568_, _24566_);
  or (_24570_, _24569_, _24564_);
  or (_24571_, _24566_, _23234_);
  and (_24572_, _24571_, _04260_);
  and (_24573_, _24572_, _24570_);
  and (_24574_, _23374_, _03809_);
  or (_24575_, _24574_, _08809_);
  or (_24577_, _24575_, _24573_);
  not (_24578_, _08815_);
  and (_24579_, _15545_, _24578_);
  and (_24580_, _24579_, \oc8051_golden_model_1.ACC [3]);
  nor (_24581_, _24579_, \oc8051_golden_model_1.ACC [3]);
  nor (_24582_, _24581_, _24580_);
  and (_24583_, _24582_, _16460_);
  nor (_24584_, _24582_, _16460_);
  nor (_24585_, _24584_, _24583_);
  and (_24586_, _16777_, _07484_);
  nor (_24588_, _16777_, _07484_);
  nor (_24589_, _24588_, _24586_);
  nor (_24590_, _24589_, _24585_);
  and (_24591_, _24589_, _24585_);
  or (_24592_, _24591_, _24590_);
  nor (_24593_, _24592_, _08821_);
  and (_24594_, _24592_, _08821_);
  nor (_24595_, _24594_, _24593_);
  nand (_24596_, _24595_, _08809_);
  and (_24597_, _24596_, _09690_);
  and (_24599_, _24597_, _24577_);
  and (_24600_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_24601_, _24600_, _08084_);
  or (_24602_, _24601_, _24449_);
  nand (_24603_, _24601_, _24449_);
  and (_24604_, _24603_, _24602_);
  nand (_24605_, _24604_, _08814_);
  nand (_24606_, _24605_, _04625_);
  or (_24607_, _24606_, _24599_);
  or (_24608_, _23234_, _04625_);
  and (_24611_, _24608_, _03206_);
  and (_24612_, _24611_, _24607_);
  and (_24613_, _23531_, _03205_);
  or (_24614_, _24613_, _06827_);
  or (_24615_, _24614_, _24612_);
  and (_24616_, _24615_, _23235_);
  or (_24617_, _24616_, _04271_);
  or (_24618_, _23234_, _06833_);
  and (_24619_, _24618_, _03820_);
  and (_24620_, _24619_, _24617_);
  not (_24622_, _16147_);
  nor (_24623_, _16472_, _24622_);
  and (_24624_, _16472_, _24622_);
  nor (_24625_, _24624_, _24623_);
  nor (_24626_, _24625_, _17129_);
  and (_24627_, _24625_, _17129_);
  nor (_24628_, _24627_, _24626_);
  nor (_24629_, _15498_, _15044_);
  and (_24630_, _15498_, _15044_);
  nor (_24631_, _24630_, _24629_);
  and (_24633_, _24631_, _15817_);
  nor (_24634_, _24631_, _15817_);
  nor (_24635_, _24634_, _24633_);
  and (_24636_, _24635_, _16790_);
  nor (_24637_, _24635_, _16790_);
  or (_24638_, _24637_, _24636_);
  and (_24639_, _24638_, _08834_);
  nor (_24640_, _24638_, _08834_);
  or (_24641_, _24640_, _24639_);
  not (_24642_, _24641_);
  nand (_24644_, _24642_, _24628_);
  or (_24645_, _24642_, _24628_);
  and (_24646_, _24645_, _03816_);
  and (_24647_, _24646_, _24644_);
  or (_24648_, _24647_, _24620_);
  and (_24649_, _24648_, _08832_);
  nor (_24650_, _11982_, _03242_);
  nor (_24651_, _08838_, _03684_);
  and (_24652_, _24651_, _24650_);
  not (_24653_, _08839_);
  and (_24655_, _15545_, _24653_);
  and (_24656_, _24655_, _07628_);
  nor (_24657_, _24655_, _07628_);
  nor (_24658_, _24657_, _24656_);
  nor (_24659_, _24658_, _16477_);
  and (_24660_, _24658_, _16477_);
  or (_24661_, _24660_, _24659_);
  and (_24662_, _24661_, _17134_);
  nor (_24663_, _24661_, _17134_);
  nor (_24664_, _24663_, _24662_);
  not (_24666_, _24664_);
  nor (_24667_, _16795_, _08846_);
  and (_24668_, _16795_, _08846_);
  nor (_24669_, _24668_, _24667_);
  nand (_24670_, _24669_, _24666_);
  or (_24671_, _24669_, _24666_);
  and (_24672_, _24671_, _08831_);
  nand (_24673_, _24672_, _24670_);
  nand (_24674_, _24673_, _24652_);
  or (_24675_, _24674_, _24649_);
  or (_24677_, _24652_, _23234_);
  and (_24678_, _24677_, _43227_);
  and (_24679_, _24678_, _24675_);
  or (_24680_, _24679_, _23218_);
  and (_43512_, _24680_, _41991_);
  not (_24681_, \oc8051_golden_model_1.PSW [1]);
  nor (_24682_, _05368_, _24681_);
  and (_24683_, _05368_, _05898_);
  or (_24684_, _24683_, _24682_);
  or (_24685_, _24684_, _04524_);
  or (_24687_, _05368_, \oc8051_golden_model_1.PSW [1]);
  and (_24688_, _12234_, _05368_);
  not (_24689_, _24688_);
  and (_24690_, _24689_, _24687_);
  or (_24691_, _24690_, _04515_);
  nand (_24692_, _05368_, _03320_);
  and (_24693_, _24692_, _24687_);
  and (_24694_, _24693_, _04499_);
  nor (_24695_, _04499_, _24681_);
  or (_24696_, _24695_, _03599_);
  or (_24698_, _24696_, _24694_);
  and (_24699_, _24698_, _03516_);
  and (_24700_, _24699_, _24691_);
  nor (_24701_, _06000_, _24681_);
  and (_24702_, _12238_, _06000_);
  or (_24703_, _24702_, _24701_);
  and (_24704_, _24703_, _03515_);
  or (_24705_, _24704_, _03597_);
  or (_24706_, _24705_, _24700_);
  and (_24707_, _24706_, _24685_);
  or (_24709_, _24707_, _03603_);
  or (_24710_, _24693_, _03611_);
  and (_24711_, _24710_, _03512_);
  and (_24712_, _24711_, _24709_);
  and (_24713_, _12224_, _06000_);
  or (_24714_, _24713_, _24701_);
  and (_24715_, _24714_, _03511_);
  or (_24716_, _24715_, _03504_);
  or (_24717_, _24716_, _24712_);
  and (_24718_, _24702_, _12253_);
  or (_24720_, _24701_, _03505_);
  or (_24721_, _24720_, _24718_);
  and (_24722_, _24721_, _24717_);
  and (_24723_, _24722_, _03501_);
  not (_24724_, _06000_);
  nor (_24725_, _12270_, _24724_);
  or (_24726_, _24701_, _24725_);
  and (_24727_, _24726_, _03500_);
  or (_24728_, _24727_, _07441_);
  or (_24729_, _24728_, _24723_);
  or (_24731_, _24684_, _06889_);
  and (_24732_, _24731_, _24729_);
  or (_24733_, _24732_, _05969_);
  and (_24734_, _06835_, _05368_);
  or (_24735_, _24682_, _05970_);
  or (_24736_, _24735_, _24734_);
  and (_24737_, _24736_, _03275_);
  and (_24738_, _24737_, _24733_);
  nor (_24739_, _12330_, _09709_);
  or (_24740_, _24739_, _24682_);
  and (_24742_, _24740_, _03644_);
  or (_24743_, _24742_, _24738_);
  and (_24744_, _24743_, _03651_);
  or (_24745_, _12220_, _09709_);
  and (_24746_, _24745_, _03649_);
  nand (_24747_, _05368_, _04347_);
  and (_24748_, _24747_, _03650_);
  or (_24749_, _24748_, _24746_);
  and (_24750_, _24749_, _24687_);
  or (_24751_, _24750_, _24744_);
  and (_24753_, _24751_, _04589_);
  or (_24754_, _12347_, _09709_);
  and (_24755_, _24687_, _03778_);
  and (_24756_, _24755_, _24754_);
  or (_24757_, _24756_, _24753_);
  and (_24758_, _24757_, _04596_);
  or (_24759_, _12219_, _09709_);
  and (_24760_, _24687_, _03655_);
  and (_24761_, _24760_, _24759_);
  or (_24762_, _24761_, _24758_);
  and (_24764_, _24762_, _04594_);
  or (_24765_, _24682_, _05699_);
  and (_24766_, _24693_, _03773_);
  and (_24767_, _24766_, _24765_);
  or (_24768_, _24767_, _24764_);
  and (_24769_, _24768_, _03787_);
  or (_24770_, _24747_, _05699_);
  and (_24771_, _24687_, _03653_);
  and (_24772_, _24771_, _24770_);
  or (_24773_, _24692_, _05699_);
  and (_24775_, _24687_, _03786_);
  and (_24776_, _24775_, _24773_);
  or (_24777_, _24776_, _03809_);
  or (_24778_, _24777_, _24772_);
  or (_24779_, _24778_, _24769_);
  or (_24780_, _24690_, _04260_);
  and (_24781_, _24780_, _03206_);
  and (_24782_, _24781_, _24779_);
  and (_24783_, _24714_, _03205_);
  or (_24784_, _24783_, _03816_);
  or (_24786_, _24784_, _24782_);
  or (_24787_, _24682_, _03820_);
  or (_24788_, _24787_, _24688_);
  and (_24789_, _24788_, _24786_);
  or (_24790_, _24789_, _43231_);
  or (_24791_, _43227_, \oc8051_golden_model_1.PSW [1]);
  and (_24792_, _24791_, _41991_);
  and (_43513_, _24792_, _24790_);
  and (_24793_, _07859_, \oc8051_golden_model_1.ACC [7]);
  nor (_24794_, _07859_, \oc8051_golden_model_1.ACC [7]);
  nor (_24796_, _24794_, _09702_);
  nor (_24797_, _24796_, _24793_);
  nand (_24798_, _24797_, _07930_);
  and (_24799_, _24793_, _07927_);
  nor (_24800_, _24799_, _07933_);
  and (_24801_, _24800_, _24798_);
  not (_24802_, \oc8051_golden_model_1.PSW [2]);
  nor (_24803_, _05368_, _24802_);
  not (_24804_, _24803_);
  or (_24805_, _12524_, _09709_);
  and (_24807_, _24805_, _24804_);
  or (_24808_, _24807_, _03275_);
  or (_24809_, _09709_, _05130_);
  and (_24810_, _24809_, _24804_);
  and (_24811_, _24810_, _07441_);
  nor (_24812_, _07962_, \oc8051_golden_model_1.ACC [7]);
  and (_24813_, _07962_, \oc8051_golden_model_1.ACC [7]);
  nor (_24814_, _24813_, _24812_);
  and (_24815_, _24814_, _10272_);
  nor (_24816_, _24814_, _10272_);
  or (_24818_, _24816_, _24815_);
  or (_24819_, _24818_, _08031_);
  nand (_24820_, _24818_, _08031_);
  and (_24821_, _24820_, _24819_);
  and (_24822_, _24821_, _08032_);
  not (_24823_, _07860_);
  and (_24824_, _10258_, _24823_);
  nor (_24825_, _10258_, _24823_);
  nor (_24826_, _24825_, _24824_);
  nor (_24827_, _24826_, _08151_);
  and (_24829_, _24826_, _08151_);
  or (_24830_, _24829_, _24827_);
  or (_24831_, _24830_, _08037_);
  nor (_24832_, _06000_, _24802_);
  and (_24833_, _12414_, _06000_);
  nor (_24834_, _24833_, _24832_);
  or (_24835_, _24834_, _03512_);
  and (_24836_, _24810_, _03597_);
  nor (_24837_, _12430_, _09709_);
  nor (_24838_, _24837_, _24803_);
  and (_24840_, _24838_, _03599_);
  and (_24841_, _05368_, \oc8051_golden_model_1.ACC [2]);
  nor (_24842_, _24841_, _24803_);
  or (_24843_, _24842_, _04500_);
  or (_24844_, _04499_, _24802_);
  and (_24845_, _24844_, _04515_);
  and (_24846_, _24845_, _24843_);
  or (_24847_, _24846_, _03515_);
  or (_24848_, _24847_, _24840_);
  not (_24849_, _24832_);
  nand (_24851_, _12416_, _06000_);
  and (_24852_, _24851_, _24849_);
  or (_24853_, _24852_, _03516_);
  and (_24854_, _24853_, _04524_);
  and (_24855_, _24854_, _24848_);
  or (_24856_, _24855_, _24836_);
  and (_24857_, _24856_, _03611_);
  and (_24858_, _24842_, _03603_);
  or (_24859_, _24858_, _03511_);
  or (_24860_, _24859_, _24857_);
  and (_24862_, _24860_, _24835_);
  or (_24863_, _24862_, _03504_);
  and (_24864_, _24849_, _10157_);
  or (_24865_, _24864_, _03505_);
  or (_24866_, _24865_, _24852_);
  and (_24867_, _24866_, _06925_);
  and (_24868_, _24867_, _24863_);
  or (_24869_, _14345_, _14236_);
  or (_24870_, _24869_, _14459_);
  or (_24871_, _24870_, _14578_);
  or (_24873_, _24871_, _14694_);
  or (_24874_, _24873_, _14811_);
  or (_24875_, _24874_, _07437_);
  nor (_24876_, _24875_, _14929_);
  or (_24877_, _24876_, _08038_);
  or (_24878_, _24877_, _24868_);
  and (_24879_, _24878_, _08128_);
  and (_24880_, _24879_, _24831_);
  or (_24881_, _24880_, _03635_);
  or (_24882_, _24881_, _24822_);
  nor (_24884_, _08273_, \oc8051_golden_model_1.ACC [7]);
  and (_24885_, _08273_, \oc8051_golden_model_1.ACC [7]);
  nor (_24886_, _24885_, _24884_);
  not (_24887_, _24886_);
  or (_24888_, _24887_, _09725_);
  nand (_24889_, _24887_, _09725_);
  and (_24890_, _24889_, _24888_);
  nand (_24891_, _24890_, _08331_);
  or (_24892_, _24890_, _08331_);
  and (_24893_, _24892_, _24891_);
  or (_24895_, _24893_, _03640_);
  and (_24896_, _24895_, _08161_);
  and (_24897_, _24896_, _24882_);
  and (_24898_, _08339_, \oc8051_golden_model_1.ACC [7]);
  nor (_24899_, _08339_, \oc8051_golden_model_1.ACC [7]);
  nor (_24900_, _24899_, _24898_);
  not (_24901_, _24900_);
  or (_24902_, _24901_, _10288_);
  nand (_24903_, _24901_, _10288_);
  and (_24904_, _24903_, _24902_);
  nand (_24906_, _24904_, _08414_);
  or (_24907_, _24904_, _08414_);
  and (_24908_, _24907_, _24906_);
  and (_24909_, _24908_, _08160_);
  or (_24910_, _24909_, _03500_);
  or (_24911_, _24910_, _24897_);
  or (_24912_, _12465_, _24724_);
  and (_24913_, _24912_, _24849_);
  or (_24914_, _24913_, _03501_);
  and (_24915_, _24914_, _06889_);
  and (_24917_, _24915_, _24911_);
  or (_24918_, _24917_, _24811_);
  and (_24919_, _24918_, _05970_);
  or (_24920_, _06714_, _09709_);
  nor (_24921_, _24803_, _05970_);
  and (_24922_, _24921_, _24920_);
  or (_24923_, _24922_, _03644_);
  or (_24924_, _24923_, _24919_);
  and (_24925_, _24924_, _24808_);
  or (_24926_, _24925_, _07455_);
  nor (_24928_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_24929_, _24928_, _07483_);
  nand (_24930_, _24929_, _07455_);
  and (_24931_, _24930_, _03651_);
  and (_24932_, _24931_, _24926_);
  nand (_24933_, _12538_, _05368_);
  nor (_24934_, _24803_, _04591_);
  and (_24935_, _24934_, _24933_);
  and (_24936_, _05368_, _06414_);
  nor (_24937_, _24936_, _24803_);
  and (_24939_, _24937_, _03650_);
  or (_24940_, _24939_, _03778_);
  or (_24941_, _24940_, _24935_);
  or (_24942_, _24941_, _24932_);
  nand (_24943_, _12544_, _05368_);
  and (_24944_, _24943_, _24804_);
  or (_24945_, _24944_, _04589_);
  and (_24946_, _24945_, _24942_);
  or (_24947_, _24946_, _03655_);
  and (_24948_, _24804_, _05792_);
  or (_24950_, _24937_, _04596_);
  or (_24951_, _24950_, _24948_);
  and (_24952_, _24951_, _24947_);
  or (_24953_, _24952_, _03773_);
  or (_24954_, _24842_, _04594_);
  or (_24955_, _24954_, _24948_);
  and (_24956_, _24955_, _04608_);
  and (_24957_, _24956_, _24953_);
  or (_24958_, _12537_, _09709_);
  nor (_24959_, _24803_, _04608_);
  and (_24961_, _24959_, _24958_);
  or (_24962_, _24961_, _03786_);
  or (_24963_, _24962_, _24957_);
  or (_24964_, _12543_, _09709_);
  and (_24965_, _24964_, _24804_);
  or (_24966_, _24965_, _04606_);
  and (_24967_, _24966_, _07933_);
  and (_24968_, _24967_, _24963_);
  or (_24969_, _24968_, _24801_);
  and (_24970_, _24969_, _08541_);
  nand (_24972_, _24813_, _08562_);
  nor (_24973_, _24812_, _10345_);
  nor (_24974_, _24973_, _24813_);
  nand (_24975_, _24974_, _08565_);
  and (_24976_, _24975_, _24972_);
  and (_24977_, _24976_, _08539_);
  or (_24978_, _24977_, _03782_);
  or (_24979_, _24978_, _24970_);
  nand (_24980_, _24885_, _08593_);
  nor (_24981_, _24887_, _10351_);
  nor (_24983_, _24981_, _24885_);
  nand (_24984_, _24983_, _08596_);
  and (_24985_, _24984_, _24980_);
  or (_24986_, _24985_, _03783_);
  and (_24987_, _24986_, _08602_);
  and (_24988_, _24987_, _24979_);
  and (_24989_, _24900_, _10357_);
  or (_24990_, _24989_, _24898_);
  and (_24991_, _24990_, _08627_);
  nor (_24992_, _24990_, _08627_);
  or (_24994_, _24992_, _24991_);
  and (_24995_, _24994_, _08569_);
  or (_24996_, _24995_, _10362_);
  or (_24997_, _24996_, _24988_);
  not (_24998_, _07946_);
  and (_24999_, _08672_, _24998_);
  or (_25000_, _24999_, _09697_);
  and (_25001_, _25000_, _10369_);
  nand (_25002_, _25001_, _24997_);
  not (_25003_, _07935_);
  nor (_25005_, _08713_, _25003_);
  and (_25006_, _08713_, _07954_);
  or (_25007_, _25006_, _10369_);
  or (_25008_, _25007_, _25005_);
  and (_25009_, _25008_, _08721_);
  and (_25010_, _25009_, _25002_);
  or (_25011_, _08762_, _08723_);
  and (_25012_, _25011_, _10379_);
  nand (_25013_, _08799_, _09691_);
  and (_25014_, _25013_, _09693_);
  or (_25016_, _25014_, _03809_);
  or (_25017_, _25016_, _25012_);
  or (_25018_, _25017_, _25010_);
  nand (_25019_, _24838_, _03809_);
  and (_25020_, _25019_, _03206_);
  and (_25021_, _25020_, _25018_);
  nor (_25022_, _24834_, _03206_);
  or (_25023_, _25022_, _03816_);
  or (_25024_, _25023_, _25021_);
  and (_25025_, _12600_, _05368_);
  or (_25027_, _24803_, _03820_);
  or (_25028_, _25027_, _25025_);
  and (_25029_, _25028_, _25024_);
  or (_25030_, _25029_, _43231_);
  or (_25031_, _43227_, \oc8051_golden_model_1.PSW [2]);
  and (_25032_, _25031_, _41991_);
  and (_43514_, _25032_, _25030_);
  nor (_25033_, _05368_, _04957_);
  and (_25034_, _05368_, _06347_);
  nor (_25035_, _25034_, _25033_);
  and (_25037_, _25035_, _03650_);
  nor (_25038_, _09709_, _04944_);
  nor (_25039_, _25038_, _25033_);
  and (_25040_, _25039_, _07441_);
  and (_25041_, _05368_, \oc8051_golden_model_1.ACC [3]);
  nor (_25042_, _25041_, _25033_);
  nor (_25043_, _25042_, _04500_);
  nor (_25044_, _04499_, _04957_);
  or (_25045_, _25044_, _25043_);
  and (_25046_, _25045_, _04515_);
  nor (_25048_, _12625_, _09709_);
  nor (_25049_, _25048_, _25033_);
  nor (_25050_, _25049_, _04515_);
  or (_25051_, _25050_, _25046_);
  and (_25052_, _25051_, _03516_);
  nor (_25053_, _06000_, _04957_);
  and (_25054_, _12638_, _06000_);
  nor (_25055_, _25054_, _25053_);
  nor (_25056_, _25055_, _03516_);
  or (_25057_, _25056_, _03597_);
  or (_25059_, _25057_, _25052_);
  nand (_25060_, _25039_, _03597_);
  and (_25061_, _25060_, _25059_);
  and (_25062_, _25061_, _03611_);
  nor (_25063_, _25042_, _03611_);
  or (_25064_, _25063_, _25062_);
  and (_25065_, _25064_, _03512_);
  and (_25066_, _12622_, _06000_);
  nor (_25067_, _25066_, _25053_);
  nor (_25068_, _25067_, _03512_);
  or (_25070_, _25068_, _03504_);
  or (_25071_, _25070_, _25065_);
  nor (_25072_, _25053_, _12653_);
  nor (_25073_, _25072_, _25055_);
  or (_25074_, _25073_, _03505_);
  and (_25075_, _25074_, _03501_);
  and (_25076_, _25075_, _25071_);
  nor (_25077_, _12671_, _24724_);
  nor (_25078_, _25077_, _25053_);
  nor (_25079_, _25078_, _03501_);
  nor (_25081_, _25079_, _07441_);
  not (_25082_, _25081_);
  nor (_25083_, _25082_, _25076_);
  nor (_25084_, _25083_, _25040_);
  nor (_25085_, _25084_, _05969_);
  and (_25086_, _06838_, _05368_);
  nor (_25087_, _25033_, _05970_);
  not (_25088_, _25087_);
  nor (_25089_, _25088_, _25086_);
  or (_25090_, _25089_, _03644_);
  nor (_25091_, _25090_, _25085_);
  nor (_25092_, _12731_, _09709_);
  nor (_25093_, _25033_, _25092_);
  nor (_25094_, _25093_, _03275_);
  or (_25095_, _25094_, _03650_);
  nor (_25096_, _25095_, _25091_);
  nor (_25097_, _25096_, _25037_);
  or (_25098_, _25097_, _03649_);
  and (_25099_, _12746_, _05368_);
  or (_25100_, _25099_, _25033_);
  or (_25103_, _25100_, _04591_);
  and (_25104_, _25103_, _04589_);
  and (_25105_, _25104_, _25098_);
  and (_25106_, _12619_, _05368_);
  nor (_25107_, _25106_, _25033_);
  nor (_25108_, _25107_, _04589_);
  nor (_25109_, _25108_, _25105_);
  nor (_25110_, _25109_, _03655_);
  nor (_25111_, _25033_, _05650_);
  not (_25112_, _25111_);
  nor (_25114_, _25035_, _04596_);
  and (_25115_, _25114_, _25112_);
  nor (_25116_, _25115_, _25110_);
  nor (_25117_, _25116_, _03773_);
  nor (_25118_, _25042_, _04594_);
  and (_25119_, _25118_, _25112_);
  nor (_25120_, _25119_, _03653_);
  not (_25121_, _25120_);
  nor (_25122_, _25121_, _25117_);
  nor (_25123_, _12745_, _09709_);
  or (_25125_, _25033_, _04608_);
  nor (_25126_, _25125_, _25123_);
  or (_25127_, _25126_, _03786_);
  nor (_25128_, _25127_, _25122_);
  nor (_25129_, _12618_, _09709_);
  nor (_25130_, _25129_, _25033_);
  nor (_25131_, _25130_, _04606_);
  or (_25132_, _25131_, _25128_);
  and (_25133_, _25132_, _04260_);
  nor (_25134_, _25049_, _04260_);
  or (_25135_, _25134_, _25133_);
  and (_25136_, _25135_, _03206_);
  nor (_25137_, _25067_, _03206_);
  or (_25138_, _25137_, _25136_);
  and (_25139_, _25138_, _03820_);
  and (_25140_, _12806_, _05368_);
  nor (_25141_, _25140_, _25033_);
  nor (_25142_, _25141_, _03820_);
  or (_25143_, _25142_, _25139_);
  or (_25144_, _25143_, _43231_);
  or (_25147_, _43227_, \oc8051_golden_model_1.PSW [3]);
  and (_25148_, _25147_, _41991_);
  and (_43515_, _25148_, _25144_);
  not (_25149_, \oc8051_golden_model_1.PSW [4]);
  nor (_25150_, _05368_, _25149_);
  nor (_25151_, _05840_, _09709_);
  nor (_25152_, _25151_, _25150_);
  and (_25153_, _25152_, _07441_);
  nor (_25154_, _06000_, _25149_);
  and (_25155_, _12853_, _06000_);
  nor (_25157_, _25155_, _25154_);
  nor (_25158_, _25157_, _03512_);
  and (_25159_, _05368_, \oc8051_golden_model_1.ACC [4]);
  nor (_25160_, _25159_, _25150_);
  nor (_25161_, _25160_, _04500_);
  nor (_25162_, _04499_, _25149_);
  or (_25163_, _25162_, _25161_);
  and (_25164_, _25163_, _04515_);
  nor (_25165_, _12820_, _09709_);
  nor (_25166_, _25165_, _25150_);
  nor (_25167_, _25166_, _04515_);
  or (_25168_, _25167_, _25164_);
  and (_25169_, _25168_, _03516_);
  and (_25170_, _12830_, _06000_);
  nor (_25171_, _25170_, _25154_);
  nor (_25172_, _25171_, _03516_);
  or (_25173_, _25172_, _03597_);
  or (_25174_, _25173_, _25169_);
  nand (_25175_, _25152_, _03597_);
  and (_25176_, _25175_, _25174_);
  and (_25179_, _25176_, _03611_);
  nor (_25180_, _25160_, _03611_);
  or (_25181_, _25180_, _25179_);
  and (_25182_, _25181_, _03512_);
  nor (_25183_, _25182_, _25158_);
  nor (_25184_, _25183_, _03504_);
  nor (_25185_, _25154_, _12860_);
  or (_25186_, _25171_, _03505_);
  nor (_25187_, _25186_, _25185_);
  nor (_25188_, _25187_, _25184_);
  nor (_25190_, _25188_, _03500_);
  nor (_25191_, _12828_, _24724_);
  nor (_25192_, _25191_, _25154_);
  nor (_25193_, _25192_, _03501_);
  nor (_25194_, _25193_, _07441_);
  not (_25195_, _25194_);
  nor (_25196_, _25195_, _25190_);
  nor (_25197_, _25196_, _25153_);
  nor (_25198_, _25197_, _05969_);
  and (_25199_, _06843_, _05368_);
  nor (_25201_, _25150_, _05970_);
  not (_25202_, _25201_);
  nor (_25203_, _25202_, _25199_);
  nor (_25204_, _25203_, _03644_);
  not (_25205_, _25204_);
  nor (_25206_, _25205_, _25198_);
  nor (_25207_, _12936_, _09709_);
  nor (_25208_, _25207_, _25150_);
  nor (_25209_, _25208_, _03275_);
  or (_25210_, _25209_, _08861_);
  or (_25212_, _25210_, _25206_);
  and (_25213_, _12951_, _05368_);
  or (_25214_, _25150_, _04591_);
  or (_25215_, _25214_, _25213_);
  and (_25216_, _06375_, _05368_);
  nor (_25217_, _25216_, _25150_);
  and (_25218_, _25217_, _03650_);
  nor (_25219_, _25218_, _03778_);
  and (_25220_, _25219_, _25215_);
  and (_25221_, _25220_, _25212_);
  and (_25222_, _12957_, _05368_);
  nor (_25223_, _25222_, _25150_);
  nor (_25224_, _25223_, _04589_);
  nor (_25225_, _25224_, _25221_);
  nor (_25226_, _25225_, _03655_);
  nor (_25227_, _25150_, _05889_);
  not (_25228_, _25227_);
  nor (_25229_, _25217_, _04596_);
  and (_25230_, _25229_, _25228_);
  nor (_25231_, _25230_, _25226_);
  nor (_25234_, _25231_, _03773_);
  nor (_25235_, _25160_, _04594_);
  and (_25236_, _25235_, _25228_);
  nor (_25237_, _25236_, _03653_);
  not (_25238_, _25237_);
  nor (_25239_, _25238_, _25234_);
  nor (_25240_, _12949_, _09709_);
  or (_25241_, _25150_, _04608_);
  nor (_25242_, _25241_, _25240_);
  or (_25243_, _25242_, _03786_);
  nor (_25245_, _25243_, _25239_);
  nor (_25246_, _12956_, _09709_);
  nor (_25247_, _25246_, _25150_);
  nor (_25248_, _25247_, _04606_);
  or (_25249_, _25248_, _25245_);
  and (_25250_, _25249_, _04260_);
  nor (_25251_, _25166_, _04260_);
  or (_25252_, _25251_, _25250_);
  and (_25253_, _25252_, _03206_);
  nor (_25254_, _25157_, _03206_);
  or (_25256_, _25254_, _25253_);
  and (_25257_, _25256_, _03820_);
  and (_25258_, _13013_, _05368_);
  nor (_25259_, _25258_, _25150_);
  nor (_25260_, _25259_, _03820_);
  or (_25261_, _25260_, _25257_);
  or (_25262_, _25261_, _43231_);
  or (_25263_, _43227_, \oc8051_golden_model_1.PSW [4]);
  and (_25264_, _25263_, _41991_);
  and (_43516_, _25264_, _25262_);
  not (_25266_, \oc8051_golden_model_1.PSW [5]);
  nor (_25267_, _05368_, _25266_);
  and (_25268_, _06842_, _05368_);
  or (_25269_, _25268_, _25267_);
  and (_25270_, _25269_, _05969_);
  and (_25271_, _05368_, \oc8051_golden_model_1.ACC [5]);
  nor (_25272_, _25271_, _25267_);
  nor (_25273_, _25272_, _04500_);
  nor (_25274_, _04499_, _25266_);
  or (_25275_, _25274_, _25273_);
  and (_25277_, _25275_, _04515_);
  nor (_25278_, _13035_, _09709_);
  nor (_25279_, _25278_, _25267_);
  nor (_25280_, _25279_, _04515_);
  or (_25281_, _25280_, _25277_);
  and (_25282_, _25281_, _03516_);
  nor (_25283_, _06000_, _25266_);
  and (_25284_, _13051_, _06000_);
  nor (_25285_, _25284_, _25283_);
  nor (_25286_, _25285_, _03516_);
  or (_25288_, _25286_, _03597_);
  or (_25289_, _25288_, _25282_);
  nor (_25290_, _05552_, _09709_);
  nor (_25291_, _25290_, _25267_);
  nand (_25292_, _25291_, _03597_);
  and (_25293_, _25292_, _25289_);
  and (_25294_, _25293_, _03611_);
  nor (_25295_, _25272_, _03611_);
  or (_25296_, _25295_, _25294_);
  and (_25297_, _25296_, _03512_);
  and (_25299_, _13032_, _06000_);
  nor (_25300_, _25299_, _25283_);
  nor (_25301_, _25300_, _03512_);
  or (_25302_, _25301_, _25297_);
  and (_25303_, _25302_, _03505_);
  nor (_25304_, _25283_, _13066_);
  nor (_25305_, _25304_, _25285_);
  and (_25306_, _25305_, _03504_);
  or (_25307_, _25306_, _25303_);
  and (_25308_, _25307_, _03501_);
  nor (_25310_, _13030_, _24724_);
  nor (_25311_, _25310_, _25283_);
  nor (_25312_, _25311_, _03501_);
  nor (_25313_, _25312_, _07441_);
  not (_25314_, _25313_);
  nor (_25315_, _25314_, _25308_);
  and (_25316_, _25291_, _07441_);
  or (_25317_, _25316_, _05969_);
  nor (_25318_, _25317_, _25315_);
  or (_25319_, _25318_, _25270_);
  and (_25321_, _25319_, _03275_);
  nor (_25322_, _13139_, _09709_);
  nor (_25323_, _25322_, _25267_);
  nor (_25324_, _25323_, _03275_);
  or (_25325_, _25324_, _08861_);
  or (_25326_, _25325_, _25321_);
  and (_25327_, _13154_, _05368_);
  or (_25328_, _25267_, _04591_);
  or (_25329_, _25328_, _25327_);
  and (_25330_, _06358_, _05368_);
  nor (_25332_, _25330_, _25267_);
  and (_25333_, _25332_, _03650_);
  nor (_25334_, _25333_, _03778_);
  and (_25335_, _25334_, _25329_);
  and (_25336_, _25335_, _25326_);
  and (_25337_, _13160_, _05368_);
  nor (_25338_, _25337_, _25267_);
  nor (_25339_, _25338_, _04589_);
  nor (_25340_, _25339_, _25336_);
  nor (_25341_, _25340_, _03655_);
  nor (_25343_, _25267_, _05601_);
  not (_25344_, _25343_);
  nor (_25345_, _25332_, _04596_);
  and (_25346_, _25345_, _25344_);
  nor (_25347_, _25346_, _25341_);
  nor (_25348_, _25347_, _03773_);
  nor (_25349_, _25272_, _04594_);
  and (_25350_, _25349_, _25344_);
  nor (_25351_, _25350_, _03653_);
  not (_25352_, _25351_);
  nor (_25353_, _25352_, _25348_);
  nor (_25354_, _13152_, _09709_);
  or (_25355_, _25267_, _04608_);
  nor (_25356_, _25355_, _25354_);
  or (_25357_, _25356_, _03786_);
  nor (_25358_, _25357_, _25353_);
  nor (_25359_, _13159_, _09709_);
  nor (_25360_, _25359_, _25267_);
  nor (_25361_, _25360_, _04606_);
  or (_25362_, _25361_, _25358_);
  and (_25365_, _25362_, _04260_);
  nor (_25366_, _25279_, _04260_);
  or (_25367_, _25366_, _25365_);
  and (_25368_, _25367_, _03206_);
  nor (_25369_, _25300_, _03206_);
  or (_25370_, _25369_, _25368_);
  and (_25371_, _25370_, _03820_);
  and (_25372_, _13217_, _05368_);
  nor (_25373_, _25372_, _25267_);
  nor (_25374_, _25373_, _03820_);
  or (_25376_, _25374_, _25371_);
  or (_25377_, _25376_, _43231_);
  or (_25378_, _43227_, \oc8051_golden_model_1.PSW [5]);
  and (_25379_, _25378_, _41991_);
  and (_43517_, _25379_, _25377_);
  not (_25380_, _08587_);
  nor (_25381_, _25380_, _08242_);
  nor (_25382_, _25381_, _03783_);
  nor (_25383_, _05368_, _15892_);
  nor (_25384_, _05442_, _09709_);
  nor (_25386_, _25384_, _25383_);
  and (_25387_, _25386_, _07441_);
  nor (_25388_, _08242_, _03640_);
  and (_25389_, _25388_, _08321_);
  nor (_25390_, _08024_, _07980_);
  nor (_25391_, _25390_, _08128_);
  or (_25392_, _08037_, _07874_);
  nor (_25393_, _25392_, _08147_);
  nor (_25394_, _06000_, _15892_);
  and (_25395_, _13251_, _06000_);
  nor (_25397_, _25395_, _25394_);
  nor (_25398_, _25397_, _03512_);
  and (_25399_, _05368_, \oc8051_golden_model_1.ACC [6]);
  nor (_25400_, _25399_, _25383_);
  nor (_25401_, _25400_, _04500_);
  nor (_25402_, _04499_, _15892_);
  or (_25403_, _25402_, _25401_);
  and (_25404_, _25403_, _04515_);
  nor (_25405_, _13235_, _09709_);
  nor (_25406_, _25405_, _25383_);
  nor (_25408_, _25406_, _04515_);
  or (_25409_, _25408_, _25404_);
  and (_25410_, _25409_, _03516_);
  and (_25411_, _13266_, _06000_);
  nor (_25412_, _25411_, _25394_);
  nor (_25413_, _25412_, _03516_);
  or (_25414_, _25413_, _03597_);
  or (_25415_, _25414_, _25410_);
  nand (_25416_, _25386_, _03597_);
  and (_25417_, _25416_, _25415_);
  and (_25419_, _25417_, _03611_);
  nor (_25420_, _25400_, _03611_);
  or (_25421_, _25420_, _25419_);
  and (_25422_, _25421_, _03512_);
  nor (_25423_, _25422_, _25398_);
  nor (_25424_, _25423_, _03504_);
  nor (_25425_, _25394_, _13281_);
  or (_25426_, _25412_, _03505_);
  or (_25427_, _25426_, _25425_);
  and (_25428_, _25427_, _08037_);
  not (_25430_, _25428_);
  nor (_25431_, _25430_, _25424_);
  or (_25432_, _25431_, _08032_);
  nor (_25433_, _25432_, _25393_);
  nor (_25434_, _25433_, _03635_);
  not (_25435_, _25434_);
  nor (_25436_, _25435_, _25391_);
  nor (_25437_, _25436_, _25389_);
  nor (_25438_, _25437_, _08160_);
  or (_25439_, _08336_, _08161_);
  nor (_25441_, _25439_, _08404_);
  or (_25442_, _25441_, _03500_);
  nor (_25443_, _25442_, _25438_);
  nor (_25444_, _13249_, _24724_);
  nor (_25445_, _25444_, _25394_);
  nor (_25446_, _25445_, _03501_);
  nor (_25447_, _25446_, _07441_);
  not (_25448_, _25447_);
  nor (_25449_, _25448_, _25443_);
  nor (_25450_, _25449_, _25387_);
  nor (_25452_, _25450_, _05969_);
  and (_25453_, _06531_, _05368_);
  nor (_25454_, _25383_, _05970_);
  not (_25455_, _25454_);
  nor (_25456_, _25455_, _25453_);
  nor (_25457_, _25456_, _03644_);
  not (_25458_, _25457_);
  nor (_25459_, _25458_, _25452_);
  nor (_25460_, _13356_, _09709_);
  nor (_25461_, _25460_, _25383_);
  nor (_25463_, _25461_, _03275_);
  or (_25464_, _25463_, _08861_);
  or (_25465_, _25464_, _25459_);
  and (_25466_, _13245_, _05368_);
  or (_25467_, _25383_, _04591_);
  or (_25468_, _25467_, _25466_);
  and (_25469_, _13363_, _05368_);
  nor (_25470_, _25469_, _25383_);
  and (_25471_, _25470_, _03650_);
  nor (_25472_, _25471_, _03778_);
  and (_25474_, _25472_, _25468_);
  and (_25475_, _25474_, _25465_);
  and (_25476_, _13374_, _05368_);
  nor (_25477_, _25476_, _25383_);
  nor (_25478_, _25477_, _04589_);
  nor (_25479_, _25478_, _25475_);
  nor (_25480_, _25479_, _03655_);
  nor (_25481_, _25383_, _05491_);
  not (_25482_, _25481_);
  nor (_25483_, _25470_, _04596_);
  and (_25485_, _25483_, _25482_);
  nor (_25486_, _25485_, _25480_);
  nor (_25487_, _25486_, _03773_);
  nor (_25488_, _25400_, _04594_);
  and (_25489_, _25488_, _25482_);
  or (_25490_, _25489_, _25487_);
  and (_25491_, _25490_, _04608_);
  nor (_25492_, _13243_, _09709_);
  nor (_25493_, _25492_, _25383_);
  nor (_25494_, _25493_, _04608_);
  or (_25496_, _25494_, _25491_);
  and (_25497_, _25496_, _04606_);
  nor (_25498_, _13373_, _09709_);
  nor (_25499_, _25498_, _25383_);
  nor (_25500_, _25499_, _04606_);
  nor (_25501_, _25500_, _07932_);
  not (_25502_, _25501_);
  nor (_25503_, _25502_, _25497_);
  not (_25504_, _07874_);
  and (_25505_, _07921_, _25504_);
  and (_25507_, _25505_, _07932_);
  or (_25508_, _25507_, _07931_);
  nor (_25509_, _25508_, _25503_);
  not (_25510_, _07931_);
  nor (_25511_, _25505_, _25510_);
  nor (_25512_, _25511_, _08539_);
  not (_25513_, _25512_);
  nor (_25514_, _25513_, _25509_);
  nor (_25515_, _08541_, _07980_);
  and (_25516_, _25515_, _08556_);
  nor (_25518_, _25516_, _03782_);
  not (_25519_, _25518_);
  nor (_25520_, _25519_, _25514_);
  nor (_25521_, _25520_, _25382_);
  nor (_25522_, _25521_, _08569_);
  not (_25523_, _08336_);
  and (_25524_, _08618_, _25523_);
  nor (_25525_, _25524_, _08602_);
  nor (_25526_, _25525_, _08635_);
  not (_25527_, _25526_);
  nor (_25528_, _25527_, _25522_);
  nor (_25529_, _08666_, _08640_);
  nor (_25530_, _25529_, _08638_);
  not (_25531_, _25530_);
  nor (_25532_, _25531_, _25528_);
  and (_25533_, _08666_, _08638_);
  nor (_25534_, _25533_, _08679_);
  not (_25535_, _25534_);
  nor (_25536_, _25535_, _25532_);
  or (_25537_, _08707_, _10369_);
  and (_25540_, _25537_, _03525_);
  not (_25541_, _25540_);
  nor (_25542_, _25541_, _25536_);
  and (_25543_, _08756_, _03524_);
  or (_25544_, _25543_, _08720_);
  nor (_25545_, _25544_, _25542_);
  nor (_25546_, _08793_, _08771_);
  nor (_25547_, _25546_, _25545_);
  and (_25548_, _25547_, _04260_);
  nor (_25549_, _25406_, _04260_);
  or (_25551_, _25549_, _25548_);
  and (_25552_, _25551_, _03206_);
  nor (_25553_, _25397_, _03206_);
  or (_25554_, _25553_, _25552_);
  and (_25555_, _25554_, _03820_);
  and (_25556_, _13425_, _05368_);
  nor (_25557_, _25383_, _25556_);
  nor (_25558_, _25557_, _03820_);
  or (_25559_, _25558_, _25555_);
  or (_25560_, _25559_, _43231_);
  or (_25562_, _43227_, \oc8051_golden_model_1.PSW [6]);
  and (_25563_, _25562_, _41991_);
  and (_43518_, _25563_, _25560_);
  not (_25564_, \oc8051_golden_model_1.PCON [0]);
  nor (_25565_, _05323_, _25564_);
  nor (_25566_, _05744_, _10403_);
  nor (_25567_, _25566_, _25565_);
  and (_25568_, _25567_, _17220_);
  and (_25569_, _05323_, _04491_);
  nor (_25570_, _25569_, _25565_);
  and (_25572_, _25570_, _07441_);
  and (_25573_, _05323_, \oc8051_golden_model_1.ACC [0]);
  nor (_25574_, _25573_, _25565_);
  nor (_25575_, _25574_, _03611_);
  nor (_25576_, _25574_, _04500_);
  nor (_25577_, _04499_, _25564_);
  or (_25578_, _25577_, _25576_);
  and (_25579_, _25578_, _04515_);
  nor (_25580_, _25567_, _04515_);
  or (_25581_, _25580_, _25579_);
  and (_25583_, _25581_, _04524_);
  nor (_25584_, _25570_, _04524_);
  nor (_25585_, _25584_, _25583_);
  nor (_25586_, _25585_, _03603_);
  or (_25587_, _25586_, _07441_);
  nor (_25588_, _25587_, _25575_);
  nor (_25589_, _25588_, _25572_);
  nor (_25590_, _25589_, _05969_);
  and (_25591_, _06836_, _05323_);
  nor (_25592_, _25565_, _05970_);
  not (_25594_, _25592_);
  nor (_25595_, _25594_, _25591_);
  nor (_25596_, _25595_, _25590_);
  nor (_25597_, _25596_, _03644_);
  nor (_25598_, _12129_, _10403_);
  or (_25599_, _25565_, _03275_);
  nor (_25600_, _25599_, _25598_);
  or (_25601_, _25600_, _03650_);
  nor (_25602_, _25601_, _25597_);
  and (_25603_, _05323_, _06366_);
  nor (_25605_, _25603_, _25565_);
  nand (_25606_, _25605_, _04591_);
  and (_25607_, _25606_, _08861_);
  nor (_25608_, _25607_, _25602_);
  and (_25609_, _12019_, _05323_);
  nor (_25610_, _25609_, _25565_);
  and (_25611_, _25610_, _03649_);
  nor (_25612_, _25611_, _25608_);
  nor (_25613_, _25612_, _03778_);
  and (_25614_, _12145_, _05323_);
  or (_25616_, _25565_, _04589_);
  nor (_25617_, _25616_, _25614_);
  or (_25618_, _25617_, _03655_);
  nor (_25619_, _25618_, _25613_);
  or (_25620_, _25605_, _04596_);
  nor (_25621_, _25620_, _25566_);
  nor (_25622_, _25621_, _25619_);
  nor (_25623_, _25622_, _03773_);
  and (_25624_, _12144_, _05323_);
  or (_25625_, _25624_, _25565_);
  and (_25627_, _25625_, _03773_);
  or (_25628_, _25627_, _25623_);
  and (_25629_, _25628_, _04608_);
  nor (_25630_, _12017_, _10403_);
  nor (_25631_, _25630_, _25565_);
  nor (_25632_, _25631_, _04608_);
  or (_25633_, _25632_, _25629_);
  and (_25634_, _25633_, _04606_);
  nor (_25635_, _12015_, _10403_);
  nor (_25636_, _25635_, _25565_);
  nor (_25638_, _25636_, _04606_);
  nor (_25639_, _25638_, _17220_);
  not (_25640_, _25639_);
  nor (_25641_, _25640_, _25634_);
  nor (_25642_, _25641_, _25568_);
  or (_25643_, _25642_, _43231_);
  or (_25644_, _43227_, \oc8051_golden_model_1.PCON [0]);
  and (_25645_, _25644_, _41991_);
  and (_43521_, _25645_, _25643_);
  and (_25646_, _06835_, _05323_);
  not (_25648_, \oc8051_golden_model_1.PCON [1]);
  nor (_25649_, _05323_, _25648_);
  nor (_25650_, _25649_, _05970_);
  not (_25651_, _25650_);
  nor (_25652_, _25651_, _25646_);
  not (_25653_, _25652_);
  and (_25654_, _05323_, _05898_);
  nor (_25655_, _25654_, _25649_);
  and (_25656_, _25655_, _07441_);
  nor (_25657_, _05323_, \oc8051_golden_model_1.PCON [1]);
  and (_25659_, _05323_, _03320_);
  nor (_25660_, _25659_, _25657_);
  and (_25661_, _25660_, _04499_);
  nor (_25662_, _04499_, _25648_);
  or (_25663_, _25662_, _25661_);
  and (_25664_, _25663_, _04515_);
  and (_25665_, _12234_, _05323_);
  nor (_25666_, _25665_, _25657_);
  and (_25667_, _25666_, _03599_);
  or (_25668_, _25667_, _25664_);
  and (_25670_, _25668_, _04524_);
  nor (_25671_, _25655_, _04524_);
  nor (_25672_, _25671_, _25670_);
  nor (_25673_, _25672_, _03603_);
  and (_25674_, _25660_, _03603_);
  nor (_25675_, _25674_, _07441_);
  not (_25676_, _25675_);
  nor (_25677_, _25676_, _25673_);
  nor (_25678_, _25677_, _25656_);
  nor (_25679_, _25678_, _05969_);
  nor (_25681_, _25679_, _03644_);
  and (_25682_, _25681_, _25653_);
  not (_25683_, _25657_);
  and (_25684_, _12330_, _05323_);
  nor (_25685_, _25684_, _03275_);
  and (_25686_, _25685_, _25683_);
  nor (_25687_, _25686_, _25682_);
  nor (_25688_, _25687_, _08861_);
  nor (_25689_, _12220_, _10403_);
  nor (_25690_, _25689_, _04591_);
  and (_25692_, _05323_, _04347_);
  nor (_25693_, _25692_, _04582_);
  nor (_25694_, _25693_, _25690_);
  nor (_25695_, _25694_, _25657_);
  nor (_25696_, _25695_, _25688_);
  nor (_25697_, _25696_, _03778_);
  nor (_25698_, _12347_, _10403_);
  nor (_25699_, _25698_, _04589_);
  and (_25700_, _25699_, _25683_);
  nor (_25701_, _25700_, _25697_);
  nor (_25703_, _25701_, _03655_);
  nor (_25704_, _12219_, _10403_);
  nor (_25705_, _25704_, _04596_);
  and (_25706_, _25705_, _25683_);
  nor (_25707_, _25706_, _25703_);
  nor (_25708_, _25707_, _03773_);
  nor (_25709_, _25649_, _05699_);
  nor (_25710_, _25709_, _04594_);
  and (_25711_, _25710_, _25660_);
  nor (_25712_, _25711_, _25708_);
  or (_25714_, _25712_, _18553_);
  and (_25715_, _25692_, _05698_);
  or (_25716_, _25657_, _04608_);
  or (_25717_, _25716_, _25715_);
  and (_25718_, _25659_, _05698_);
  or (_25719_, _25657_, _04606_);
  or (_25720_, _25719_, _25718_);
  and (_25721_, _25720_, _04260_);
  and (_25722_, _25721_, _25717_);
  and (_25723_, _25722_, _25714_);
  nor (_25724_, _25666_, _04260_);
  nor (_25725_, _25724_, _25723_);
  and (_25726_, _25725_, _03820_);
  nor (_25727_, _25665_, _25649_);
  nor (_25728_, _25727_, _03820_);
  or (_25729_, _25728_, _25726_);
  or (_25730_, _25729_, _43231_);
  or (_25731_, _43227_, \oc8051_golden_model_1.PCON [1]);
  and (_25732_, _25731_, _41991_);
  and (_43522_, _25732_, _25730_);
  not (_25735_, \oc8051_golden_model_1.PCON [2]);
  nor (_25736_, _05323_, _25735_);
  nor (_25737_, _12543_, _10403_);
  nor (_25738_, _25737_, _25736_);
  nor (_25739_, _25738_, _04606_);
  and (_25740_, _06839_, _05323_);
  nor (_25741_, _25740_, _25736_);
  or (_25742_, _25741_, _05970_);
  and (_25743_, _05323_, \oc8051_golden_model_1.ACC [2]);
  nor (_25744_, _25743_, _25736_);
  nor (_25746_, _25744_, _03611_);
  nor (_25747_, _25744_, _04500_);
  nor (_25748_, _04499_, _25735_);
  or (_25749_, _25748_, _25747_);
  and (_25750_, _25749_, _04515_);
  nor (_25751_, _12430_, _10403_);
  nor (_25752_, _25751_, _25736_);
  nor (_25753_, _25752_, _04515_);
  or (_25754_, _25753_, _25750_);
  and (_25755_, _25754_, _04524_);
  nor (_25757_, _10403_, _05130_);
  nor (_25758_, _25757_, _25736_);
  nor (_25759_, _25758_, _04524_);
  nor (_25760_, _25759_, _25755_);
  nor (_25761_, _25760_, _03603_);
  or (_25762_, _25761_, _07441_);
  nor (_25763_, _25762_, _25746_);
  and (_25764_, _25758_, _07441_);
  or (_25765_, _25764_, _05969_);
  or (_25766_, _25765_, _25763_);
  and (_25768_, _25766_, _03275_);
  and (_25769_, _25768_, _25742_);
  nor (_25770_, _12524_, _10403_);
  or (_25771_, _25736_, _03275_);
  nor (_25772_, _25771_, _25770_);
  or (_25773_, _25772_, _03650_);
  nor (_25774_, _25773_, _25769_);
  and (_25775_, _05323_, _06414_);
  nor (_25776_, _25775_, _25736_);
  nand (_25777_, _25776_, _04591_);
  and (_25779_, _25777_, _08861_);
  nor (_25780_, _25779_, _25774_);
  and (_25781_, _12538_, _05323_);
  nor (_25782_, _25781_, _25736_);
  and (_25783_, _25782_, _03649_);
  nor (_25784_, _25783_, _25780_);
  nor (_25785_, _25784_, _03778_);
  and (_25786_, _12544_, _05323_);
  or (_25787_, _25736_, _04589_);
  nor (_25788_, _25787_, _25786_);
  or (_25790_, _25788_, _03655_);
  nor (_25791_, _25790_, _25785_);
  nor (_25792_, _25736_, _05793_);
  not (_25793_, _25792_);
  nor (_25794_, _25776_, _04596_);
  and (_25795_, _25794_, _25793_);
  nor (_25796_, _25795_, _25791_);
  nor (_25797_, _25796_, _03773_);
  nor (_25798_, _25744_, _04594_);
  and (_25799_, _25798_, _25793_);
  nor (_25801_, _25799_, _03653_);
  not (_25802_, _25801_);
  nor (_25803_, _25802_, _25797_);
  nor (_25804_, _12537_, _10403_);
  or (_25805_, _25736_, _04608_);
  nor (_25806_, _25805_, _25804_);
  or (_25807_, _25806_, _03786_);
  nor (_25808_, _25807_, _25803_);
  nor (_25809_, _25808_, _25739_);
  nor (_25810_, _25809_, _03809_);
  nor (_25812_, _25752_, _04260_);
  or (_25813_, _25812_, _03816_);
  nor (_25814_, _25813_, _25810_);
  and (_25815_, _12600_, _05323_);
  or (_25816_, _25736_, _03820_);
  nor (_25817_, _25816_, _25815_);
  nor (_25818_, _25817_, _25814_);
  or (_25819_, _25818_, _43231_);
  or (_25820_, _43227_, \oc8051_golden_model_1.PCON [2]);
  and (_25821_, _25820_, _41991_);
  and (_43523_, _25821_, _25819_);
  not (_25823_, \oc8051_golden_model_1.PCON [3]);
  nor (_25824_, _05323_, _25823_);
  nor (_25825_, _12618_, _10403_);
  nor (_25826_, _25825_, _25824_);
  nor (_25827_, _25826_, _04606_);
  and (_25828_, _05323_, \oc8051_golden_model_1.ACC [3]);
  nor (_25829_, _25828_, _25824_);
  nor (_25830_, _25829_, _04500_);
  nor (_25831_, _04499_, _25823_);
  or (_25833_, _25831_, _25830_);
  and (_25834_, _25833_, _04515_);
  nor (_25835_, _12625_, _10403_);
  nor (_25836_, _25835_, _25824_);
  nor (_25837_, _25836_, _04515_);
  or (_25838_, _25837_, _25834_);
  and (_25839_, _25838_, _04524_);
  nor (_25840_, _10403_, _04944_);
  nor (_25841_, _25840_, _25824_);
  nor (_25842_, _25841_, _04524_);
  nor (_25844_, _25842_, _25839_);
  nor (_25845_, _25844_, _03603_);
  nor (_25846_, _25829_, _03611_);
  nor (_25847_, _25846_, _07441_);
  not (_25848_, _25847_);
  nor (_25849_, _25848_, _25845_);
  and (_25850_, _25841_, _07441_);
  or (_25851_, _25850_, _05969_);
  or (_25852_, _25851_, _25849_);
  and (_25853_, _06838_, _05323_);
  nor (_25855_, _25853_, _25824_);
  or (_25856_, _25855_, _05970_);
  and (_25857_, _25856_, _03275_);
  and (_25858_, _25857_, _25852_);
  nor (_25859_, _12731_, _10403_);
  or (_25860_, _25824_, _03275_);
  nor (_25861_, _25860_, _25859_);
  or (_25862_, _25861_, _03650_);
  nor (_25863_, _25862_, _25858_);
  and (_25864_, _05323_, _06347_);
  nor (_25866_, _25864_, _25824_);
  nand (_25867_, _25866_, _04591_);
  and (_25868_, _25867_, _08861_);
  nor (_25869_, _25868_, _25863_);
  and (_25870_, _12746_, _05323_);
  nor (_25871_, _25870_, _25824_);
  and (_25872_, _25871_, _03649_);
  nor (_25873_, _25872_, _25869_);
  nor (_25874_, _25873_, _03778_);
  and (_25875_, _12619_, _05323_);
  or (_25877_, _25824_, _04589_);
  nor (_25878_, _25877_, _25875_);
  or (_25879_, _25878_, _03655_);
  nor (_25880_, _25879_, _25874_);
  nor (_25881_, _25824_, _05650_);
  not (_25882_, _25881_);
  nor (_25883_, _25866_, _04596_);
  and (_25884_, _25883_, _25882_);
  nor (_25885_, _25884_, _25880_);
  nor (_25886_, _25885_, _03773_);
  nor (_25888_, _25829_, _04594_);
  and (_25889_, _25888_, _25882_);
  or (_25890_, _25889_, _25886_);
  and (_25891_, _25890_, _04608_);
  nor (_25892_, _12745_, _10403_);
  nor (_25893_, _25892_, _25824_);
  nor (_25894_, _25893_, _04608_);
  or (_25895_, _25894_, _25891_);
  and (_25896_, _25895_, _04606_);
  nor (_25897_, _25896_, _25827_);
  nor (_25899_, _25897_, _03809_);
  nor (_25900_, _25836_, _04260_);
  or (_25901_, _25900_, _03816_);
  nor (_25902_, _25901_, _25899_);
  and (_25903_, _12806_, _05323_);
  nor (_25904_, _25903_, _25824_);
  and (_25905_, _25904_, _03816_);
  nor (_25906_, _25905_, _25902_);
  or (_25907_, _25906_, _43231_);
  or (_25908_, _43227_, \oc8051_golden_model_1.PCON [3]);
  and (_25910_, _25908_, _41991_);
  and (_43524_, _25910_, _25907_);
  not (_25911_, \oc8051_golden_model_1.PCON [4]);
  nor (_25912_, _05323_, _25911_);
  nor (_25913_, _12956_, _10403_);
  nor (_25914_, _25913_, _25912_);
  nor (_25915_, _25914_, _04606_);
  and (_25916_, _12957_, _05323_);
  nor (_25917_, _25916_, _25912_);
  nor (_25918_, _25917_, _04589_);
  and (_25920_, _06375_, _05323_);
  nor (_25921_, _25920_, _25912_);
  and (_25922_, _25921_, _03650_);
  and (_25923_, _05323_, \oc8051_golden_model_1.ACC [4]);
  nor (_25924_, _25923_, _25912_);
  nor (_25925_, _25924_, _03611_);
  nor (_25926_, _25924_, _04500_);
  nor (_25927_, _04499_, _25911_);
  or (_25928_, _25927_, _25926_);
  and (_25929_, _25928_, _04515_);
  nor (_25931_, _12820_, _10403_);
  nor (_25932_, _25931_, _25912_);
  nor (_25933_, _25932_, _04515_);
  or (_25934_, _25933_, _25929_);
  and (_25935_, _25934_, _04524_);
  nor (_25936_, _05840_, _10403_);
  nor (_25937_, _25936_, _25912_);
  nor (_25938_, _25937_, _04524_);
  nor (_25939_, _25938_, _25935_);
  nor (_25940_, _25939_, _03603_);
  or (_25942_, _25940_, _07441_);
  nor (_25943_, _25942_, _25925_);
  and (_25944_, _25937_, _07441_);
  nor (_25945_, _25944_, _25943_);
  nor (_25946_, _25945_, _05969_);
  and (_25947_, _06843_, _05323_);
  nor (_25948_, _25912_, _05970_);
  not (_25949_, _25948_);
  nor (_25950_, _25949_, _25947_);
  or (_25951_, _25950_, _03644_);
  nor (_25953_, _25951_, _25946_);
  nor (_25954_, _12936_, _10403_);
  nor (_25955_, _25954_, _25912_);
  nor (_25956_, _25955_, _03275_);
  or (_25957_, _25956_, _03650_);
  nor (_25958_, _25957_, _25953_);
  nor (_25959_, _25958_, _25922_);
  or (_25960_, _25959_, _03649_);
  and (_25961_, _12951_, _05323_);
  or (_25962_, _25961_, _25912_);
  or (_25964_, _25962_, _04591_);
  and (_25965_, _25964_, _04589_);
  and (_25966_, _25965_, _25960_);
  nor (_25967_, _25966_, _25918_);
  nor (_25968_, _25967_, _03655_);
  nor (_25969_, _25912_, _05889_);
  not (_25970_, _25969_);
  nor (_25971_, _25921_, _04596_);
  and (_25972_, _25971_, _25970_);
  nor (_25973_, _25972_, _25968_);
  nor (_25975_, _25973_, _03773_);
  nor (_25976_, _25924_, _04594_);
  and (_25977_, _25976_, _25970_);
  or (_25978_, _25977_, _25975_);
  and (_25979_, _25978_, _04608_);
  nor (_25980_, _12949_, _10403_);
  nor (_25981_, _25980_, _25912_);
  nor (_25982_, _25981_, _04608_);
  or (_25983_, _25982_, _25979_);
  and (_25984_, _25983_, _04606_);
  nor (_25986_, _25984_, _25915_);
  nor (_25987_, _25986_, _03809_);
  nor (_25988_, _25932_, _04260_);
  or (_25989_, _25988_, _03816_);
  nor (_25990_, _25989_, _25987_);
  and (_25991_, _13013_, _05323_);
  or (_25992_, _25912_, _03820_);
  nor (_25993_, _25992_, _25991_);
  nor (_25994_, _25993_, _25990_);
  or (_25995_, _25994_, _43231_);
  or (_25997_, _43227_, \oc8051_golden_model_1.PCON [4]);
  and (_25998_, _25997_, _41991_);
  and (_43525_, _25998_, _25995_);
  not (_25999_, \oc8051_golden_model_1.PCON [5]);
  nor (_26000_, _05323_, _25999_);
  nor (_26001_, _13159_, _10403_);
  nor (_26002_, _26001_, _26000_);
  nor (_26003_, _26002_, _04606_);
  and (_26004_, _13160_, _05323_);
  nor (_26005_, _26004_, _26000_);
  nor (_26007_, _26005_, _04589_);
  and (_26008_, _06842_, _05323_);
  or (_26009_, _26008_, _26000_);
  and (_26010_, _26009_, _05969_);
  and (_26011_, _05323_, \oc8051_golden_model_1.ACC [5]);
  nor (_26012_, _26011_, _26000_);
  nor (_26013_, _26012_, _03611_);
  nor (_26014_, _26012_, _04500_);
  nor (_26015_, _04499_, _25999_);
  or (_26016_, _26015_, _26014_);
  and (_26018_, _26016_, _04515_);
  nor (_26019_, _13035_, _10403_);
  nor (_26020_, _26019_, _26000_);
  nor (_26021_, _26020_, _04515_);
  or (_26022_, _26021_, _26018_);
  and (_26023_, _26022_, _04524_);
  nor (_26024_, _05552_, _10403_);
  nor (_26025_, _26024_, _26000_);
  nor (_26026_, _26025_, _04524_);
  nor (_26027_, _26026_, _26023_);
  nor (_26029_, _26027_, _03603_);
  or (_26030_, _26029_, _07441_);
  nor (_26031_, _26030_, _26013_);
  and (_26032_, _26025_, _07441_);
  or (_26033_, _26032_, _05969_);
  nor (_26034_, _26033_, _26031_);
  or (_26035_, _26034_, _26010_);
  and (_26036_, _26035_, _03275_);
  nor (_26037_, _13139_, _10403_);
  nor (_26038_, _26037_, _26000_);
  nor (_26040_, _26038_, _03275_);
  or (_26041_, _26040_, _08861_);
  or (_26042_, _26041_, _26036_);
  and (_26043_, _13154_, _05323_);
  or (_26044_, _26000_, _04591_);
  or (_26045_, _26044_, _26043_);
  and (_26046_, _06358_, _05323_);
  nor (_26047_, _26046_, _26000_);
  and (_26048_, _26047_, _03650_);
  nor (_26049_, _26048_, _03778_);
  and (_26051_, _26049_, _26045_);
  and (_26052_, _26051_, _26042_);
  nor (_26053_, _26052_, _26007_);
  nor (_26054_, _26053_, _03655_);
  nor (_26055_, _26000_, _05601_);
  not (_26056_, _26055_);
  nor (_26057_, _26047_, _04596_);
  and (_26058_, _26057_, _26056_);
  nor (_26059_, _26058_, _26054_);
  nor (_26060_, _26059_, _03773_);
  nor (_26062_, _26012_, _04594_);
  and (_26063_, _26062_, _26056_);
  nor (_26064_, _26063_, _03653_);
  not (_26065_, _26064_);
  nor (_26066_, _26065_, _26060_);
  nor (_26067_, _13152_, _10403_);
  or (_26068_, _26000_, _04608_);
  nor (_26069_, _26068_, _26067_);
  or (_26070_, _26069_, _03786_);
  nor (_26071_, _26070_, _26066_);
  nor (_26072_, _26071_, _26003_);
  nor (_26073_, _26072_, _03809_);
  nor (_26074_, _26020_, _04260_);
  or (_26075_, _26074_, _03816_);
  nor (_26076_, _26075_, _26073_);
  and (_26077_, _13217_, _05323_);
  or (_26078_, _26000_, _03820_);
  nor (_26079_, _26078_, _26077_);
  nor (_26080_, _26079_, _26076_);
  or (_26081_, _26080_, _43231_);
  or (_26084_, _43227_, \oc8051_golden_model_1.PCON [5]);
  and (_26085_, _26084_, _41991_);
  and (_43526_, _26085_, _26081_);
  not (_26086_, \oc8051_golden_model_1.PCON [6]);
  nor (_26087_, _05323_, _26086_);
  nor (_26088_, _13373_, _10403_);
  nor (_26089_, _26088_, _26087_);
  nor (_26090_, _26089_, _04606_);
  and (_26091_, _13374_, _05323_);
  nor (_26092_, _26091_, _26087_);
  nor (_26094_, _26092_, _04589_);
  and (_26095_, _06531_, _05323_);
  or (_26096_, _26095_, _26087_);
  and (_26097_, _26096_, _05969_);
  and (_26098_, _05323_, \oc8051_golden_model_1.ACC [6]);
  nor (_26099_, _26098_, _26087_);
  nor (_26100_, _26099_, _04500_);
  nor (_26101_, _04499_, _26086_);
  or (_26102_, _26101_, _26100_);
  and (_26103_, _26102_, _04515_);
  nor (_26105_, _13235_, _10403_);
  nor (_26106_, _26105_, _26087_);
  nor (_26107_, _26106_, _04515_);
  or (_26108_, _26107_, _26103_);
  and (_26109_, _26108_, _04524_);
  nor (_26110_, _05442_, _10403_);
  nor (_26111_, _26110_, _26087_);
  nor (_26112_, _26111_, _04524_);
  nor (_26113_, _26112_, _26109_);
  nor (_26114_, _26113_, _03603_);
  nor (_26116_, _26099_, _03611_);
  nor (_26117_, _26116_, _07441_);
  not (_26118_, _26117_);
  nor (_26119_, _26118_, _26114_);
  and (_26120_, _26111_, _07441_);
  or (_26121_, _26120_, _05969_);
  nor (_26122_, _26121_, _26119_);
  or (_26123_, _26122_, _26097_);
  and (_26124_, _26123_, _03275_);
  nor (_26125_, _13356_, _10403_);
  nor (_26127_, _26125_, _26087_);
  nor (_26128_, _26127_, _03275_);
  or (_26129_, _26128_, _08861_);
  or (_26130_, _26129_, _26124_);
  and (_26131_, _13245_, _05323_);
  or (_26132_, _26087_, _04591_);
  or (_26133_, _26132_, _26131_);
  and (_26134_, _13363_, _05323_);
  nor (_26135_, _26134_, _26087_);
  and (_26136_, _26135_, _03650_);
  nor (_26138_, _26136_, _03778_);
  and (_26139_, _26138_, _26133_);
  and (_26140_, _26139_, _26130_);
  nor (_26141_, _26140_, _26094_);
  nor (_26142_, _26141_, _03655_);
  nor (_26143_, _26087_, _05491_);
  not (_26144_, _26143_);
  nor (_26145_, _26135_, _04596_);
  and (_26146_, _26145_, _26144_);
  nor (_26147_, _26146_, _26142_);
  nor (_26149_, _26147_, _03773_);
  nor (_26150_, _26099_, _04594_);
  and (_26151_, _26150_, _26144_);
  or (_26152_, _26151_, _26149_);
  and (_26153_, _26152_, _04608_);
  nor (_26154_, _13243_, _10403_);
  nor (_26155_, _26154_, _26087_);
  nor (_26156_, _26155_, _04608_);
  or (_26157_, _26156_, _26153_);
  and (_26158_, _26157_, _04606_);
  nor (_26160_, _26158_, _26090_);
  nor (_26161_, _26160_, _03809_);
  nor (_26162_, _26106_, _04260_);
  or (_26163_, _26162_, _03816_);
  nor (_26164_, _26163_, _26161_);
  and (_26165_, _13425_, _05323_);
  or (_26166_, _26087_, _03820_);
  nor (_26167_, _26166_, _26165_);
  nor (_26168_, _26167_, _26164_);
  or (_26169_, _26168_, _43231_);
  or (_26171_, _43227_, \oc8051_golden_model_1.PCON [6]);
  and (_26172_, _26171_, _41991_);
  and (_43527_, _26172_, _26169_);
  not (_26173_, \oc8051_golden_model_1.SBUF [0]);
  nor (_26174_, _05330_, _26173_);
  nor (_26175_, _05744_, _10485_);
  nor (_26176_, _26175_, _26174_);
  and (_26177_, _26176_, _17220_);
  and (_26178_, _05330_, \oc8051_golden_model_1.ACC [0]);
  nor (_26179_, _26178_, _26174_);
  nor (_26180_, _26179_, _03611_);
  nor (_26181_, _26180_, _07441_);
  nor (_26182_, _26176_, _04515_);
  nor (_26183_, _04499_, _26173_);
  nor (_26184_, _26179_, _04500_);
  nor (_26185_, _26184_, _26183_);
  nor (_26186_, _26185_, _03599_);
  or (_26187_, _26186_, _03597_);
  nor (_26188_, _26187_, _26182_);
  or (_26189_, _26188_, _03603_);
  and (_26192_, _26189_, _26181_);
  and (_26193_, _05330_, _04491_);
  and (_26194_, _06889_, _04524_);
  or (_26195_, _26194_, _26174_);
  nor (_26196_, _26195_, _26193_);
  nor (_26197_, _26196_, _26192_);
  nor (_26198_, _26197_, _05969_);
  and (_26199_, _06836_, _05330_);
  nor (_26200_, _26174_, _05970_);
  not (_26201_, _26200_);
  nor (_26203_, _26201_, _26199_);
  nor (_26204_, _26203_, _26198_);
  nor (_26205_, _26204_, _03644_);
  nor (_26206_, _12129_, _10485_);
  or (_26207_, _26174_, _03275_);
  nor (_26208_, _26207_, _26206_);
  or (_26209_, _26208_, _03650_);
  nor (_26210_, _26209_, _26205_);
  and (_26211_, _05330_, _06366_);
  nor (_26212_, _26211_, _26174_);
  nand (_26214_, _26212_, _04591_);
  and (_26215_, _26214_, _08861_);
  nor (_26216_, _26215_, _26210_);
  and (_26217_, _12019_, _05330_);
  nor (_26218_, _26217_, _26174_);
  and (_26219_, _26218_, _03649_);
  nor (_26220_, _26219_, _26216_);
  nor (_26221_, _26220_, _03778_);
  and (_26222_, _12145_, _05330_);
  or (_26223_, _26174_, _04589_);
  nor (_26225_, _26223_, _26222_);
  or (_26226_, _26225_, _03655_);
  nor (_26227_, _26226_, _26221_);
  or (_26228_, _26212_, _04596_);
  nor (_26229_, _26228_, _26175_);
  nor (_26230_, _26229_, _26227_);
  nor (_26231_, _26230_, _03773_);
  nor (_26232_, _26174_, _05744_);
  or (_26233_, _26232_, _04594_);
  nor (_26234_, _26233_, _26179_);
  or (_26236_, _26234_, _26231_);
  and (_26237_, _26236_, _04608_);
  nor (_26238_, _12017_, _10485_);
  nor (_26239_, _26238_, _26174_);
  nor (_26240_, _26239_, _04608_);
  or (_26241_, _26240_, _26237_);
  and (_26242_, _26241_, _04606_);
  nor (_26243_, _12015_, _10485_);
  nor (_26244_, _26243_, _26174_);
  nor (_26245_, _26244_, _04606_);
  nor (_26247_, _26245_, _17220_);
  not (_26248_, _26247_);
  nor (_26249_, _26248_, _26242_);
  nor (_26250_, _26249_, _26177_);
  or (_26251_, _26250_, _43231_);
  or (_26252_, _43227_, \oc8051_golden_model_1.SBUF [0]);
  and (_26253_, _26252_, _41991_);
  and (_43530_, _26253_, _26251_);
  and (_26254_, _06835_, _05330_);
  not (_26255_, \oc8051_golden_model_1.SBUF [1]);
  nor (_26257_, _05330_, _26255_);
  nor (_26258_, _26257_, _05970_);
  not (_26259_, _26258_);
  nor (_26260_, _26259_, _26254_);
  not (_26261_, _26260_);
  and (_26262_, _05330_, _05898_);
  nor (_26263_, _26262_, _26257_);
  and (_26264_, _26263_, _07441_);
  nor (_26265_, _05330_, \oc8051_golden_model_1.SBUF [1]);
  and (_26266_, _05330_, _03320_);
  nor (_26268_, _26266_, _26265_);
  and (_26269_, _26268_, _04499_);
  nor (_26270_, _04499_, _26255_);
  or (_26271_, _26270_, _26269_);
  and (_26272_, _26271_, _04515_);
  and (_26273_, _12234_, _05330_);
  nor (_26274_, _26273_, _26265_);
  and (_26275_, _26274_, _03599_);
  or (_26276_, _26275_, _26272_);
  and (_26277_, _26276_, _04524_);
  nor (_26279_, _26263_, _04524_);
  nor (_26280_, _26279_, _26277_);
  nor (_26281_, _26280_, _03603_);
  and (_26282_, _26268_, _03603_);
  nor (_26283_, _26282_, _07441_);
  not (_26284_, _26283_);
  nor (_26285_, _26284_, _26281_);
  nor (_26286_, _26285_, _26264_);
  nor (_26287_, _26286_, _05969_);
  nor (_26288_, _26287_, _03644_);
  and (_26290_, _26288_, _26261_);
  not (_26291_, _26265_);
  and (_26292_, _12330_, _05330_);
  nor (_26293_, _26292_, _03275_);
  and (_26294_, _26293_, _26291_);
  nor (_26295_, _26294_, _26290_);
  nor (_26296_, _26295_, _08861_);
  nor (_26297_, _12220_, _10485_);
  nor (_26298_, _26297_, _04591_);
  and (_26299_, _05330_, _04347_);
  nor (_26301_, _26299_, _04582_);
  or (_26302_, _26301_, _26298_);
  and (_26303_, _26302_, _26291_);
  nor (_26304_, _26303_, _26296_);
  nor (_26305_, _26304_, _03778_);
  nor (_26306_, _12347_, _10485_);
  nor (_26307_, _26306_, _04589_);
  and (_26308_, _26307_, _26291_);
  nor (_26309_, _26308_, _26305_);
  nor (_26310_, _26309_, _03655_);
  nor (_26312_, _12219_, _10485_);
  nor (_26313_, _26312_, _04596_);
  and (_26314_, _26313_, _26291_);
  nor (_26315_, _26314_, _26310_);
  nor (_26316_, _26315_, _03773_);
  nor (_26317_, _26257_, _05699_);
  nor (_26318_, _26317_, _04594_);
  and (_26319_, _26318_, _26268_);
  nor (_26320_, _26319_, _26316_);
  or (_26321_, _26320_, _18553_);
  and (_26323_, _26299_, _05698_);
  nor (_26324_, _26323_, _04608_);
  and (_26325_, _26324_, _26291_);
  nand (_26326_, _26266_, _05698_);
  nor (_26327_, _26265_, _04606_);
  and (_26328_, _26327_, _26326_);
  or (_26329_, _26328_, _03809_);
  nor (_26330_, _26329_, _26325_);
  and (_26331_, _26330_, _26321_);
  nor (_26332_, _26274_, _04260_);
  nor (_26334_, _26332_, _26331_);
  and (_26335_, _26334_, _03820_);
  nor (_26336_, _26273_, _26257_);
  nor (_26337_, _26336_, _03820_);
  or (_26338_, _26337_, _26335_);
  or (_26339_, _26338_, _43231_);
  or (_26340_, _43227_, \oc8051_golden_model_1.SBUF [1]);
  and (_26341_, _26340_, _41991_);
  and (_43531_, _26341_, _26339_);
  not (_26342_, \oc8051_golden_model_1.SBUF [2]);
  nor (_26344_, _05330_, _26342_);
  nor (_26345_, _12543_, _10485_);
  nor (_26346_, _26345_, _26344_);
  nor (_26347_, _26346_, _04606_);
  nor (_26348_, _10485_, _05130_);
  nor (_26349_, _26348_, _26344_);
  and (_26350_, _26349_, _07441_);
  nor (_26351_, _12430_, _10485_);
  nor (_26352_, _26351_, _26344_);
  nor (_26353_, _26352_, _04515_);
  nor (_26355_, _04499_, _26342_);
  and (_26356_, _05330_, \oc8051_golden_model_1.ACC [2]);
  nor (_26357_, _26356_, _26344_);
  nor (_26358_, _26357_, _04500_);
  nor (_26359_, _26358_, _26355_);
  nor (_26360_, _26359_, _03599_);
  or (_26361_, _26360_, _26353_);
  and (_26362_, _26361_, _04524_);
  nor (_26363_, _26349_, _04524_);
  or (_26364_, _26363_, _26362_);
  and (_26366_, _26364_, _03611_);
  nor (_26367_, _26357_, _03611_);
  nor (_26368_, _26367_, _07441_);
  not (_26369_, _26368_);
  nor (_26370_, _26369_, _26366_);
  nor (_26371_, _26370_, _26350_);
  nor (_26372_, _26371_, _05969_);
  and (_26373_, _06839_, _05330_);
  nor (_26374_, _26344_, _05970_);
  not (_26375_, _26374_);
  nor (_26377_, _26375_, _26373_);
  nor (_26378_, _26377_, _26372_);
  nor (_26379_, _26378_, _03644_);
  nor (_26380_, _12524_, _10485_);
  or (_26381_, _26344_, _03275_);
  nor (_26382_, _26381_, _26380_);
  or (_26383_, _26382_, _03650_);
  nor (_26384_, _26383_, _26379_);
  and (_26385_, _05330_, _06414_);
  nor (_26386_, _26385_, _26344_);
  nand (_26388_, _26386_, _04591_);
  and (_26389_, _26388_, _08861_);
  nor (_26390_, _26389_, _26384_);
  and (_26391_, _12538_, _05330_);
  nor (_26392_, _26391_, _26344_);
  and (_26393_, _26392_, _03649_);
  nor (_26394_, _26393_, _26390_);
  nor (_26395_, _26394_, _03778_);
  and (_26396_, _12544_, _05330_);
  or (_26397_, _26344_, _04589_);
  nor (_26399_, _26397_, _26396_);
  or (_26400_, _26399_, _03655_);
  nor (_26401_, _26400_, _26395_);
  nor (_26402_, _26344_, _05793_);
  not (_26403_, _26402_);
  nor (_26404_, _26386_, _04596_);
  and (_26405_, _26404_, _26403_);
  nor (_26406_, _26405_, _26401_);
  nor (_26407_, _26406_, _03773_);
  nor (_26408_, _26357_, _04594_);
  and (_26410_, _26408_, _26403_);
  nor (_26411_, _26410_, _03653_);
  not (_26412_, _26411_);
  nor (_26413_, _26412_, _26407_);
  nor (_26414_, _12537_, _10485_);
  or (_26415_, _26344_, _04608_);
  nor (_26416_, _26415_, _26414_);
  or (_26417_, _26416_, _03786_);
  nor (_26418_, _26417_, _26413_);
  nor (_26419_, _26418_, _26347_);
  nor (_26421_, _26419_, _03809_);
  nor (_26422_, _26352_, _04260_);
  or (_26423_, _26422_, _03816_);
  nor (_26424_, _26423_, _26421_);
  and (_26425_, _12600_, _05330_);
  or (_26426_, _26344_, _03820_);
  nor (_26427_, _26426_, _26425_);
  nor (_26428_, _26427_, _26424_);
  or (_26429_, _26428_, _43231_);
  or (_26430_, _43227_, \oc8051_golden_model_1.SBUF [2]);
  and (_26432_, _26430_, _41991_);
  and (_43532_, _26432_, _26429_);
  not (_26433_, \oc8051_golden_model_1.SBUF [3]);
  nor (_26434_, _05330_, _26433_);
  nor (_26435_, _12618_, _10485_);
  nor (_26436_, _26435_, _26434_);
  nor (_26437_, _26436_, _04606_);
  and (_26438_, _12619_, _05330_);
  nor (_26439_, _26438_, _26434_);
  nor (_26440_, _26439_, _04589_);
  and (_26442_, _06838_, _05330_);
  or (_26443_, _26442_, _26434_);
  and (_26444_, _26443_, _05969_);
  and (_26445_, _05330_, \oc8051_golden_model_1.ACC [3]);
  nor (_26446_, _26445_, _26434_);
  nor (_26447_, _26446_, _03611_);
  nor (_26448_, _26446_, _04500_);
  nor (_26449_, _04499_, _26433_);
  or (_26450_, _26449_, _26448_);
  and (_26451_, _26450_, _04515_);
  nor (_26453_, _12625_, _10485_);
  nor (_26454_, _26453_, _26434_);
  nor (_26455_, _26454_, _04515_);
  or (_26456_, _26455_, _26451_);
  and (_26457_, _26456_, _04524_);
  nor (_26458_, _10485_, _04944_);
  nor (_26459_, _26458_, _26434_);
  nor (_26460_, _26459_, _04524_);
  nor (_26461_, _26460_, _26457_);
  nor (_26462_, _26461_, _03603_);
  or (_26464_, _26462_, _07441_);
  nor (_26465_, _26464_, _26447_);
  and (_26466_, _26459_, _07441_);
  or (_26467_, _26466_, _05969_);
  nor (_26468_, _26467_, _26465_);
  or (_26469_, _26468_, _26444_);
  and (_26470_, _26469_, _03275_);
  nor (_26471_, _12731_, _10485_);
  nor (_26472_, _26471_, _26434_);
  nor (_26473_, _26472_, _03275_);
  or (_26475_, _26473_, _08861_);
  or (_26476_, _26475_, _26470_);
  and (_26477_, _12746_, _05330_);
  or (_26478_, _26434_, _04591_);
  or (_26479_, _26478_, _26477_);
  and (_26480_, _05330_, _06347_);
  nor (_26481_, _26480_, _26434_);
  and (_26482_, _26481_, _03650_);
  nor (_26483_, _26482_, _03778_);
  and (_26484_, _26483_, _26479_);
  and (_26486_, _26484_, _26476_);
  nor (_26487_, _26486_, _26440_);
  nor (_26488_, _26487_, _03655_);
  nor (_26489_, _26434_, _05650_);
  not (_26490_, _26489_);
  nor (_26491_, _26481_, _04596_);
  and (_26492_, _26491_, _26490_);
  nor (_26493_, _26492_, _26488_);
  nor (_26494_, _26493_, _03773_);
  nor (_26495_, _26446_, _04594_);
  and (_26497_, _26495_, _26490_);
  nor (_26498_, _26497_, _03653_);
  not (_26499_, _26498_);
  nor (_26500_, _26499_, _26494_);
  nor (_26501_, _12745_, _10485_);
  or (_26502_, _26434_, _04608_);
  nor (_26503_, _26502_, _26501_);
  or (_26504_, _26503_, _03786_);
  nor (_26505_, _26504_, _26500_);
  nor (_26506_, _26505_, _26437_);
  nor (_26508_, _26506_, _03809_);
  nor (_26509_, _26454_, _04260_);
  or (_26510_, _26509_, _03816_);
  nor (_26511_, _26510_, _26508_);
  and (_26512_, _12806_, _05330_);
  or (_26513_, _26434_, _03820_);
  nor (_26514_, _26513_, _26512_);
  nor (_26515_, _26514_, _26511_);
  or (_26516_, _26515_, _43231_);
  or (_26517_, _43227_, \oc8051_golden_model_1.SBUF [3]);
  and (_26519_, _26517_, _41991_);
  and (_43533_, _26519_, _26516_);
  not (_26520_, \oc8051_golden_model_1.SBUF [4]);
  nor (_26521_, _05330_, _26520_);
  nor (_26522_, _12956_, _10485_);
  nor (_26523_, _26522_, _26521_);
  nor (_26524_, _26523_, _04606_);
  and (_26525_, _12957_, _05330_);
  nor (_26526_, _26525_, _26521_);
  nor (_26527_, _26526_, _04589_);
  and (_26529_, _06375_, _05330_);
  nor (_26530_, _26529_, _26521_);
  and (_26531_, _26530_, _03650_);
  and (_26532_, _05330_, \oc8051_golden_model_1.ACC [4]);
  nor (_26533_, _26532_, _26521_);
  nor (_26534_, _26533_, _03611_);
  nor (_26535_, _26533_, _04500_);
  nor (_26536_, _04499_, _26520_);
  or (_26537_, _26536_, _26535_);
  and (_26538_, _26537_, _04515_);
  nor (_26540_, _12820_, _10485_);
  nor (_26541_, _26540_, _26521_);
  nor (_26542_, _26541_, _04515_);
  or (_26543_, _26542_, _26538_);
  and (_26544_, _26543_, _04524_);
  nor (_26545_, _05840_, _10485_);
  nor (_26546_, _26545_, _26521_);
  nor (_26547_, _26546_, _04524_);
  nor (_26548_, _26547_, _26544_);
  nor (_26549_, _26548_, _03603_);
  or (_26551_, _26549_, _07441_);
  nor (_26552_, _26551_, _26534_);
  and (_26553_, _26546_, _07441_);
  nor (_26554_, _26553_, _26552_);
  nor (_26555_, _26554_, _05969_);
  and (_26556_, _06843_, _05330_);
  nor (_26557_, _26521_, _05970_);
  not (_26558_, _26557_);
  nor (_26559_, _26558_, _26556_);
  or (_26560_, _26559_, _03644_);
  nor (_26562_, _26560_, _26555_);
  nor (_26563_, _12936_, _10485_);
  nor (_26564_, _26563_, _26521_);
  nor (_26565_, _26564_, _03275_);
  or (_26566_, _26565_, _03650_);
  nor (_26567_, _26566_, _26562_);
  nor (_26568_, _26567_, _26531_);
  or (_26569_, _26568_, _03649_);
  and (_26570_, _12951_, _05330_);
  or (_26571_, _26570_, _26521_);
  or (_26573_, _26571_, _04591_);
  and (_26574_, _26573_, _04589_);
  and (_26575_, _26574_, _26569_);
  nor (_26576_, _26575_, _26527_);
  nor (_26577_, _26576_, _03655_);
  nor (_26578_, _26521_, _05889_);
  not (_26579_, _26578_);
  nor (_26580_, _26530_, _04596_);
  and (_26581_, _26580_, _26579_);
  nor (_26582_, _26581_, _26577_);
  nor (_26584_, _26582_, _03773_);
  nor (_26585_, _26533_, _04594_);
  and (_26586_, _26585_, _26579_);
  nor (_26587_, _26586_, _03653_);
  not (_26588_, _26587_);
  nor (_26589_, _26588_, _26584_);
  nor (_26590_, _12949_, _10485_);
  or (_26591_, _26521_, _04608_);
  nor (_26592_, _26591_, _26590_);
  or (_26593_, _26592_, _03786_);
  nor (_26595_, _26593_, _26589_);
  nor (_26596_, _26595_, _26524_);
  nor (_26597_, _26596_, _03809_);
  nor (_26598_, _26541_, _04260_);
  or (_26599_, _26598_, _03816_);
  nor (_26600_, _26599_, _26597_);
  and (_26601_, _13013_, _05330_);
  or (_26602_, _26521_, _03820_);
  nor (_26603_, _26602_, _26601_);
  nor (_26604_, _26603_, _26600_);
  or (_26606_, _26604_, _43231_);
  or (_26607_, _43227_, \oc8051_golden_model_1.SBUF [4]);
  and (_26608_, _26607_, _41991_);
  and (_43534_, _26608_, _26606_);
  not (_26609_, \oc8051_golden_model_1.SBUF [5]);
  nor (_26610_, _05330_, _26609_);
  nor (_26611_, _13159_, _10485_);
  nor (_26612_, _26611_, _26610_);
  nor (_26613_, _26612_, _04606_);
  and (_26614_, _13160_, _05330_);
  nor (_26616_, _26614_, _26610_);
  nor (_26617_, _26616_, _04589_);
  and (_26618_, _06842_, _05330_);
  or (_26619_, _26618_, _26610_);
  and (_26620_, _26619_, _05969_);
  and (_26621_, _05330_, \oc8051_golden_model_1.ACC [5]);
  nor (_26622_, _26621_, _26610_);
  nor (_26623_, _26622_, _04500_);
  nor (_26624_, _04499_, _26609_);
  or (_26625_, _26624_, _26623_);
  and (_26626_, _26625_, _04515_);
  nor (_26627_, _13035_, _10485_);
  nor (_26628_, _26627_, _26610_);
  nor (_26629_, _26628_, _04515_);
  or (_26630_, _26629_, _26626_);
  and (_26631_, _26630_, _04524_);
  nor (_26632_, _05552_, _10485_);
  nor (_26633_, _26632_, _26610_);
  nor (_26634_, _26633_, _04524_);
  nor (_26635_, _26634_, _26631_);
  nor (_26638_, _26635_, _03603_);
  nor (_26639_, _26622_, _03611_);
  nor (_26640_, _26639_, _07441_);
  not (_26641_, _26640_);
  nor (_26642_, _26641_, _26638_);
  and (_26643_, _26633_, _07441_);
  or (_26644_, _26643_, _05969_);
  nor (_26645_, _26644_, _26642_);
  or (_26646_, _26645_, _26620_);
  and (_26647_, _26646_, _03275_);
  nor (_26649_, _13139_, _10485_);
  nor (_26650_, _26649_, _26610_);
  nor (_26651_, _26650_, _03275_);
  or (_26652_, _26651_, _08861_);
  or (_26653_, _26652_, _26647_);
  and (_26654_, _13154_, _05330_);
  or (_26655_, _26610_, _04591_);
  or (_26656_, _26655_, _26654_);
  and (_26657_, _06358_, _05330_);
  nor (_26658_, _26657_, _26610_);
  and (_26660_, _26658_, _03650_);
  nor (_26661_, _26660_, _03778_);
  and (_26662_, _26661_, _26656_);
  and (_26663_, _26662_, _26653_);
  nor (_26664_, _26663_, _26617_);
  nor (_26665_, _26664_, _03655_);
  nor (_26666_, _26610_, _05601_);
  not (_26667_, _26666_);
  nor (_26668_, _26658_, _04596_);
  and (_26669_, _26668_, _26667_);
  nor (_26671_, _26669_, _26665_);
  nor (_26672_, _26671_, _03773_);
  nor (_26673_, _26622_, _04594_);
  and (_26674_, _26673_, _26667_);
  nor (_26675_, _26674_, _03653_);
  not (_26676_, _26675_);
  nor (_26677_, _26676_, _26672_);
  nor (_26678_, _13152_, _10485_);
  or (_26679_, _26610_, _04608_);
  nor (_26680_, _26679_, _26678_);
  or (_26682_, _26680_, _03786_);
  nor (_26683_, _26682_, _26677_);
  nor (_26684_, _26683_, _26613_);
  nor (_26685_, _26684_, _03809_);
  nor (_26686_, _26628_, _04260_);
  or (_26687_, _26686_, _03816_);
  nor (_26688_, _26687_, _26685_);
  and (_26689_, _13217_, _05330_);
  or (_26690_, _26610_, _03820_);
  nor (_26691_, _26690_, _26689_);
  nor (_26693_, _26691_, _26688_);
  or (_26694_, _26693_, _43231_);
  or (_26695_, _43227_, \oc8051_golden_model_1.SBUF [5]);
  and (_26696_, _26695_, _41991_);
  and (_43535_, _26696_, _26694_);
  not (_26697_, \oc8051_golden_model_1.SBUF [6]);
  nor (_26698_, _05330_, _26697_);
  nor (_26699_, _13373_, _10485_);
  nor (_26700_, _26699_, _26698_);
  nor (_26701_, _26700_, _04606_);
  and (_26703_, _13374_, _05330_);
  nor (_26704_, _26703_, _26698_);
  nor (_26705_, _26704_, _04589_);
  and (_26706_, _06531_, _05330_);
  or (_26707_, _26706_, _26698_);
  and (_26708_, _26707_, _05969_);
  and (_26709_, _05330_, \oc8051_golden_model_1.ACC [6]);
  nor (_26710_, _26709_, _26698_);
  nor (_26711_, _26710_, _03611_);
  nor (_26712_, _26710_, _04500_);
  nor (_26714_, _04499_, _26697_);
  or (_26715_, _26714_, _26712_);
  and (_26716_, _26715_, _04515_);
  nor (_26717_, _13235_, _10485_);
  nor (_26718_, _26717_, _26698_);
  nor (_26719_, _26718_, _04515_);
  or (_26720_, _26719_, _26716_);
  and (_26721_, _26720_, _04524_);
  nor (_26722_, _05442_, _10485_);
  nor (_26723_, _26722_, _26698_);
  nor (_26725_, _26723_, _04524_);
  nor (_26726_, _26725_, _26721_);
  nor (_26727_, _26726_, _03603_);
  or (_26728_, _26727_, _07441_);
  nor (_26729_, _26728_, _26711_);
  and (_26730_, _26723_, _07441_);
  or (_26731_, _26730_, _05969_);
  nor (_26732_, _26731_, _26729_);
  or (_26733_, _26732_, _26708_);
  and (_26734_, _26733_, _03275_);
  nor (_26736_, _13356_, _10485_);
  nor (_26737_, _26736_, _26698_);
  nor (_26738_, _26737_, _03275_);
  or (_26739_, _26738_, _08861_);
  or (_26740_, _26739_, _26734_);
  and (_26741_, _13245_, _05330_);
  or (_26742_, _26698_, _04591_);
  or (_26743_, _26742_, _26741_);
  and (_26744_, _13363_, _05330_);
  nor (_26745_, _26744_, _26698_);
  and (_26747_, _26745_, _03650_);
  nor (_26748_, _26747_, _03778_);
  and (_26749_, _26748_, _26743_);
  and (_26750_, _26749_, _26740_);
  nor (_26751_, _26750_, _26705_);
  nor (_26752_, _26751_, _03655_);
  nor (_26753_, _26698_, _05491_);
  not (_26754_, _26753_);
  nor (_26755_, _26745_, _04596_);
  and (_26756_, _26755_, _26754_);
  nor (_26758_, _26756_, _26752_);
  nor (_26759_, _26758_, _03773_);
  nor (_26760_, _26710_, _04594_);
  and (_26761_, _26760_, _26754_);
  nor (_26762_, _26761_, _03653_);
  not (_26763_, _26762_);
  nor (_26764_, _26763_, _26759_);
  nor (_26765_, _13243_, _10485_);
  or (_26766_, _26698_, _04608_);
  nor (_26767_, _26766_, _26765_);
  or (_26769_, _26767_, _03786_);
  nor (_26770_, _26769_, _26764_);
  nor (_26771_, _26770_, _26701_);
  nor (_26772_, _26771_, _03809_);
  nor (_26773_, _26718_, _04260_);
  or (_26774_, _26773_, _03816_);
  nor (_26775_, _26774_, _26772_);
  and (_26776_, _13425_, _05330_);
  or (_26777_, _26698_, _03820_);
  nor (_26778_, _26777_, _26776_);
  nor (_26780_, _26778_, _26775_);
  or (_26781_, _26780_, _43231_);
  or (_26782_, _43227_, \oc8051_golden_model_1.SBUF [6]);
  and (_26783_, _26782_, _41991_);
  and (_43536_, _26783_, _26781_);
  not (_26784_, \oc8051_golden_model_1.SCON [0]);
  nor (_26785_, _05345_, _26784_);
  and (_26786_, _12145_, _05345_);
  nor (_26787_, _26786_, _26785_);
  nor (_26788_, _26787_, _04589_);
  and (_26790_, _05345_, _06366_);
  nor (_26791_, _26790_, _26785_);
  and (_26792_, _26791_, _03650_);
  and (_26793_, _05345_, _04491_);
  nor (_26794_, _26793_, _26785_);
  and (_26795_, _26794_, _07441_);
  and (_26796_, _05345_, \oc8051_golden_model_1.ACC [0]);
  nor (_26797_, _26796_, _26785_);
  nor (_26798_, _26797_, _04500_);
  nor (_26799_, _04499_, _26784_);
  or (_26801_, _26799_, _26798_);
  and (_26802_, _26801_, _04515_);
  nor (_26803_, _05744_, _10566_);
  nor (_26804_, _26803_, _26785_);
  nor (_26805_, _26804_, _04515_);
  or (_26806_, _26805_, _26802_);
  and (_26807_, _26806_, _03516_);
  nor (_26808_, _05976_, _26784_);
  and (_26809_, _12035_, _05976_);
  nor (_26810_, _26809_, _26808_);
  nor (_26812_, _26810_, _03516_);
  nor (_26813_, _26812_, _26807_);
  nor (_26814_, _26813_, _03597_);
  nor (_26815_, _26794_, _04524_);
  or (_26816_, _26815_, _26814_);
  and (_26817_, _26816_, _03611_);
  nor (_26818_, _26797_, _03611_);
  or (_26819_, _26818_, _26817_);
  and (_26820_, _26819_, _03512_);
  and (_26821_, _26785_, _03511_);
  or (_26823_, _26821_, _26820_);
  and (_26824_, _26823_, _03505_);
  nor (_26825_, _26804_, _03505_);
  or (_26826_, _26825_, _26824_);
  and (_26827_, _26826_, _03501_);
  nor (_26828_, _12066_, _10603_);
  nor (_26829_, _26828_, _26808_);
  nor (_26830_, _26829_, _03501_);
  or (_26831_, _26830_, _07441_);
  nor (_26832_, _26831_, _26827_);
  nor (_26834_, _26832_, _26795_);
  nor (_26835_, _26834_, _05969_);
  and (_26836_, _06836_, _05345_);
  nor (_26837_, _26785_, _05970_);
  not (_26838_, _26837_);
  nor (_26839_, _26838_, _26836_);
  or (_26840_, _26839_, _03644_);
  nor (_26841_, _26840_, _26835_);
  nor (_26842_, _12129_, _10566_);
  nor (_26843_, _26842_, _26785_);
  nor (_26845_, _26843_, _03275_);
  or (_26846_, _26845_, _03650_);
  nor (_26847_, _26846_, _26841_);
  nor (_26848_, _26847_, _26792_);
  or (_26849_, _26848_, _03649_);
  and (_26850_, _12019_, _05345_);
  or (_26851_, _26850_, _26785_);
  or (_26852_, _26851_, _04591_);
  and (_26853_, _26852_, _04589_);
  and (_26854_, _26853_, _26849_);
  nor (_26856_, _26854_, _26788_);
  nor (_26857_, _26856_, _03655_);
  or (_26858_, _26791_, _04596_);
  nor (_26859_, _26858_, _26803_);
  nor (_26860_, _26859_, _26857_);
  nor (_26861_, _26860_, _03773_);
  and (_26862_, _12144_, _05345_);
  or (_26863_, _26862_, _26785_);
  and (_26864_, _26863_, _03773_);
  or (_26865_, _26864_, _26861_);
  and (_26867_, _26865_, _04608_);
  nor (_26868_, _12017_, _10566_);
  nor (_26869_, _26868_, _26785_);
  nor (_26870_, _26869_, _04608_);
  or (_26871_, _26870_, _26867_);
  and (_26872_, _26871_, _04606_);
  nor (_26873_, _12015_, _10566_);
  nor (_26874_, _26873_, _26785_);
  nor (_26875_, _26874_, _04606_);
  or (_26876_, _26875_, _26872_);
  and (_26878_, _26876_, _04260_);
  nor (_26879_, _26804_, _04260_);
  or (_26880_, _26879_, _26878_);
  and (_26881_, _26880_, _03206_);
  and (_26882_, _26785_, _03205_);
  nor (_26883_, _26882_, _03816_);
  not (_26884_, _26883_);
  nor (_26885_, _26884_, _26881_);
  and (_26886_, _26804_, _03816_);
  or (_26887_, _26886_, _26885_);
  nand (_26889_, _26887_, _43227_);
  or (_26890_, _43227_, \oc8051_golden_model_1.SCON [0]);
  and (_26891_, _26890_, _41991_);
  and (_43537_, _26891_, _26889_);
  not (_26892_, \oc8051_golden_model_1.SCON [1]);
  nor (_26893_, _05345_, _26892_);
  and (_26894_, _06835_, _05345_);
  or (_26895_, _26894_, _26893_);
  and (_26896_, _26895_, _05969_);
  nor (_26897_, _05345_, \oc8051_golden_model_1.SCON [1]);
  and (_26899_, _05345_, _03320_);
  nor (_26900_, _26899_, _26897_);
  and (_26901_, _26900_, _04499_);
  nor (_26902_, _04499_, _26892_);
  or (_26903_, _26902_, _26901_);
  and (_26904_, _26903_, _04515_);
  and (_26905_, _12234_, _05345_);
  nor (_26906_, _26905_, _26897_);
  and (_26907_, _26906_, _03599_);
  or (_26908_, _26907_, _26904_);
  and (_26910_, _26908_, _03516_);
  nor (_26911_, _05976_, _26892_);
  and (_26912_, _12238_, _05976_);
  nor (_26913_, _26912_, _26911_);
  nor (_26914_, _26913_, _03516_);
  or (_26915_, _26914_, _26910_);
  and (_26916_, _26915_, _04524_);
  and (_26917_, _05345_, _05898_);
  nor (_26918_, _26917_, _26893_);
  nor (_26919_, _26918_, _04524_);
  or (_26920_, _26919_, _26916_);
  and (_26921_, _26920_, _03611_);
  and (_26922_, _26900_, _03603_);
  or (_26923_, _26922_, _26921_);
  and (_26924_, _26923_, _03512_);
  and (_26925_, _12224_, _05976_);
  nor (_26926_, _26925_, _26911_);
  nor (_26927_, _26926_, _03512_);
  or (_26928_, _26927_, _26924_);
  and (_26929_, _26928_, _03505_);
  and (_26932_, _26912_, _12253_);
  or (_26933_, _26932_, _26911_);
  and (_26934_, _26933_, _03504_);
  or (_26935_, _26934_, _26929_);
  and (_26936_, _26935_, _03501_);
  nor (_26937_, _12270_, _10603_);
  nor (_26938_, _26911_, _26937_);
  nor (_26939_, _26938_, _03501_);
  or (_26940_, _26939_, _07441_);
  nor (_26941_, _26940_, _26936_);
  and (_26943_, _26918_, _07441_);
  or (_26944_, _26943_, _05969_);
  nor (_26945_, _26944_, _26941_);
  or (_26946_, _26945_, _26896_);
  and (_26947_, _26946_, _03275_);
  nor (_26948_, _12330_, _10566_);
  nor (_26949_, _26948_, _26893_);
  nor (_26950_, _26949_, _03275_);
  nor (_26951_, _26950_, _26947_);
  nor (_26952_, _26951_, _08861_);
  nor (_26954_, _12220_, _10566_);
  nor (_26955_, _26954_, _04591_);
  and (_26956_, _05345_, _04347_);
  nor (_26957_, _26956_, _04582_);
  nor (_26958_, _26957_, _26955_);
  nor (_26959_, _26958_, _26897_);
  nor (_26960_, _26959_, _26952_);
  nor (_26961_, _26960_, _03778_);
  not (_26962_, _26897_);
  nor (_26963_, _12347_, _10566_);
  nor (_26965_, _26963_, _04589_);
  and (_26966_, _26965_, _26962_);
  nor (_26967_, _26966_, _26961_);
  nor (_26968_, _26967_, _03655_);
  nor (_26969_, _12219_, _10566_);
  nor (_26970_, _26969_, _04596_);
  and (_26971_, _26970_, _26962_);
  nor (_26972_, _26971_, _26968_);
  nor (_26973_, _26972_, _03773_);
  nor (_26974_, _26893_, _05699_);
  nor (_26976_, _26974_, _04594_);
  and (_26977_, _26976_, _26900_);
  nor (_26978_, _26977_, _26973_);
  or (_26979_, _26978_, _18553_);
  and (_26980_, _26899_, _05698_);
  nor (_26981_, _26980_, _04606_);
  and (_26982_, _26981_, _26962_);
  nor (_26983_, _26982_, _03809_);
  and (_26984_, _26956_, _05698_);
  or (_26985_, _26897_, _04608_);
  or (_26987_, _26985_, _26984_);
  and (_26988_, _26987_, _26983_);
  and (_26989_, _26988_, _26979_);
  nor (_26990_, _26906_, _04260_);
  or (_26991_, _26990_, _03205_);
  nor (_26992_, _26991_, _26989_);
  nor (_26993_, _26926_, _03206_);
  or (_26994_, _26993_, _03816_);
  nor (_26995_, _26994_, _26992_);
  nor (_26996_, _26905_, _26893_);
  and (_26998_, _26996_, _03816_);
  nor (_26999_, _26998_, _26995_);
  or (_27000_, _26999_, _43231_);
  or (_27001_, _43227_, \oc8051_golden_model_1.SCON [1]);
  and (_27002_, _27001_, _41991_);
  and (_43540_, _27002_, _27000_);
  not (_27003_, \oc8051_golden_model_1.SCON [2]);
  nor (_27004_, _05345_, _27003_);
  and (_27005_, _05345_, _06414_);
  nor (_27006_, _27005_, _27004_);
  and (_27008_, _27006_, _03650_);
  nor (_27009_, _10566_, _05130_);
  nor (_27010_, _27009_, _27004_);
  and (_27011_, _27010_, _07441_);
  and (_27012_, _05345_, \oc8051_golden_model_1.ACC [2]);
  nor (_27013_, _27012_, _27004_);
  nor (_27014_, _27013_, _04500_);
  nor (_27015_, _04499_, _27003_);
  or (_27016_, _27015_, _27014_);
  and (_27017_, _27016_, _04515_);
  nor (_27019_, _12430_, _10566_);
  nor (_27020_, _27019_, _27004_);
  nor (_27021_, _27020_, _04515_);
  or (_27022_, _27021_, _27017_);
  and (_27023_, _27022_, _03516_);
  nor (_27024_, _05976_, _27003_);
  and (_27025_, _12416_, _05976_);
  nor (_27026_, _27025_, _27024_);
  nor (_27027_, _27026_, _03516_);
  or (_27028_, _27027_, _27023_);
  and (_27029_, _27028_, _04524_);
  nor (_27030_, _27010_, _04524_);
  or (_27031_, _27030_, _27029_);
  and (_27032_, _27031_, _03611_);
  nor (_27033_, _27013_, _03611_);
  or (_27034_, _27033_, _27032_);
  and (_27035_, _27034_, _03512_);
  and (_27036_, _12414_, _05976_);
  nor (_27037_, _27036_, _27024_);
  nor (_27038_, _27037_, _03512_);
  or (_27041_, _27038_, _27035_);
  and (_27042_, _27041_, _03505_);
  and (_27043_, _27025_, _12447_);
  or (_27044_, _27043_, _27024_);
  and (_27045_, _27044_, _03504_);
  or (_27046_, _27045_, _27042_);
  and (_27047_, _27046_, _03501_);
  nor (_27048_, _12465_, _10603_);
  nor (_27049_, _27048_, _27024_);
  nor (_27050_, _27049_, _03501_);
  nor (_27052_, _27050_, _07441_);
  not (_27053_, _27052_);
  nor (_27054_, _27053_, _27047_);
  nor (_27055_, _27054_, _27011_);
  nor (_27056_, _27055_, _05969_);
  and (_27057_, _06839_, _05345_);
  nor (_27058_, _27004_, _05970_);
  not (_27059_, _27058_);
  nor (_27060_, _27059_, _27057_);
  or (_27061_, _27060_, _03644_);
  nor (_27063_, _27061_, _27056_);
  nor (_27064_, _12524_, _10566_);
  nor (_27065_, _27004_, _27064_);
  nor (_27066_, _27065_, _03275_);
  or (_27067_, _27066_, _03650_);
  nor (_27068_, _27067_, _27063_);
  nor (_27069_, _27068_, _27008_);
  or (_27070_, _27069_, _03649_);
  and (_27071_, _12538_, _05345_);
  or (_27072_, _27071_, _27004_);
  or (_27074_, _27072_, _04591_);
  and (_27075_, _27074_, _04589_);
  and (_27076_, _27075_, _27070_);
  and (_27077_, _12544_, _05345_);
  nor (_27078_, _27077_, _27004_);
  nor (_27079_, _27078_, _04589_);
  nor (_27080_, _27079_, _27076_);
  nor (_27081_, _27080_, _03655_);
  nor (_27082_, _27004_, _05793_);
  not (_27083_, _27082_);
  nor (_27085_, _27006_, _04596_);
  and (_27086_, _27085_, _27083_);
  nor (_27087_, _27086_, _27081_);
  nor (_27088_, _27087_, _03773_);
  nor (_27089_, _27013_, _04594_);
  and (_27090_, _27089_, _27083_);
  or (_27091_, _27090_, _27088_);
  and (_27092_, _27091_, _04608_);
  nor (_27093_, _12537_, _10566_);
  nor (_27094_, _27093_, _27004_);
  nor (_27096_, _27094_, _04608_);
  or (_27097_, _27096_, _27092_);
  and (_27098_, _27097_, _04606_);
  nor (_27099_, _12543_, _10566_);
  nor (_27100_, _27099_, _27004_);
  nor (_27101_, _27100_, _04606_);
  or (_27102_, _27101_, _27098_);
  and (_27103_, _27102_, _04260_);
  nor (_27104_, _27020_, _04260_);
  or (_27105_, _27104_, _27103_);
  and (_27107_, _27105_, _03206_);
  nor (_27108_, _27037_, _03206_);
  or (_27109_, _27108_, _27107_);
  and (_27110_, _27109_, _03820_);
  and (_27111_, _12600_, _05345_);
  nor (_27112_, _27111_, _27004_);
  nor (_27113_, _27112_, _03820_);
  or (_27114_, _27113_, _27110_);
  or (_27115_, _27114_, _43231_);
  or (_27116_, _43227_, \oc8051_golden_model_1.SCON [2]);
  and (_27118_, _27116_, _41991_);
  and (_43541_, _27118_, _27115_);
  not (_27119_, \oc8051_golden_model_1.SCON [3]);
  nor (_27120_, _05345_, _27119_);
  and (_27121_, _05345_, _06347_);
  nor (_27122_, _27121_, _27120_);
  and (_27123_, _27122_, _03650_);
  nor (_27124_, _10566_, _04944_);
  nor (_27125_, _27124_, _27120_);
  and (_27126_, _27125_, _07441_);
  and (_27128_, _05345_, \oc8051_golden_model_1.ACC [3]);
  nor (_27129_, _27128_, _27120_);
  nor (_27130_, _27129_, _04500_);
  nor (_27131_, _04499_, _27119_);
  or (_27132_, _27131_, _27130_);
  and (_27133_, _27132_, _04515_);
  nor (_27134_, _12625_, _10566_);
  nor (_27135_, _27134_, _27120_);
  nor (_27136_, _27135_, _04515_);
  or (_27137_, _27136_, _27133_);
  and (_27139_, _27137_, _03516_);
  nor (_27140_, _05976_, _27119_);
  and (_27141_, _12638_, _05976_);
  nor (_27142_, _27141_, _27140_);
  nor (_27143_, _27142_, _03516_);
  or (_27144_, _27143_, _03597_);
  or (_27145_, _27144_, _27139_);
  nand (_27146_, _27125_, _03597_);
  and (_27147_, _27146_, _27145_);
  and (_27148_, _27147_, _03611_);
  nor (_27150_, _27129_, _03611_);
  or (_27151_, _27150_, _27148_);
  and (_27152_, _27151_, _03512_);
  and (_27153_, _12622_, _05976_);
  nor (_27154_, _27153_, _27140_);
  nor (_27155_, _27154_, _03512_);
  or (_27156_, _27155_, _03504_);
  or (_27157_, _27156_, _27152_);
  nor (_27158_, _27140_, _12653_);
  nor (_27159_, _27158_, _27142_);
  or (_27161_, _27159_, _03505_);
  and (_27162_, _27161_, _03501_);
  and (_27163_, _27162_, _27157_);
  nor (_27164_, _12671_, _10603_);
  nor (_27165_, _27164_, _27140_);
  nor (_27166_, _27165_, _03501_);
  nor (_27167_, _27166_, _07441_);
  not (_27168_, _27167_);
  nor (_27169_, _27168_, _27163_);
  nor (_27170_, _27169_, _27126_);
  nor (_27172_, _27170_, _05969_);
  and (_27173_, _06838_, _05345_);
  nor (_27174_, _27120_, _05970_);
  not (_27175_, _27174_);
  nor (_27176_, _27175_, _27173_);
  or (_27177_, _27176_, _03644_);
  nor (_27178_, _27177_, _27172_);
  nor (_27179_, _12731_, _10566_);
  nor (_27180_, _27120_, _27179_);
  nor (_27181_, _27180_, _03275_);
  or (_27183_, _27181_, _03650_);
  nor (_27184_, _27183_, _27178_);
  nor (_27185_, _27184_, _27123_);
  or (_27186_, _27185_, _03649_);
  and (_27187_, _12746_, _05345_);
  or (_27188_, _27187_, _27120_);
  or (_27189_, _27188_, _04591_);
  and (_27190_, _27189_, _04589_);
  and (_27191_, _27190_, _27186_);
  and (_27192_, _12619_, _05345_);
  nor (_27194_, _27192_, _27120_);
  nor (_27195_, _27194_, _04589_);
  nor (_27196_, _27195_, _27191_);
  nor (_27197_, _27196_, _03655_);
  nor (_27198_, _27120_, _05650_);
  not (_27199_, _27198_);
  nor (_27200_, _27122_, _04596_);
  and (_27201_, _27200_, _27199_);
  nor (_27202_, _27201_, _27197_);
  nor (_27203_, _27202_, _03773_);
  nor (_27205_, _27129_, _04594_);
  and (_27206_, _27205_, _27199_);
  nor (_27207_, _27206_, _03653_);
  not (_27208_, _27207_);
  nor (_27209_, _27208_, _27203_);
  nor (_27210_, _12745_, _10566_);
  or (_27211_, _27120_, _04608_);
  nor (_27212_, _27211_, _27210_);
  or (_27213_, _27212_, _03786_);
  nor (_27214_, _27213_, _27209_);
  nor (_27216_, _12618_, _10566_);
  nor (_27217_, _27216_, _27120_);
  nor (_27218_, _27217_, _04606_);
  or (_27219_, _27218_, _27214_);
  and (_27220_, _27219_, _04260_);
  nor (_27221_, _27135_, _04260_);
  or (_27222_, _27221_, _27220_);
  and (_27223_, _27222_, _03206_);
  nor (_27224_, _27154_, _03206_);
  or (_27225_, _27224_, _27223_);
  and (_27227_, _27225_, _03820_);
  and (_27228_, _12806_, _05345_);
  nor (_27229_, _27228_, _27120_);
  nor (_27230_, _27229_, _03820_);
  or (_27231_, _27230_, _27227_);
  or (_27232_, _27231_, _43231_);
  or (_27233_, _43227_, \oc8051_golden_model_1.SCON [3]);
  and (_27234_, _27233_, _41991_);
  and (_43542_, _27234_, _27232_);
  not (_27235_, \oc8051_golden_model_1.SCON [4]);
  nor (_27237_, _05345_, _27235_);
  nor (_27238_, _05840_, _10566_);
  nor (_27239_, _27238_, _27237_);
  and (_27240_, _27239_, _07441_);
  nor (_27241_, _05976_, _27235_);
  and (_27242_, _12853_, _05976_);
  nor (_27243_, _27242_, _27241_);
  nor (_27244_, _27243_, _03512_);
  and (_27245_, _05345_, \oc8051_golden_model_1.ACC [4]);
  nor (_27246_, _27245_, _27237_);
  nor (_27247_, _27246_, _04500_);
  nor (_27248_, _04499_, _27235_);
  or (_27249_, _27248_, _27247_);
  and (_27250_, _27249_, _04515_);
  nor (_27251_, _12820_, _10566_);
  nor (_27252_, _27251_, _27237_);
  nor (_27253_, _27252_, _04515_);
  or (_27254_, _27253_, _27250_);
  and (_27255_, _27254_, _03516_);
  and (_27256_, _12830_, _05976_);
  nor (_27259_, _27256_, _27241_);
  nor (_27260_, _27259_, _03516_);
  or (_27261_, _27260_, _03597_);
  or (_27262_, _27261_, _27255_);
  nand (_27263_, _27239_, _03597_);
  and (_27264_, _27263_, _27262_);
  and (_27265_, _27264_, _03611_);
  nor (_27266_, _27246_, _03611_);
  or (_27267_, _27266_, _27265_);
  and (_27268_, _27267_, _03512_);
  nor (_27270_, _27268_, _27244_);
  nor (_27271_, _27270_, _03504_);
  nor (_27272_, _27241_, _12860_);
  or (_27273_, _27259_, _03505_);
  nor (_27274_, _27273_, _27272_);
  nor (_27275_, _27274_, _27271_);
  nor (_27276_, _27275_, _03500_);
  nor (_27277_, _12828_, _10603_);
  nor (_27278_, _27277_, _27241_);
  nor (_27279_, _27278_, _03501_);
  nor (_27281_, _27279_, _07441_);
  not (_27282_, _27281_);
  nor (_27283_, _27282_, _27276_);
  nor (_27284_, _27283_, _27240_);
  nor (_27285_, _27284_, _05969_);
  and (_27286_, _06843_, _05345_);
  nor (_27287_, _27237_, _05970_);
  not (_27288_, _27287_);
  nor (_27289_, _27288_, _27286_);
  nor (_27290_, _27289_, _03644_);
  not (_27292_, _27290_);
  nor (_27293_, _27292_, _27285_);
  nor (_27294_, _12936_, _10566_);
  nor (_27295_, _27294_, _27237_);
  nor (_27296_, _27295_, _03275_);
  or (_27297_, _27296_, _08861_);
  or (_27298_, _27297_, _27293_);
  and (_27299_, _12951_, _05345_);
  or (_27300_, _27237_, _04591_);
  or (_27301_, _27300_, _27299_);
  and (_27303_, _06375_, _05345_);
  nor (_27304_, _27303_, _27237_);
  and (_27305_, _27304_, _03650_);
  nor (_27306_, _27305_, _03778_);
  and (_27307_, _27306_, _27301_);
  and (_27308_, _27307_, _27298_);
  and (_27309_, _12957_, _05345_);
  nor (_27310_, _27309_, _27237_);
  nor (_27311_, _27310_, _04589_);
  nor (_27312_, _27311_, _27308_);
  nor (_27314_, _27312_, _03655_);
  nor (_27315_, _27237_, _05889_);
  not (_27316_, _27315_);
  nor (_27317_, _27304_, _04596_);
  and (_27318_, _27317_, _27316_);
  nor (_27319_, _27318_, _27314_);
  nor (_27320_, _27319_, _03773_);
  nor (_27321_, _27246_, _04594_);
  and (_27322_, _27321_, _27316_);
  nor (_27323_, _27322_, _03653_);
  not (_27325_, _27323_);
  nor (_27326_, _27325_, _27320_);
  nor (_27327_, _12949_, _10566_);
  or (_27328_, _27237_, _04608_);
  nor (_27329_, _27328_, _27327_);
  or (_27330_, _27329_, _03786_);
  nor (_27331_, _27330_, _27326_);
  nor (_27332_, _12956_, _10566_);
  nor (_27333_, _27332_, _27237_);
  nor (_27334_, _27333_, _04606_);
  or (_27336_, _27334_, _27331_);
  and (_27337_, _27336_, _04260_);
  nor (_27338_, _27252_, _04260_);
  or (_27339_, _27338_, _27337_);
  and (_27340_, _27339_, _03206_);
  nor (_27341_, _27243_, _03206_);
  or (_27342_, _27341_, _27340_);
  and (_27343_, _27342_, _03820_);
  and (_27344_, _13013_, _05345_);
  nor (_27345_, _27344_, _27237_);
  nor (_27347_, _27345_, _03820_);
  or (_27348_, _27347_, _27343_);
  or (_27349_, _27348_, _43231_);
  or (_27350_, _43227_, \oc8051_golden_model_1.SCON [4]);
  and (_27351_, _27350_, _41991_);
  and (_43543_, _27351_, _27349_);
  not (_27352_, \oc8051_golden_model_1.SCON [5]);
  nor (_27353_, _05345_, _27352_);
  and (_27354_, _06842_, _05345_);
  or (_27355_, _27354_, _27353_);
  and (_27357_, _27355_, _05969_);
  and (_27358_, _05345_, \oc8051_golden_model_1.ACC [5]);
  nor (_27359_, _27358_, _27353_);
  nor (_27360_, _27359_, _04500_);
  nor (_27361_, _04499_, _27352_);
  or (_27362_, _27361_, _27360_);
  and (_27363_, _27362_, _04515_);
  nor (_27364_, _13035_, _10566_);
  nor (_27365_, _27364_, _27353_);
  nor (_27366_, _27365_, _04515_);
  or (_27368_, _27366_, _27363_);
  and (_27369_, _27368_, _03516_);
  nor (_27370_, _05976_, _27352_);
  and (_27371_, _13051_, _05976_);
  nor (_27372_, _27371_, _27370_);
  nor (_27373_, _27372_, _03516_);
  or (_27374_, _27373_, _03597_);
  or (_27375_, _27374_, _27369_);
  nor (_27376_, _05552_, _10566_);
  nor (_27377_, _27376_, _27353_);
  nand (_27379_, _27377_, _03597_);
  and (_27380_, _27379_, _27375_);
  and (_27381_, _27380_, _03611_);
  nor (_27382_, _27359_, _03611_);
  or (_27383_, _27382_, _27381_);
  and (_27384_, _27383_, _03512_);
  and (_27385_, _13032_, _05976_);
  nor (_27386_, _27385_, _27370_);
  nor (_27387_, _27386_, _03512_);
  or (_27388_, _27387_, _27384_);
  and (_27390_, _27388_, _03505_);
  nor (_27391_, _27370_, _13066_);
  nor (_27392_, _27391_, _27372_);
  and (_27393_, _27392_, _03504_);
  or (_27394_, _27393_, _27390_);
  and (_27395_, _27394_, _03501_);
  nor (_27396_, _13030_, _10603_);
  nor (_27397_, _27396_, _27370_);
  nor (_27398_, _27397_, _03501_);
  nor (_27399_, _27398_, _07441_);
  not (_27401_, _27399_);
  nor (_27402_, _27401_, _27395_);
  and (_27403_, _27377_, _07441_);
  or (_27404_, _27403_, _05969_);
  nor (_27405_, _27404_, _27402_);
  or (_27406_, _27405_, _27357_);
  and (_27407_, _27406_, _03275_);
  nor (_27408_, _13139_, _10566_);
  nor (_27409_, _27408_, _27353_);
  nor (_27410_, _27409_, _03275_);
  or (_27412_, _27410_, _08861_);
  or (_27413_, _27412_, _27407_);
  and (_27414_, _13154_, _05345_);
  or (_27415_, _27353_, _04591_);
  or (_27416_, _27415_, _27414_);
  and (_27417_, _06358_, _05345_);
  nor (_27418_, _27417_, _27353_);
  and (_27419_, _27418_, _03650_);
  nor (_27420_, _27419_, _03778_);
  and (_27421_, _27420_, _27416_);
  and (_27423_, _27421_, _27413_);
  and (_27424_, _13160_, _05345_);
  nor (_27425_, _27424_, _27353_);
  nor (_27426_, _27425_, _04589_);
  nor (_27427_, _27426_, _27423_);
  nor (_27428_, _27427_, _03655_);
  nor (_27429_, _27353_, _05601_);
  not (_27430_, _27429_);
  nor (_27431_, _27418_, _04596_);
  and (_27432_, _27431_, _27430_);
  nor (_27434_, _27432_, _27428_);
  nor (_27435_, _27434_, _03773_);
  nor (_27436_, _27359_, _04594_);
  and (_27437_, _27436_, _27430_);
  nor (_27438_, _27437_, _03653_);
  not (_27439_, _27438_);
  nor (_27440_, _27439_, _27435_);
  nor (_27441_, _13152_, _10566_);
  or (_27442_, _27353_, _04608_);
  nor (_27443_, _27442_, _27441_);
  or (_27445_, _27443_, _03786_);
  nor (_27446_, _27445_, _27440_);
  nor (_27447_, _13159_, _10566_);
  nor (_27448_, _27447_, _27353_);
  nor (_27449_, _27448_, _04606_);
  or (_27450_, _27449_, _27446_);
  and (_27451_, _27450_, _04260_);
  nor (_27452_, _27365_, _04260_);
  or (_27453_, _27452_, _27451_);
  and (_27454_, _27453_, _03206_);
  nor (_27456_, _27386_, _03206_);
  or (_27457_, _27456_, _27454_);
  and (_27458_, _27457_, _03820_);
  and (_27459_, _13217_, _05345_);
  nor (_27460_, _27459_, _27353_);
  nor (_27461_, _27460_, _03820_);
  or (_27462_, _27461_, _27458_);
  or (_27463_, _27462_, _43231_);
  or (_27464_, _43227_, \oc8051_golden_model_1.SCON [5]);
  and (_27465_, _27464_, _41991_);
  and (_43544_, _27465_, _27463_);
  not (_27467_, \oc8051_golden_model_1.SCON [6]);
  nor (_27468_, _05345_, _27467_);
  and (_27469_, _06531_, _05345_);
  or (_27470_, _27469_, _27468_);
  and (_27471_, _27470_, _05969_);
  and (_27472_, _05345_, \oc8051_golden_model_1.ACC [6]);
  nor (_27473_, _27472_, _27468_);
  nor (_27474_, _27473_, _04500_);
  nor (_27475_, _04499_, _27467_);
  or (_27477_, _27475_, _27474_);
  and (_27478_, _27477_, _04515_);
  nor (_27479_, _13235_, _10566_);
  nor (_27480_, _27479_, _27468_);
  nor (_27481_, _27480_, _04515_);
  or (_27482_, _27481_, _27478_);
  and (_27483_, _27482_, _03516_);
  nor (_27484_, _05976_, _27467_);
  and (_27485_, _13266_, _05976_);
  nor (_27486_, _27485_, _27484_);
  nor (_27488_, _27486_, _03516_);
  or (_27489_, _27488_, _03597_);
  or (_27490_, _27489_, _27483_);
  nor (_27491_, _05442_, _10566_);
  nor (_27492_, _27491_, _27468_);
  nand (_27493_, _27492_, _03597_);
  and (_27494_, _27493_, _27490_);
  and (_27495_, _27494_, _03611_);
  nor (_27496_, _27473_, _03611_);
  or (_27497_, _27496_, _27495_);
  and (_27499_, _27497_, _03512_);
  and (_27500_, _13251_, _05976_);
  nor (_27501_, _27500_, _27484_);
  nor (_27502_, _27501_, _03512_);
  or (_27503_, _27502_, _03504_);
  or (_27504_, _27503_, _27499_);
  nor (_27505_, _27484_, _13281_);
  nor (_27506_, _27505_, _27486_);
  or (_27507_, _27506_, _03505_);
  and (_27508_, _27507_, _03501_);
  and (_27509_, _27508_, _27504_);
  nor (_27510_, _13249_, _10603_);
  nor (_27511_, _27510_, _27484_);
  nor (_27512_, _27511_, _03501_);
  nor (_27513_, _27512_, _07441_);
  not (_27514_, _27513_);
  nor (_27515_, _27514_, _27509_);
  and (_27516_, _27492_, _07441_);
  or (_27517_, _27516_, _05969_);
  nor (_27518_, _27517_, _27515_);
  or (_27521_, _27518_, _27471_);
  and (_27522_, _27521_, _03275_);
  nor (_27523_, _13356_, _10566_);
  nor (_27524_, _27523_, _27468_);
  nor (_27525_, _27524_, _03275_);
  or (_27526_, _27525_, _08861_);
  or (_27527_, _27526_, _27522_);
  and (_27528_, _13245_, _05345_);
  or (_27529_, _27468_, _04591_);
  or (_27530_, _27529_, _27528_);
  and (_27532_, _13363_, _05345_);
  nor (_27533_, _27532_, _27468_);
  and (_27534_, _27533_, _03650_);
  nor (_27535_, _27534_, _03778_);
  and (_27536_, _27535_, _27530_);
  and (_27537_, _27536_, _27527_);
  and (_27538_, _13374_, _05345_);
  nor (_27539_, _27538_, _27468_);
  nor (_27540_, _27539_, _04589_);
  nor (_27541_, _27540_, _27537_);
  nor (_27543_, _27541_, _03655_);
  nor (_27544_, _27468_, _05491_);
  not (_27545_, _27544_);
  nor (_27546_, _27533_, _04596_);
  and (_27547_, _27546_, _27545_);
  nor (_27548_, _27547_, _27543_);
  nor (_27549_, _27548_, _03773_);
  nor (_27550_, _27473_, _04594_);
  and (_27551_, _27550_, _27545_);
  nor (_27552_, _27551_, _03653_);
  not (_27554_, _27552_);
  nor (_27555_, _27554_, _27549_);
  nor (_27556_, _13243_, _10566_);
  or (_27557_, _27468_, _04608_);
  nor (_27558_, _27557_, _27556_);
  or (_27559_, _27558_, _03786_);
  nor (_27560_, _27559_, _27555_);
  nor (_27561_, _13373_, _10566_);
  nor (_27562_, _27561_, _27468_);
  nor (_27563_, _27562_, _04606_);
  or (_27565_, _27563_, _27560_);
  and (_27566_, _27565_, _04260_);
  nor (_27567_, _27480_, _04260_);
  or (_27568_, _27567_, _27566_);
  and (_27569_, _27568_, _03206_);
  nor (_27570_, _27501_, _03206_);
  or (_27571_, _27570_, _27569_);
  and (_27572_, _27571_, _03820_);
  and (_27573_, _13425_, _05345_);
  nor (_27574_, _27573_, _27468_);
  nor (_27576_, _27574_, _03820_);
  or (_27577_, _27576_, _27572_);
  or (_27578_, _27577_, _43231_);
  or (_27579_, _43227_, \oc8051_golden_model_1.SCON [6]);
  and (_27580_, _27579_, _41991_);
  and (_43545_, _27580_, _27578_);
  nor (_27581_, _05315_, _04079_);
  nor (_27582_, _05744_, _10686_);
  nor (_27583_, _27582_, _27581_);
  and (_27584_, _27583_, _17220_);
  and (_27586_, _27583_, _03599_);
  and (_27587_, _05315_, \oc8051_golden_model_1.ACC [0]);
  nor (_27588_, _27587_, _27581_);
  nor (_27589_, _27588_, _04500_);
  nor (_27590_, _04499_, _04079_);
  or (_27591_, _27590_, _03599_);
  nor (_27592_, _27591_, _27589_);
  nor (_27593_, _27592_, _27586_);
  and (_27594_, _27593_, _04524_);
  or (_27595_, _27594_, _04080_);
  and (_27597_, _27595_, _03611_);
  nor (_27598_, _27588_, _03611_);
  or (_27599_, _27598_, _27597_);
  and (_27600_, _27599_, _04650_);
  nor (_27601_, _07441_, _04540_);
  not (_27602_, _27601_);
  nor (_27603_, _27602_, _27600_);
  not (_27604_, _27581_);
  and (_27605_, _05315_, _04491_);
  nor (_27606_, _27605_, _06889_);
  and (_27608_, _27606_, _27604_);
  nor (_27609_, _27608_, _27603_);
  nor (_27610_, _27609_, _05969_);
  and (_27611_, _06836_, _05315_);
  nor (_27612_, _27581_, _05970_);
  not (_27613_, _27612_);
  nor (_27614_, _27613_, _27611_);
  nor (_27615_, _27614_, _27610_);
  nor (_27616_, _27615_, _03644_);
  nor (_27617_, _12129_, _10686_);
  or (_27619_, _27581_, _03275_);
  nor (_27620_, _27619_, _27617_);
  or (_27621_, _27620_, _03650_);
  nor (_27622_, _27621_, _27616_);
  and (_27623_, _05315_, _06366_);
  nor (_27624_, _27623_, _27581_);
  nand (_27625_, _27624_, _04591_);
  and (_27626_, _27625_, _08861_);
  nor (_27627_, _27626_, _27622_);
  and (_27628_, _12019_, _05315_);
  nor (_27630_, _27628_, _27581_);
  and (_27631_, _27630_, _03649_);
  nor (_27632_, _27631_, _27627_);
  nor (_27633_, _27632_, _03778_);
  and (_27634_, _12145_, _05315_);
  or (_27635_, _27581_, _04589_);
  nor (_27636_, _27635_, _27634_);
  or (_27637_, _27636_, _03655_);
  nor (_27638_, _27637_, _27633_);
  or (_27639_, _27624_, _04596_);
  nor (_27641_, _27639_, _27582_);
  nor (_27642_, _27641_, _27638_);
  nor (_27643_, _27642_, _03773_);
  and (_27644_, _12144_, _05315_);
  or (_27645_, _27644_, _27581_);
  and (_27646_, _27645_, _03773_);
  or (_27647_, _27646_, _27643_);
  and (_27648_, _27647_, _04608_);
  nor (_27649_, _12017_, _10686_);
  nor (_27650_, _27649_, _27581_);
  nor (_27652_, _27650_, _04608_);
  or (_27653_, _27652_, _27648_);
  and (_27654_, _27653_, _04606_);
  nor (_27655_, _12015_, _10686_);
  nor (_27656_, _27655_, _27581_);
  nor (_27657_, _27656_, _04606_);
  nor (_27658_, _27657_, _17220_);
  not (_27659_, _27658_);
  nor (_27660_, _27659_, _27654_);
  nor (_27661_, _27660_, _27584_);
  and (_27663_, _27661_, _43227_);
  nor (_27664_, \oc8051_golden_model_1.SP [0], rst);
  nor (_27665_, _27664_, _00000_);
  or (_43548_, _27665_, _27663_);
  nor (_27666_, _05315_, _04365_);
  and (_27667_, _12234_, _05315_);
  nor (_27668_, _27667_, _27666_);
  nor (_27669_, _27668_, _03820_);
  not (_27670_, _10796_);
  and (_27671_, _03227_, _04365_);
  not (_27673_, _03227_);
  nor (_27674_, _05315_, \oc8051_golden_model_1.SP [1]);
  and (_27675_, _05315_, _03320_);
  nor (_27676_, _27675_, _27674_);
  and (_27677_, _27676_, _04499_);
  nor (_27678_, _04499_, _04365_);
  or (_27679_, _27678_, _27677_);
  and (_27680_, _27679_, _04868_);
  and (_27681_, _03947_, _04365_);
  or (_27682_, _27681_, _27680_);
  and (_27684_, _27682_, _04515_);
  nor (_27685_, _27674_, _27667_);
  and (_27686_, _27685_, _03599_);
  or (_27687_, _27686_, _27684_);
  and (_27688_, _27687_, _03257_);
  nor (_27689_, _03257_, \oc8051_golden_model_1.SP [1]);
  or (_27690_, _27689_, _03597_);
  or (_27691_, _27690_, _27688_);
  nand (_27692_, _04647_, _03597_);
  and (_27693_, _27692_, _27691_);
  and (_27695_, _27693_, _03611_);
  and (_27696_, _27676_, _03603_);
  or (_27697_, _27696_, _27695_);
  and (_27698_, _27697_, _04650_);
  or (_27699_, _27698_, _10729_);
  nor (_27700_, _27699_, _04649_);
  nor (_27701_, _04856_, _04365_);
  or (_27702_, _27701_, _07441_);
  nor (_27703_, _27702_, _27700_);
  or (_27704_, _10686_, _05898_);
  nor (_27706_, _27674_, _06889_);
  and (_27707_, _27706_, _27704_);
  nor (_27708_, _27707_, _05969_);
  not (_27709_, _27708_);
  nor (_27710_, _27709_, _27703_);
  and (_27711_, _06835_, _05315_);
  nor (_27712_, _27666_, _05970_);
  not (_27713_, _27712_);
  nor (_27714_, _27713_, _27711_);
  nor (_27715_, _27714_, _03644_);
  not (_27717_, _27715_);
  nor (_27718_, _27717_, _27710_);
  nor (_27719_, _12330_, _10686_);
  or (_27720_, _27719_, _27666_);
  and (_27721_, _27720_, _03644_);
  nor (_27722_, _27721_, _27718_);
  nor (_27723_, _27722_, _03650_);
  and (_27724_, _05315_, _06249_);
  or (_27725_, _27724_, _27666_);
  and (_27726_, _27725_, _03650_);
  or (_27728_, _27726_, _27723_);
  and (_27729_, _27728_, _27673_);
  or (_27730_, _27729_, _27671_);
  and (_27731_, _27730_, _04591_);
  nor (_27732_, _12220_, _10686_);
  or (_27733_, _27732_, _04591_);
  nor (_27734_, _27733_, _27674_);
  nor (_27735_, _27734_, _27731_);
  nor (_27736_, _27735_, _03778_);
  nor (_27737_, _12347_, _10686_);
  or (_27739_, _27737_, _04589_);
  nor (_27740_, _27739_, _27674_);
  nor (_27741_, _27740_, _27736_);
  nor (_27742_, _27741_, _03655_);
  nor (_27743_, _12219_, _10686_);
  or (_27744_, _27743_, _04596_);
  nor (_27745_, _27744_, _27674_);
  nor (_27746_, _27745_, _27742_);
  nor (_27747_, _27746_, _10777_);
  and (_27748_, _03238_, _04365_);
  nor (_27750_, _27666_, _05699_);
  nor (_27751_, _27750_, _04594_);
  and (_27752_, _27751_, _27676_);
  nor (_27753_, _27752_, _27748_);
  not (_27754_, _27753_);
  nor (_27755_, _27754_, _27747_);
  nor (_27756_, _27755_, _18553_);
  nor (_27757_, _12346_, _10686_);
  or (_27758_, _27757_, _27666_);
  and (_27759_, _27758_, _03786_);
  nor (_27761_, _12218_, _10686_);
  or (_27762_, _27761_, _27666_);
  and (_27763_, _27762_, _03653_);
  nor (_27764_, _27763_, _27759_);
  not (_27765_, _27764_);
  nor (_27766_, _27765_, _27756_);
  nor (_27767_, _27766_, _27670_);
  nor (_27768_, _10796_, \oc8051_golden_model_1.SP [1]);
  nor (_27769_, _27768_, _03521_);
  not (_27770_, _27769_);
  nor (_27772_, _27770_, _27767_);
  nor (_27773_, _04372_, _03809_);
  not (_27774_, _27773_);
  nor (_27775_, _27774_, _27772_);
  and (_27776_, _27685_, _03809_);
  nor (_27777_, _27776_, _05047_);
  not (_27778_, _27777_);
  nor (_27779_, _27778_, _27775_);
  nor (_27780_, _04625_, _04365_);
  nor (_27781_, _27780_, _03816_);
  not (_27783_, _27781_);
  nor (_27784_, _27783_, _27779_);
  nor (_27785_, _27784_, _27669_);
  nor (_27786_, _27785_, _43231_);
  nor (_27787_, \oc8051_golden_model_1.SP [1], rst);
  nor (_27788_, _27787_, _00000_);
  or (_43549_, _27788_, _27786_);
  and (_27789_, _05213_, _03248_);
  and (_27790_, _05213_, _03238_);
  nor (_27791_, _27790_, _03653_);
  nor (_27792_, _05315_, _06069_);
  and (_27793_, _12544_, _05315_);
  nor (_27794_, _27793_, _27792_);
  nor (_27795_, _27794_, _04589_);
  and (_27796_, _13449_, _03227_);
  not (_27797_, _27792_);
  nor (_27798_, _10686_, _05130_);
  nor (_27799_, _27798_, _06889_);
  and (_27800_, _27799_, _27797_);
  nor (_27801_, _13449_, _03253_);
  nor (_27804_, _04499_, _06069_);
  and (_27805_, _05315_, \oc8051_golden_model_1.ACC [2]);
  nor (_27806_, _27805_, _27792_);
  nor (_27807_, _27806_, _04500_);
  or (_27808_, _27807_, _27804_);
  and (_27809_, _27808_, _04868_);
  and (_27810_, _05213_, _03947_);
  nor (_27811_, _27810_, _27809_);
  nor (_27812_, _27811_, _03599_);
  nor (_27813_, _12430_, _10686_);
  nor (_27815_, _27813_, _27792_);
  nor (_27816_, _27815_, _04515_);
  or (_27817_, _27816_, _27812_);
  and (_27818_, _27817_, _03257_);
  nor (_27819_, _13449_, _03257_);
  or (_27820_, _27819_, _03597_);
  or (_27821_, _27820_, _27818_);
  nand (_27822_, _06101_, _03597_);
  and (_27823_, _27822_, _27821_);
  and (_27824_, _27823_, _03611_);
  nor (_27826_, _27806_, _03611_);
  or (_27827_, _27826_, _27824_);
  and (_27828_, _27827_, _04650_);
  or (_27829_, _27828_, _05156_);
  and (_27830_, _27829_, _03253_);
  or (_27831_, _27830_, _27801_);
  and (_27832_, _27831_, _03278_);
  nor (_27833_, _13449_, _03278_);
  nor (_27834_, _27833_, _07441_);
  not (_27835_, _27834_);
  nor (_27837_, _27835_, _27832_);
  nor (_27838_, _27837_, _27800_);
  nor (_27839_, _27838_, _05969_);
  and (_27840_, _06839_, _05315_);
  nor (_27841_, _27792_, _05970_);
  not (_27842_, _27841_);
  nor (_27843_, _27842_, _27840_);
  or (_27844_, _27843_, _03644_);
  nor (_27845_, _27844_, _27839_);
  nor (_27846_, _12524_, _10686_);
  nor (_27848_, _27846_, _27792_);
  nor (_27849_, _27848_, _03275_);
  or (_27850_, _27849_, _03650_);
  or (_27851_, _27850_, _27845_);
  and (_27852_, _05315_, _06414_);
  nor (_27853_, _27852_, _27792_);
  nand (_27854_, _27853_, _03650_);
  and (_27855_, _27854_, _27851_);
  nor (_27856_, _27855_, _03227_);
  nor (_27857_, _27856_, _27796_);
  nor (_27859_, _27857_, _03649_);
  and (_27860_, _12538_, _05315_);
  or (_27861_, _27792_, _04591_);
  nor (_27862_, _27861_, _27860_);
  or (_27863_, _27862_, _03778_);
  nor (_27864_, _27863_, _27859_);
  nor (_27865_, _27864_, _27795_);
  nor (_27866_, _27865_, _03655_);
  and (_27867_, _27797_, _05792_);
  not (_27868_, _27867_);
  nor (_27870_, _27853_, _04596_);
  and (_27871_, _27870_, _27868_);
  nor (_27872_, _27871_, _27866_);
  nor (_27873_, _27872_, _10777_);
  nor (_27874_, _27806_, _04594_);
  and (_27875_, _27874_, _27868_);
  nor (_27876_, _27875_, _27873_);
  and (_27877_, _27876_, _27791_);
  nor (_27878_, _12537_, _10686_);
  nor (_27879_, _27878_, _27792_);
  and (_27881_, _27879_, _03653_);
  nor (_27882_, _27881_, _27877_);
  nor (_27883_, _27882_, _03786_);
  nor (_27884_, _12543_, _10686_);
  or (_27885_, _27792_, _04606_);
  nor (_27886_, _27885_, _27884_);
  or (_27887_, _27886_, _03792_);
  nor (_27888_, _27887_, _27883_);
  and (_27889_, _13449_, _03792_);
  or (_27890_, _27889_, _27888_);
  and (_27892_, _27890_, _06475_);
  or (_27893_, _27892_, _27789_);
  and (_27894_, _27893_, _03522_);
  and (_27895_, _13449_, _03521_);
  or (_27896_, _27895_, _03809_);
  nor (_27897_, _27896_, _27894_);
  and (_27898_, _27815_, _03809_);
  or (_27899_, _27898_, _05047_);
  nor (_27900_, _27899_, _27897_);
  nor (_27901_, _13449_, _04625_);
  nor (_27903_, _27901_, _03816_);
  not (_27904_, _27903_);
  nor (_27905_, _27904_, _27900_);
  and (_27906_, _12600_, _05315_);
  nor (_27907_, _27906_, _27792_);
  and (_27908_, _27907_, _03816_);
  nor (_27909_, _27908_, _27905_);
  and (_27910_, _27909_, _43227_);
  nor (_27911_, \oc8051_golden_model_1.SP [2], rst);
  nor (_27912_, _27911_, _00000_);
  or (_43550_, _27912_, _27910_);
  nor (_27914_, _05216_, _04625_);
  and (_27915_, _05216_, _03248_);
  nor (_27916_, _05315_, _03596_);
  and (_27917_, _12619_, _05315_);
  nor (_27918_, _27917_, _27916_);
  nor (_27919_, _27918_, _04589_);
  nor (_27920_, _05216_, _04856_);
  nor (_27921_, _04499_, _03596_);
  and (_27922_, _05315_, \oc8051_golden_model_1.ACC [3]);
  nor (_27924_, _27922_, _27916_);
  nor (_27925_, _27924_, _04500_);
  or (_27926_, _27925_, _27921_);
  and (_27927_, _27926_, _04868_);
  and (_27928_, _05216_, _03947_);
  nor (_27929_, _27928_, _27927_);
  nor (_27930_, _27929_, _03599_);
  nor (_27931_, _12625_, _10686_);
  nor (_27932_, _27931_, _27916_);
  nor (_27933_, _27932_, _04515_);
  or (_27935_, _27933_, _27930_);
  and (_27936_, _27935_, _03257_);
  nor (_27937_, _13453_, _03257_);
  or (_27938_, _27937_, _03597_);
  or (_27939_, _27938_, _27936_);
  nand (_27940_, _06076_, _03597_);
  and (_27941_, _27940_, _27939_);
  and (_27942_, _27941_, _03611_);
  nor (_27943_, _27924_, _03611_);
  or (_27944_, _27943_, _27942_);
  and (_27946_, _27944_, _04650_);
  or (_27947_, _27946_, _10729_);
  nor (_27948_, _27947_, _04992_);
  nor (_27949_, _27948_, _27920_);
  nor (_27950_, _27949_, _06888_);
  nor (_27951_, _10686_, _04944_);
  nor (_27952_, _27951_, _27916_);
  nor (_27953_, _27952_, _04131_);
  nor (_27954_, _27953_, _06889_);
  nor (_27955_, _27954_, _27950_);
  not (_27957_, _04131_);
  nor (_27958_, _27952_, _27957_);
  nor (_27959_, _27958_, _05969_);
  not (_27960_, _27959_);
  nor (_27961_, _27960_, _27955_);
  and (_27962_, _06838_, _05315_);
  nor (_27963_, _27916_, _05970_);
  not (_27964_, _27963_);
  nor (_27965_, _27964_, _27962_);
  nor (_27966_, _27965_, _03644_);
  not (_27968_, _27966_);
  nor (_27969_, _27968_, _27961_);
  nor (_27970_, _12731_, _10686_);
  nor (_27971_, _27970_, _27916_);
  nor (_27972_, _27971_, _03275_);
  or (_27973_, _27972_, _27969_);
  and (_27974_, _27973_, _04582_);
  and (_27975_, _05315_, _06347_);
  nor (_27976_, _27975_, _27916_);
  nor (_27977_, _27976_, _04582_);
  or (_27979_, _27977_, _27974_);
  and (_27980_, _27979_, _27673_);
  and (_27981_, _05216_, _03227_);
  or (_27982_, _27981_, _03649_);
  nor (_27983_, _27982_, _27980_);
  and (_27984_, _12746_, _05315_);
  or (_27985_, _27916_, _04591_);
  nor (_27986_, _27985_, _27984_);
  or (_27987_, _27986_, _03778_);
  nor (_27988_, _27987_, _27983_);
  nor (_27990_, _27988_, _27919_);
  nor (_27991_, _27990_, _03655_);
  nor (_27992_, _27916_, _05650_);
  not (_27993_, _27992_);
  nor (_27994_, _27976_, _04596_);
  and (_27995_, _27994_, _27993_);
  nor (_27996_, _27995_, _27991_);
  nor (_27997_, _27996_, _10777_);
  nor (_27998_, _27924_, _04594_);
  and (_27999_, _27998_, _27993_);
  and (_28001_, _05216_, _03238_);
  nor (_28002_, _28001_, _27999_);
  and (_28003_, _28002_, _04608_);
  not (_28004_, _28003_);
  nor (_28005_, _28004_, _27997_);
  nor (_28006_, _12745_, _10686_);
  nor (_28007_, _28006_, _27916_);
  and (_28008_, _28007_, _03653_);
  nor (_28009_, _28008_, _28005_);
  nor (_28010_, _28009_, _03786_);
  nor (_28012_, _12618_, _10686_);
  or (_28013_, _27916_, _04606_);
  nor (_28014_, _28013_, _28012_);
  or (_28015_, _28014_, _03792_);
  nor (_28016_, _28015_, _28010_);
  nor (_28017_, _06073_, _03596_);
  nor (_28018_, _28017_, _06074_);
  nor (_28019_, _28018_, _10680_);
  or (_28020_, _28019_, _28016_);
  and (_28021_, _28020_, _06475_);
  or (_28023_, _28021_, _27915_);
  and (_28024_, _28023_, _03522_);
  nor (_28025_, _28018_, _03522_);
  or (_28026_, _28025_, _28024_);
  and (_28027_, _28026_, _04260_);
  nor (_28028_, _27932_, _04260_);
  nor (_28029_, _28028_, _05047_);
  not (_28030_, _28029_);
  nor (_28031_, _28030_, _28027_);
  nor (_28032_, _28031_, _27914_);
  and (_28034_, _28032_, _03820_);
  and (_28035_, _12806_, _05315_);
  nor (_28036_, _28035_, _27916_);
  nor (_28037_, _28036_, _03820_);
  or (_28038_, _28037_, _28034_);
  or (_28039_, _28038_, _43231_);
  or (_28040_, _43227_, \oc8051_golden_model_1.SP [3]);
  and (_28041_, _28040_, _41991_);
  and (_43551_, _28041_, _28039_);
  nor (_28042_, _04952_, \oc8051_golden_model_1.SP [4]);
  nor (_28044_, _28042_, _10672_);
  nor (_28045_, _28044_, _04625_);
  nor (_28046_, _05315_, _10714_);
  and (_28047_, _12957_, _05315_);
  nor (_28048_, _28047_, _28046_);
  nor (_28049_, _28048_, _04589_);
  nor (_28050_, _05840_, _10686_);
  nor (_28051_, _28050_, _28046_);
  nor (_28052_, _28051_, _06889_);
  or (_28053_, _28052_, _05969_);
  and (_28055_, _04953_, \oc8051_golden_model_1.SP [4]);
  nor (_28056_, _04953_, \oc8051_golden_model_1.SP [4]);
  nor (_28057_, _28056_, _28055_);
  and (_28058_, _28057_, _03510_);
  nor (_28059_, _04499_, _10714_);
  and (_28060_, _05315_, \oc8051_golden_model_1.ACC [4]);
  nor (_28061_, _28060_, _28046_);
  nor (_28062_, _28061_, _04500_);
  or (_28063_, _28062_, _28059_);
  and (_28064_, _28063_, _04868_);
  and (_28066_, _28044_, _03947_);
  nor (_28067_, _28066_, _28064_);
  nor (_28068_, _28067_, _03599_);
  nor (_28069_, _12820_, _10686_);
  nor (_28070_, _28069_, _28046_);
  nor (_28071_, _28070_, _04515_);
  or (_28072_, _28071_, _28068_);
  and (_28073_, _28072_, _03257_);
  not (_28074_, _28044_);
  nor (_28075_, _28074_, _03257_);
  or (_28077_, _28075_, _28073_);
  and (_28078_, _28077_, _04524_);
  and (_28079_, _10715_, _04079_);
  nor (_28080_, _06075_, _10714_);
  nor (_28081_, _28080_, _28079_);
  nor (_28082_, _28081_, _04524_);
  or (_28083_, _28082_, _28078_);
  and (_28084_, _28083_, _03611_);
  nor (_28085_, _28061_, _03611_);
  or (_28086_, _28085_, _28084_);
  and (_28088_, _28086_, _04650_);
  or (_28089_, _28088_, _10729_);
  nor (_28090_, _28089_, _28058_);
  nor (_28091_, _28044_, _04856_);
  or (_28092_, _28091_, _07441_);
  nor (_28093_, _28092_, _28090_);
  nor (_28094_, _28093_, _28053_);
  and (_28095_, _06843_, _05315_);
  nor (_28096_, _28046_, _05970_);
  not (_28097_, _28096_);
  nor (_28099_, _28097_, _28095_);
  or (_28100_, _28099_, _03644_);
  nor (_28101_, _28100_, _28094_);
  nor (_28102_, _12936_, _10686_);
  nor (_28103_, _28102_, _28046_);
  nor (_28104_, _28103_, _03275_);
  or (_28105_, _28104_, _03650_);
  or (_28106_, _28105_, _28101_);
  and (_28107_, _06375_, _05315_);
  nor (_28108_, _28107_, _28046_);
  nand (_28110_, _28108_, _03650_);
  and (_28111_, _28110_, _28106_);
  nor (_28112_, _28111_, _03227_);
  and (_28113_, _28074_, _03227_);
  nor (_28114_, _28113_, _28112_);
  nor (_28115_, _28114_, _03649_);
  and (_28116_, _12951_, _05315_);
  or (_28117_, _28046_, _04591_);
  nor (_28118_, _28117_, _28116_);
  or (_28119_, _28118_, _03778_);
  nor (_28121_, _28119_, _28115_);
  nor (_28122_, _28121_, _28049_);
  nor (_28123_, _28122_, _03655_);
  nor (_28124_, _28046_, _05889_);
  not (_28125_, _28124_);
  nor (_28126_, _28108_, _04596_);
  and (_28127_, _28126_, _28125_);
  nor (_28128_, _28127_, _28123_);
  nor (_28129_, _28128_, _10777_);
  nor (_28130_, _28061_, _04594_);
  and (_28132_, _28130_, _28125_);
  and (_28133_, _28044_, _03238_);
  nor (_28134_, _28133_, _28132_);
  and (_28135_, _28134_, _04608_);
  not (_28136_, _28135_);
  nor (_28137_, _28136_, _28129_);
  nor (_28138_, _12949_, _10686_);
  nor (_28139_, _28138_, _28046_);
  and (_28140_, _28139_, _03653_);
  nor (_28141_, _28140_, _28137_);
  nor (_28143_, _28141_, _03786_);
  nor (_28144_, _12956_, _10686_);
  or (_28145_, _28046_, _04606_);
  nor (_28146_, _28145_, _28144_);
  or (_28147_, _28146_, _03792_);
  nor (_28148_, _28147_, _28143_);
  nor (_28149_, _06074_, _10714_);
  nor (_28150_, _28149_, _10715_);
  nor (_28151_, _28150_, _10680_);
  or (_28152_, _28151_, _28148_);
  and (_28154_, _28152_, _06475_);
  and (_28155_, _28044_, _03248_);
  or (_28156_, _28155_, _28154_);
  and (_28157_, _28156_, _03522_);
  nor (_28158_, _28150_, _03522_);
  or (_28159_, _28158_, _28157_);
  and (_28160_, _28159_, _04260_);
  nor (_28161_, _28070_, _04260_);
  nor (_28162_, _28161_, _05047_);
  not (_28163_, _28162_);
  nor (_28165_, _28163_, _28160_);
  nor (_28166_, _28165_, _28045_);
  and (_28167_, _28166_, _03820_);
  and (_28168_, _13013_, _05315_);
  nor (_28169_, _28168_, _28046_);
  nor (_28170_, _28169_, _03820_);
  or (_28171_, _28170_, _28167_);
  or (_28172_, _28171_, _43231_);
  or (_28173_, _43227_, \oc8051_golden_model_1.SP [4]);
  and (_28174_, _28173_, _41991_);
  and (_43552_, _28174_, _28172_);
  nor (_28176_, _10672_, \oc8051_golden_model_1.SP [5]);
  nor (_28177_, _28176_, _10673_);
  nor (_28178_, _28177_, _04625_);
  and (_28179_, _28177_, _03238_);
  nor (_28180_, _28179_, _03653_);
  nor (_28181_, _05315_, _10713_);
  and (_28182_, _13160_, _05315_);
  nor (_28183_, _28182_, _28181_);
  nor (_28184_, _28183_, _04589_);
  nor (_28186_, _05552_, _10686_);
  nor (_28187_, _28186_, _28181_);
  nor (_28188_, _28187_, _06889_);
  or (_28189_, _28188_, _05969_);
  nor (_28190_, _04499_, _10713_);
  and (_28191_, _05315_, \oc8051_golden_model_1.ACC [5]);
  nor (_28192_, _28191_, _28181_);
  nor (_28193_, _28192_, _04500_);
  or (_28194_, _28193_, _28190_);
  and (_28195_, _28194_, _04868_);
  and (_28197_, _28177_, _03947_);
  nor (_28198_, _28197_, _28195_);
  nor (_28199_, _28198_, _03599_);
  nor (_28200_, _13035_, _10686_);
  nor (_28201_, _28200_, _28181_);
  nor (_28202_, _28201_, _04515_);
  or (_28203_, _28202_, _28199_);
  and (_28204_, _28203_, _03257_);
  not (_28205_, _28177_);
  nor (_28206_, _28205_, _03257_);
  or (_28208_, _28206_, _28204_);
  and (_28209_, _28208_, _04524_);
  and (_28210_, _10716_, _04079_);
  nor (_28211_, _28079_, _10713_);
  nor (_28212_, _28211_, _28210_);
  nor (_28213_, _28212_, _04524_);
  or (_28214_, _28213_, _28209_);
  and (_28215_, _28214_, _03611_);
  nor (_28216_, _28192_, _03611_);
  or (_28217_, _28216_, _28215_);
  and (_28219_, _28217_, _04650_);
  and (_28220_, _10673_, \oc8051_golden_model_1.SP [0]);
  nor (_28221_, _28055_, \oc8051_golden_model_1.SP [5]);
  nor (_28222_, _28221_, _28220_);
  and (_28223_, _28222_, _03510_);
  nor (_28224_, _28223_, _10729_);
  not (_28225_, _28224_);
  nor (_28226_, _28225_, _28219_);
  nor (_28227_, _28177_, _04856_);
  or (_28228_, _28227_, _07441_);
  nor (_28229_, _28228_, _28226_);
  nor (_28230_, _28229_, _28189_);
  and (_28231_, _06842_, _05315_);
  nor (_28232_, _28181_, _05970_);
  not (_28233_, _28232_);
  nor (_28234_, _28233_, _28231_);
  or (_28235_, _28234_, _03644_);
  nor (_28236_, _28235_, _28230_);
  nor (_28237_, _13139_, _10686_);
  nor (_28238_, _28237_, _28181_);
  nor (_28241_, _28238_, _03275_);
  or (_28242_, _28241_, _03650_);
  or (_28243_, _28242_, _28236_);
  and (_28244_, _06358_, _05315_);
  nor (_28245_, _28244_, _28181_);
  nand (_28246_, _28245_, _03650_);
  and (_28247_, _28246_, _28243_);
  nor (_28248_, _28247_, _03227_);
  and (_28249_, _28205_, _03227_);
  nor (_28250_, _28249_, _28248_);
  nor (_28252_, _28250_, _03649_);
  and (_28253_, _13154_, _05315_);
  or (_28254_, _28181_, _04591_);
  nor (_28255_, _28254_, _28253_);
  or (_28256_, _28255_, _03778_);
  nor (_28257_, _28256_, _28252_);
  nor (_28258_, _28257_, _28184_);
  nor (_28259_, _28258_, _03655_);
  nor (_28260_, _28181_, _05601_);
  not (_28261_, _28260_);
  nor (_28263_, _28245_, _04596_);
  and (_28264_, _28263_, _28261_);
  nor (_28265_, _28264_, _28259_);
  nor (_28266_, _28265_, _10777_);
  nor (_28267_, _28192_, _04594_);
  and (_28268_, _28267_, _28261_);
  nor (_28269_, _28268_, _28266_);
  and (_28270_, _28269_, _28180_);
  nor (_28271_, _13152_, _10686_);
  nor (_28272_, _28271_, _28181_);
  and (_28274_, _28272_, _03653_);
  nor (_28275_, _28274_, _28270_);
  nor (_28276_, _28275_, _03786_);
  nor (_28277_, _13159_, _10686_);
  or (_28278_, _28181_, _04606_);
  nor (_28279_, _28278_, _28277_);
  or (_28280_, _28279_, _03792_);
  nor (_28281_, _28280_, _28276_);
  nor (_28282_, _10715_, _10713_);
  nor (_28283_, _28282_, _10716_);
  nor (_28285_, _28283_, _10680_);
  or (_28286_, _28285_, _28281_);
  and (_28287_, _28286_, _06475_);
  and (_28288_, _28177_, _03248_);
  or (_28289_, _28288_, _28287_);
  and (_28290_, _28289_, _03522_);
  nor (_28291_, _28283_, _03522_);
  or (_28292_, _28291_, _28290_);
  and (_28293_, _28292_, _04260_);
  nor (_28294_, _28201_, _04260_);
  nor (_28296_, _28294_, _05047_);
  not (_28297_, _28296_);
  nor (_28298_, _28297_, _28293_);
  nor (_28299_, _28298_, _28178_);
  nor (_28300_, _28299_, _03816_);
  and (_28301_, _13217_, _05315_);
  nor (_28302_, _28301_, _28181_);
  and (_28303_, _28302_, _03816_);
  nor (_28304_, _28303_, _28300_);
  or (_28305_, _28304_, _43231_);
  or (_28307_, _43227_, \oc8051_golden_model_1.SP [5]);
  and (_28308_, _28307_, _41991_);
  and (_43553_, _28308_, _28305_);
  nor (_28309_, _05315_, _10712_);
  and (_28310_, _13374_, _05315_);
  nor (_28311_, _28310_, _28309_);
  nor (_28312_, _28311_, _04589_);
  and (_28313_, _06531_, _05315_);
  or (_28314_, _28313_, _28309_);
  and (_28315_, _28314_, _05969_);
  nor (_28317_, _04499_, _10712_);
  and (_28318_, _05315_, \oc8051_golden_model_1.ACC [6]);
  nor (_28319_, _28318_, _28309_);
  nor (_28320_, _28319_, _04500_);
  or (_28321_, _28320_, _28317_);
  and (_28322_, _28321_, _04868_);
  nor (_28323_, _10673_, \oc8051_golden_model_1.SP [6]);
  nor (_28324_, _28323_, _10674_);
  and (_28325_, _28324_, _03947_);
  nor (_28326_, _28325_, _28322_);
  nor (_28328_, _28326_, _03599_);
  nor (_28329_, _13235_, _10686_);
  nor (_28330_, _28329_, _28309_);
  nor (_28331_, _28330_, _04515_);
  or (_28332_, _28331_, _28328_);
  and (_28333_, _28332_, _03257_);
  not (_28334_, _28324_);
  nor (_28335_, _28334_, _03257_);
  or (_28336_, _28335_, _28333_);
  and (_28337_, _28336_, _04524_);
  nor (_28339_, _28210_, _10712_);
  nor (_28340_, _28339_, _10718_);
  nor (_28341_, _28340_, _04524_);
  or (_28342_, _28341_, _28337_);
  and (_28343_, _28342_, _03611_);
  nor (_28344_, _28319_, _03611_);
  or (_28345_, _28344_, _28343_);
  and (_28346_, _28345_, _04650_);
  nor (_28347_, _28220_, \oc8051_golden_model_1.SP [6]);
  nor (_28348_, _28347_, _10730_);
  and (_28350_, _28348_, _03510_);
  nor (_28351_, _28350_, _28346_);
  nor (_28352_, _28351_, _10729_);
  nor (_28353_, _28334_, _04856_);
  nor (_28354_, _28353_, _07441_);
  not (_28355_, _28354_);
  nor (_28356_, _28355_, _28352_);
  not (_28357_, _28309_);
  nor (_28358_, _05442_, _10686_);
  nor (_28359_, _28358_, _06889_);
  and (_28361_, _28359_, _28357_);
  or (_28362_, _28361_, _05969_);
  nor (_28363_, _28362_, _28356_);
  or (_28364_, _28363_, _28315_);
  and (_28365_, _28364_, _03275_);
  nor (_28366_, _13356_, _10686_);
  nor (_28367_, _28366_, _28309_);
  nor (_28368_, _28367_, _03275_);
  or (_28369_, _28368_, _03650_);
  or (_28370_, _28369_, _28365_);
  and (_28372_, _13363_, _05315_);
  nor (_28373_, _28372_, _28309_);
  nand (_28374_, _28373_, _03650_);
  and (_28375_, _28374_, _28370_);
  nor (_28376_, _28375_, _03227_);
  and (_28377_, _28334_, _03227_);
  nor (_28378_, _28377_, _28376_);
  nor (_28379_, _28378_, _03649_);
  and (_28380_, _13245_, _05315_);
  or (_28381_, _28309_, _04591_);
  nor (_28383_, _28381_, _28380_);
  or (_28384_, _28383_, _03778_);
  nor (_28385_, _28384_, _28379_);
  nor (_28386_, _28385_, _28312_);
  nor (_28387_, _28386_, _03655_);
  and (_28388_, _28357_, _05490_);
  not (_28389_, _28388_);
  nor (_28390_, _28373_, _04596_);
  and (_28391_, _28390_, _28389_);
  nor (_28392_, _28391_, _28387_);
  nor (_28394_, _28392_, _10777_);
  and (_28395_, _28324_, _03238_);
  or (_28396_, _28388_, _04594_);
  nor (_28397_, _28396_, _28319_);
  nor (_28398_, _28397_, _28395_);
  and (_28399_, _28398_, _04608_);
  not (_28400_, _28399_);
  nor (_28401_, _28400_, _28394_);
  nor (_28402_, _13243_, _10686_);
  nor (_28403_, _28402_, _28309_);
  and (_28405_, _28403_, _03653_);
  nor (_28406_, _28405_, _28401_);
  and (_28407_, _28406_, _04606_);
  nor (_28408_, _13373_, _10686_);
  nor (_28409_, _28408_, _28309_);
  nor (_28410_, _28409_, _04606_);
  or (_28411_, _28410_, _28407_);
  and (_28412_, _28411_, _10680_);
  nor (_28413_, _10716_, _10712_);
  nor (_28414_, _28413_, _10717_);
  not (_28415_, _28414_);
  nor (_28416_, _28415_, _03248_);
  nor (_28417_, _28416_, _10796_);
  nor (_28418_, _28417_, _28412_);
  and (_28419_, _28334_, _03248_);
  or (_28420_, _28419_, _03521_);
  nor (_28421_, _28420_, _28418_);
  and (_28422_, _28415_, _03521_);
  or (_28423_, _28422_, _03809_);
  nor (_28424_, _28423_, _28421_);
  and (_28427_, _28330_, _03809_);
  nor (_28428_, _28427_, _05047_);
  not (_28429_, _28428_);
  nor (_28430_, _28429_, _28424_);
  nor (_28431_, _28334_, _04625_);
  nor (_28432_, _28431_, _03816_);
  not (_28433_, _28432_);
  nor (_28434_, _28433_, _28430_);
  and (_28435_, _13425_, _05315_);
  or (_28436_, _28309_, _03820_);
  nor (_28438_, _28436_, _28435_);
  nor (_28439_, _28438_, _28434_);
  or (_28440_, _28439_, _43231_);
  or (_28441_, _43227_, \oc8051_golden_model_1.SP [6]);
  and (_28442_, _28441_, _41991_);
  and (_43554_, _28442_, _28440_);
  not (_28443_, \oc8051_golden_model_1.TCON [0]);
  nor (_28444_, _05353_, _28443_);
  nor (_28445_, _05744_, _10824_);
  nor (_28446_, _28445_, _28444_);
  and (_28448_, _28446_, _03816_);
  and (_28449_, _12145_, _05353_);
  nor (_28450_, _28449_, _28444_);
  nor (_28451_, _28450_, _04589_);
  and (_28452_, _05353_, _06366_);
  nor (_28453_, _28452_, _28444_);
  and (_28454_, _28453_, _03650_);
  and (_28455_, _05353_, _04491_);
  nor (_28456_, _28455_, _28444_);
  and (_28457_, _28456_, _07441_);
  and (_28459_, _05353_, \oc8051_golden_model_1.ACC [0]);
  nor (_28460_, _28459_, _28444_);
  nor (_28461_, _28460_, _04500_);
  nor (_28462_, _04499_, _28443_);
  or (_28463_, _28462_, _28461_);
  and (_28464_, _28463_, _04515_);
  nor (_28465_, _28446_, _04515_);
  or (_28466_, _28465_, _28464_);
  and (_28467_, _28466_, _03516_);
  nor (_28468_, _05997_, _28443_);
  and (_28470_, _12035_, _05997_);
  nor (_28471_, _28470_, _28468_);
  nor (_28472_, _28471_, _03516_);
  nor (_28473_, _28472_, _28467_);
  nor (_28474_, _28473_, _03597_);
  nor (_28475_, _28456_, _04524_);
  or (_28476_, _28475_, _28474_);
  and (_28477_, _28476_, _03611_);
  nor (_28478_, _28460_, _03611_);
  or (_28479_, _28478_, _28477_);
  and (_28481_, _28479_, _03512_);
  and (_28482_, _28444_, _03511_);
  or (_28483_, _28482_, _28481_);
  and (_28484_, _28483_, _03505_);
  nor (_28485_, _28446_, _03505_);
  or (_28486_, _28485_, _28484_);
  and (_28487_, _28486_, _03501_);
  nor (_28488_, _12066_, _10861_);
  nor (_28489_, _28488_, _28468_);
  nor (_28490_, _28489_, _03501_);
  or (_28492_, _28490_, _07441_);
  nor (_28493_, _28492_, _28487_);
  nor (_28494_, _28493_, _28457_);
  nor (_28495_, _28494_, _05969_);
  and (_28496_, _06836_, _05353_);
  nor (_28497_, _28444_, _05970_);
  not (_28498_, _28497_);
  nor (_28499_, _28498_, _28496_);
  or (_28500_, _28499_, _03644_);
  nor (_28501_, _28500_, _28495_);
  nor (_28503_, _12129_, _10824_);
  nor (_28504_, _28503_, _28444_);
  nor (_28505_, _28504_, _03275_);
  or (_28506_, _28505_, _03650_);
  nor (_28507_, _28506_, _28501_);
  nor (_28508_, _28507_, _28454_);
  or (_28509_, _28508_, _03649_);
  and (_28510_, _12019_, _05353_);
  or (_28511_, _28510_, _28444_);
  or (_28512_, _28511_, _04591_);
  and (_28514_, _28512_, _04589_);
  and (_28515_, _28514_, _28509_);
  nor (_28516_, _28515_, _28451_);
  nor (_28517_, _28516_, _03655_);
  or (_28518_, _28453_, _04596_);
  nor (_28519_, _28518_, _28445_);
  nor (_28520_, _28519_, _28517_);
  nor (_28521_, _28520_, _03773_);
  and (_28522_, _12144_, _05353_);
  or (_28523_, _28522_, _28444_);
  and (_28525_, _28523_, _03773_);
  or (_28526_, _28525_, _28521_);
  and (_28527_, _28526_, _04608_);
  nor (_28528_, _12017_, _10824_);
  nor (_28529_, _28528_, _28444_);
  nor (_28530_, _28529_, _04608_);
  or (_28531_, _28530_, _28527_);
  and (_28532_, _28531_, _04606_);
  nor (_28533_, _12015_, _10824_);
  nor (_28534_, _28533_, _28444_);
  nor (_28536_, _28534_, _04606_);
  or (_28537_, _28536_, _28532_);
  and (_28538_, _28537_, _04260_);
  nor (_28539_, _28446_, _04260_);
  or (_28540_, _28539_, _28538_);
  and (_28541_, _28540_, _03206_);
  and (_28542_, _28444_, _03205_);
  nor (_28543_, _28542_, _03816_);
  not (_28544_, _28543_);
  nor (_28545_, _28544_, _28541_);
  nor (_28547_, _28545_, _28448_);
  or (_28548_, _28547_, _43231_);
  or (_28549_, _43227_, \oc8051_golden_model_1.TCON [0]);
  and (_28550_, _28549_, _41991_);
  and (_43555_, _28550_, _28548_);
  and (_28551_, _10824_, \oc8051_golden_model_1.TCON [1]);
  and (_28552_, _05353_, _05898_);
  or (_28553_, _28552_, _28551_);
  or (_28554_, _28553_, _04524_);
  or (_28555_, _05353_, \oc8051_golden_model_1.TCON [1]);
  and (_28557_, _12234_, _05353_);
  not (_28558_, _28557_);
  and (_28559_, _28558_, _28555_);
  or (_28560_, _28559_, _04515_);
  nand (_28561_, _05353_, _03320_);
  and (_28562_, _28561_, _28555_);
  and (_28563_, _28562_, _04499_);
  and (_28564_, _04500_, \oc8051_golden_model_1.TCON [1]);
  or (_28565_, _28564_, _03599_);
  or (_28566_, _28565_, _28563_);
  and (_28568_, _28566_, _03516_);
  and (_28569_, _28568_, _28560_);
  and (_28570_, _10861_, \oc8051_golden_model_1.TCON [1]);
  and (_28571_, _12238_, _05997_);
  or (_28572_, _28571_, _28570_);
  and (_28573_, _28572_, _03515_);
  or (_28574_, _28573_, _03597_);
  or (_28575_, _28574_, _28569_);
  and (_28576_, _28575_, _28554_);
  or (_28577_, _28576_, _03603_);
  or (_28579_, _28562_, _03611_);
  and (_28580_, _28579_, _03512_);
  and (_28581_, _28580_, _28577_);
  and (_28582_, _12224_, _05997_);
  or (_28583_, _28582_, _28570_);
  and (_28584_, _28583_, _03511_);
  or (_28585_, _28584_, _03504_);
  or (_28586_, _28585_, _28581_);
  and (_28587_, _28571_, _12253_);
  or (_28588_, _28570_, _03505_);
  or (_28590_, _28588_, _28587_);
  and (_28591_, _28590_, _28586_);
  and (_28592_, _28591_, _03501_);
  nor (_28593_, _12270_, _10861_);
  or (_28594_, _28570_, _28593_);
  and (_28595_, _28594_, _03500_);
  or (_28596_, _28595_, _07441_);
  or (_28597_, _28596_, _28592_);
  or (_28598_, _28553_, _06889_);
  and (_28599_, _28598_, _28597_);
  or (_28601_, _28599_, _05969_);
  and (_28602_, _06835_, _05353_);
  or (_28603_, _28551_, _05970_);
  or (_28604_, _28603_, _28602_);
  and (_28605_, _28604_, _03275_);
  and (_28606_, _28605_, _28601_);
  nor (_28607_, _12330_, _10824_);
  or (_28608_, _28607_, _28551_);
  and (_28609_, _28608_, _03644_);
  or (_28610_, _28609_, _28606_);
  and (_28612_, _28610_, _03651_);
  or (_28613_, _12220_, _10824_);
  and (_28614_, _28613_, _03649_);
  nand (_28615_, _05353_, _04347_);
  and (_28616_, _28615_, _03650_);
  or (_28617_, _28616_, _28614_);
  and (_28618_, _28617_, _28555_);
  or (_28619_, _28618_, _28612_);
  and (_28620_, _28619_, _04589_);
  or (_28621_, _12347_, _10824_);
  and (_28623_, _28555_, _03778_);
  and (_28624_, _28623_, _28621_);
  or (_28625_, _28624_, _28620_);
  and (_28626_, _28625_, _04596_);
  or (_28627_, _12219_, _10824_);
  and (_28628_, _28555_, _03655_);
  and (_28629_, _28628_, _28627_);
  or (_28630_, _28629_, _28626_);
  and (_28631_, _28630_, _04594_);
  or (_28632_, _28551_, _05699_);
  and (_28634_, _28562_, _03773_);
  and (_28635_, _28634_, _28632_);
  or (_28636_, _28635_, _28631_);
  and (_28637_, _28636_, _03787_);
  or (_28638_, _28615_, _05699_);
  and (_28639_, _28555_, _03653_);
  and (_28640_, _28639_, _28638_);
  or (_28641_, _28561_, _05699_);
  and (_28642_, _28555_, _03786_);
  and (_28643_, _28642_, _28641_);
  or (_28645_, _28643_, _03809_);
  or (_28646_, _28645_, _28640_);
  or (_28647_, _28646_, _28637_);
  or (_28648_, _28559_, _04260_);
  and (_28649_, _28648_, _03206_);
  and (_28650_, _28649_, _28647_);
  and (_28651_, _28583_, _03205_);
  or (_28652_, _28651_, _03816_);
  or (_28653_, _28652_, _28650_);
  or (_28654_, _28551_, _03820_);
  or (_28656_, _28654_, _28557_);
  and (_28657_, _28656_, _28653_);
  and (_28658_, _28657_, _43227_);
  nor (_28659_, \oc8051_golden_model_1.TCON [1], rst);
  nor (_28660_, _28659_, _00000_);
  or (_43556_, _28660_, _28658_);
  not (_28661_, \oc8051_golden_model_1.TCON [2]);
  nor (_28662_, _05353_, _28661_);
  and (_28663_, _05353_, _06414_);
  nor (_28664_, _28663_, _28662_);
  and (_28666_, _28664_, _03650_);
  nor (_28667_, _10824_, _05130_);
  nor (_28668_, _28667_, _28662_);
  and (_28669_, _28668_, _07441_);
  nor (_28670_, _28668_, _04524_);
  nor (_28671_, _05997_, _28661_);
  and (_28672_, _12416_, _05997_);
  nor (_28673_, _28672_, _28671_);
  and (_28674_, _28673_, _03515_);
  nor (_28675_, _12430_, _10824_);
  nor (_28677_, _28675_, _28662_);
  nor (_28678_, _28677_, _04515_);
  nor (_28679_, _04499_, _28661_);
  and (_28680_, _05353_, \oc8051_golden_model_1.ACC [2]);
  nor (_28681_, _28680_, _28662_);
  nor (_28682_, _28681_, _04500_);
  nor (_28683_, _28682_, _28679_);
  nor (_28684_, _28683_, _03599_);
  or (_28685_, _28684_, _03515_);
  nor (_28686_, _28685_, _28678_);
  nor (_28688_, _28686_, _28674_);
  and (_28689_, _28688_, _04524_);
  or (_28690_, _28689_, _28670_);
  and (_28691_, _28690_, _03611_);
  nor (_28692_, _28681_, _03611_);
  or (_28693_, _28692_, _28691_);
  and (_28694_, _28693_, _03512_);
  and (_28695_, _12414_, _05997_);
  nor (_28696_, _28695_, _28671_);
  nor (_28697_, _28696_, _03512_);
  or (_28699_, _28697_, _03504_);
  or (_28700_, _28699_, _28694_);
  nor (_28701_, _28671_, _12447_);
  nor (_28702_, _28701_, _28673_);
  or (_28703_, _28702_, _03505_);
  and (_28704_, _28703_, _03501_);
  and (_28705_, _28704_, _28700_);
  nor (_28706_, _12465_, _10861_);
  nor (_28707_, _28706_, _28671_);
  nor (_28708_, _28707_, _03501_);
  nor (_28710_, _28708_, _07441_);
  not (_28711_, _28710_);
  nor (_28712_, _28711_, _28705_);
  nor (_28713_, _28712_, _28669_);
  nor (_28714_, _28713_, _05969_);
  and (_28715_, _06839_, _05353_);
  nor (_28716_, _28662_, _05970_);
  not (_28717_, _28716_);
  nor (_28718_, _28717_, _28715_);
  or (_28719_, _28718_, _03644_);
  nor (_28721_, _28719_, _28714_);
  nor (_28722_, _12524_, _10824_);
  nor (_28723_, _28662_, _28722_);
  nor (_28724_, _28723_, _03275_);
  or (_28725_, _28724_, _03650_);
  nor (_28726_, _28725_, _28721_);
  nor (_28727_, _28726_, _28666_);
  or (_28728_, _28727_, _03649_);
  and (_28729_, _12538_, _05353_);
  or (_28730_, _28729_, _28662_);
  or (_28732_, _28730_, _04591_);
  and (_28733_, _28732_, _04589_);
  and (_28734_, _28733_, _28728_);
  and (_28735_, _12544_, _05353_);
  nor (_28736_, _28735_, _28662_);
  nor (_28737_, _28736_, _04589_);
  nor (_28738_, _28737_, _28734_);
  nor (_28739_, _28738_, _03655_);
  nor (_28740_, _28662_, _05793_);
  not (_28741_, _28740_);
  nor (_28743_, _28664_, _04596_);
  and (_28744_, _28743_, _28741_);
  nor (_28745_, _28744_, _28739_);
  nor (_28746_, _28745_, _03773_);
  nor (_28747_, _28681_, _04594_);
  and (_28748_, _28747_, _28741_);
  or (_28749_, _28748_, _28746_);
  and (_28750_, _28749_, _04608_);
  nor (_28751_, _12537_, _10824_);
  nor (_28752_, _28751_, _28662_);
  nor (_28754_, _28752_, _04608_);
  or (_28755_, _28754_, _28750_);
  and (_28756_, _28755_, _04606_);
  nor (_28757_, _12543_, _10824_);
  nor (_28758_, _28757_, _28662_);
  nor (_28759_, _28758_, _04606_);
  or (_28760_, _28759_, _28756_);
  and (_28761_, _28760_, _04260_);
  nor (_28762_, _28677_, _04260_);
  or (_28763_, _28762_, _28761_);
  and (_28765_, _28763_, _03206_);
  nor (_28766_, _28696_, _03206_);
  nor (_28767_, _28766_, _03816_);
  not (_28768_, _28767_);
  nor (_28769_, _28768_, _28765_);
  and (_28770_, _12600_, _05353_);
  or (_28771_, _28662_, _03820_);
  nor (_28772_, _28771_, _28770_);
  nor (_28773_, _28772_, _28769_);
  or (_28774_, _28773_, _43231_);
  or (_28776_, _43227_, \oc8051_golden_model_1.TCON [2]);
  and (_28777_, _28776_, _41991_);
  and (_43557_, _28777_, _28774_);
  not (_28778_, \oc8051_golden_model_1.TCON [3]);
  nor (_28779_, _05353_, _28778_);
  and (_28780_, _05353_, _06347_);
  nor (_28781_, _28780_, _28779_);
  and (_28782_, _28781_, _03650_);
  nor (_28783_, _10824_, _04944_);
  nor (_28784_, _28783_, _28779_);
  and (_28786_, _28784_, _07441_);
  and (_28787_, _05353_, \oc8051_golden_model_1.ACC [3]);
  nor (_28788_, _28787_, _28779_);
  nor (_28789_, _28788_, _04500_);
  nor (_28790_, _04499_, _28778_);
  or (_28791_, _28790_, _28789_);
  and (_28792_, _28791_, _04515_);
  nor (_28793_, _12625_, _10824_);
  nor (_28794_, _28793_, _28779_);
  nor (_28795_, _28794_, _04515_);
  or (_28797_, _28795_, _28792_);
  and (_28798_, _28797_, _03516_);
  nor (_28799_, _05997_, _28778_);
  and (_28800_, _12638_, _05997_);
  nor (_28801_, _28800_, _28799_);
  nor (_28802_, _28801_, _03516_);
  or (_28803_, _28802_, _03597_);
  or (_28804_, _28803_, _28798_);
  nand (_28805_, _28784_, _03597_);
  and (_28806_, _28805_, _28804_);
  and (_28808_, _28806_, _03611_);
  nor (_28809_, _28788_, _03611_);
  or (_28810_, _28809_, _28808_);
  and (_28811_, _28810_, _03512_);
  and (_28812_, _12622_, _05997_);
  nor (_28813_, _28812_, _28799_);
  nor (_28814_, _28813_, _03512_);
  or (_28815_, _28814_, _28811_);
  and (_28816_, _28815_, _03505_);
  nor (_28817_, _28799_, _12653_);
  nor (_28818_, _28817_, _28801_);
  and (_28819_, _28818_, _03504_);
  or (_28820_, _28819_, _28816_);
  and (_28821_, _28820_, _03501_);
  nor (_28822_, _12671_, _10861_);
  nor (_28823_, _28822_, _28799_);
  nor (_28824_, _28823_, _03501_);
  nor (_28825_, _28824_, _07441_);
  not (_28826_, _28825_);
  nor (_28827_, _28826_, _28821_);
  nor (_28829_, _28827_, _28786_);
  nor (_28830_, _28829_, _05969_);
  and (_28831_, _06838_, _05353_);
  nor (_28832_, _28779_, _05970_);
  not (_28833_, _28832_);
  nor (_28834_, _28833_, _28831_);
  or (_28835_, _28834_, _03644_);
  nor (_28836_, _28835_, _28830_);
  nor (_28837_, _12731_, _10824_);
  nor (_28838_, _28779_, _28837_);
  nor (_28840_, _28838_, _03275_);
  or (_28841_, _28840_, _03650_);
  nor (_28842_, _28841_, _28836_);
  nor (_28843_, _28842_, _28782_);
  or (_28844_, _28843_, _03649_);
  and (_28845_, _12746_, _05353_);
  or (_28846_, _28845_, _28779_);
  or (_28847_, _28846_, _04591_);
  and (_28848_, _28847_, _04589_);
  and (_28849_, _28848_, _28844_);
  and (_28851_, _12619_, _05353_);
  nor (_28852_, _28851_, _28779_);
  nor (_28853_, _28852_, _04589_);
  nor (_28854_, _28853_, _28849_);
  nor (_28855_, _28854_, _03655_);
  nor (_28856_, _28779_, _05650_);
  not (_28857_, _28856_);
  nor (_28858_, _28781_, _04596_);
  and (_28859_, _28858_, _28857_);
  nor (_28860_, _28859_, _28855_);
  nor (_28862_, _28860_, _03773_);
  nor (_28863_, _28788_, _04594_);
  and (_28864_, _28863_, _28857_);
  or (_28865_, _28864_, _28862_);
  and (_28866_, _28865_, _04608_);
  nor (_28867_, _12745_, _10824_);
  nor (_28868_, _28867_, _28779_);
  nor (_28869_, _28868_, _04608_);
  or (_28870_, _28869_, _28866_);
  and (_28871_, _28870_, _04606_);
  nor (_28873_, _12618_, _10824_);
  nor (_28874_, _28873_, _28779_);
  nor (_28875_, _28874_, _04606_);
  or (_28876_, _28875_, _28871_);
  and (_28877_, _28876_, _04260_);
  nor (_28878_, _28794_, _04260_);
  or (_28879_, _28878_, _28877_);
  and (_28880_, _28879_, _03206_);
  nor (_28881_, _28813_, _03206_);
  or (_28882_, _28881_, _28880_);
  and (_28884_, _28882_, _03820_);
  and (_28885_, _12806_, _05353_);
  nor (_28886_, _28885_, _28779_);
  nor (_28887_, _28886_, _03820_);
  or (_28888_, _28887_, _28884_);
  or (_28889_, _28888_, _43231_);
  or (_28890_, _43227_, \oc8051_golden_model_1.TCON [3]);
  and (_28891_, _28890_, _41991_);
  and (_43560_, _28891_, _28889_);
  not (_28892_, \oc8051_golden_model_1.TCON [4]);
  nor (_28894_, _05353_, _28892_);
  nor (_28895_, _05840_, _10824_);
  nor (_28896_, _28895_, _28894_);
  and (_28897_, _28896_, _07441_);
  nor (_28898_, _05997_, _28892_);
  and (_28899_, _12853_, _05997_);
  nor (_28900_, _28899_, _28898_);
  nor (_28901_, _28900_, _03512_);
  and (_28902_, _05353_, \oc8051_golden_model_1.ACC [4]);
  nor (_28903_, _28902_, _28894_);
  nor (_28905_, _28903_, _04500_);
  nor (_28906_, _04499_, _28892_);
  or (_28907_, _28906_, _28905_);
  and (_28908_, _28907_, _04515_);
  nor (_28909_, _12820_, _10824_);
  nor (_28910_, _28909_, _28894_);
  nor (_28911_, _28910_, _04515_);
  or (_28912_, _28911_, _28908_);
  and (_28913_, _28912_, _03516_);
  and (_28914_, _12830_, _05997_);
  nor (_28916_, _28914_, _28898_);
  nor (_28917_, _28916_, _03516_);
  or (_28918_, _28917_, _03597_);
  or (_28919_, _28918_, _28913_);
  nand (_28920_, _28896_, _03597_);
  and (_28921_, _28920_, _28919_);
  and (_28922_, _28921_, _03611_);
  nor (_28923_, _28903_, _03611_);
  or (_28924_, _28923_, _28922_);
  and (_28925_, _28924_, _03512_);
  nor (_28927_, _28925_, _28901_);
  nor (_28928_, _28927_, _03504_);
  nor (_28929_, _28898_, _12860_);
  or (_28930_, _28916_, _03505_);
  nor (_28931_, _28930_, _28929_);
  nor (_28932_, _28931_, _28928_);
  nor (_28933_, _28932_, _03500_);
  nor (_28934_, _12828_, _10861_);
  nor (_28935_, _28934_, _28898_);
  nor (_28936_, _28935_, _03501_);
  nor (_28938_, _28936_, _07441_);
  not (_28939_, _28938_);
  nor (_28940_, _28939_, _28933_);
  nor (_28941_, _28940_, _28897_);
  nor (_28942_, _28941_, _05969_);
  and (_28943_, _06843_, _05353_);
  nor (_28944_, _28894_, _05970_);
  not (_28945_, _28944_);
  nor (_28946_, _28945_, _28943_);
  nor (_28947_, _28946_, _03644_);
  not (_28948_, _28947_);
  nor (_28949_, _28948_, _28942_);
  nor (_28950_, _12936_, _10824_);
  nor (_28951_, _28950_, _28894_);
  nor (_28952_, _28951_, _03275_);
  or (_28953_, _28952_, _08861_);
  or (_28954_, _28953_, _28949_);
  and (_28955_, _12951_, _05353_);
  or (_28956_, _28894_, _04591_);
  or (_28957_, _28956_, _28955_);
  and (_28960_, _06375_, _05353_);
  nor (_28961_, _28960_, _28894_);
  and (_28962_, _28961_, _03650_);
  nor (_28963_, _28962_, _03778_);
  and (_28964_, _28963_, _28957_);
  and (_28965_, _28964_, _28954_);
  and (_28966_, _12957_, _05353_);
  nor (_28967_, _28966_, _28894_);
  nor (_28968_, _28967_, _04589_);
  nor (_28969_, _28968_, _28965_);
  nor (_28971_, _28969_, _03655_);
  nor (_28972_, _28894_, _05889_);
  not (_28973_, _28972_);
  nor (_28974_, _28961_, _04596_);
  and (_28975_, _28974_, _28973_);
  nor (_28976_, _28975_, _28971_);
  nor (_28977_, _28976_, _03773_);
  nor (_28978_, _28903_, _04594_);
  and (_28979_, _28978_, _28973_);
  or (_28980_, _28979_, _28977_);
  and (_28982_, _28980_, _04608_);
  nor (_28983_, _12949_, _10824_);
  nor (_28984_, _28983_, _28894_);
  nor (_28985_, _28984_, _04608_);
  or (_28986_, _28985_, _28982_);
  and (_28987_, _28986_, _04606_);
  nor (_28988_, _12956_, _10824_);
  nor (_28989_, _28988_, _28894_);
  nor (_28990_, _28989_, _04606_);
  or (_28991_, _28990_, _28987_);
  and (_28993_, _28991_, _04260_);
  nor (_28994_, _28910_, _04260_);
  or (_28995_, _28994_, _28993_);
  and (_28996_, _28995_, _03206_);
  nor (_28997_, _28900_, _03206_);
  or (_28998_, _28997_, _28996_);
  and (_28999_, _28998_, _03820_);
  and (_29000_, _13013_, _05353_);
  nor (_29001_, _29000_, _28894_);
  nor (_29002_, _29001_, _03820_);
  or (_29004_, _29002_, _28999_);
  or (_29005_, _29004_, _43231_);
  or (_29006_, _43227_, \oc8051_golden_model_1.TCON [4]);
  and (_29007_, _29006_, _41991_);
  and (_43561_, _29007_, _29005_);
  not (_29008_, \oc8051_golden_model_1.TCON [5]);
  nor (_29009_, _05353_, _29008_);
  and (_29010_, _06842_, _05353_);
  or (_29011_, _29010_, _29009_);
  and (_29012_, _29011_, _05969_);
  and (_29014_, _05353_, \oc8051_golden_model_1.ACC [5]);
  nor (_29015_, _29014_, _29009_);
  nor (_29016_, _29015_, _04500_);
  nor (_29017_, _04499_, _29008_);
  or (_29018_, _29017_, _29016_);
  and (_29019_, _29018_, _04515_);
  nor (_29020_, _13035_, _10824_);
  nor (_29021_, _29020_, _29009_);
  nor (_29022_, _29021_, _04515_);
  or (_29023_, _29022_, _29019_);
  and (_29025_, _29023_, _03516_);
  nor (_29026_, _05997_, _29008_);
  and (_29027_, _13051_, _05997_);
  nor (_29028_, _29027_, _29026_);
  nor (_29029_, _29028_, _03516_);
  or (_29030_, _29029_, _03597_);
  or (_29031_, _29030_, _29025_);
  nor (_29032_, _05552_, _10824_);
  nor (_29033_, _29032_, _29009_);
  nand (_29034_, _29033_, _03597_);
  and (_29036_, _29034_, _29031_);
  and (_29037_, _29036_, _03611_);
  nor (_29038_, _29015_, _03611_);
  or (_29039_, _29038_, _29037_);
  and (_29040_, _29039_, _03512_);
  and (_29041_, _13032_, _05997_);
  nor (_29042_, _29041_, _29026_);
  nor (_29043_, _29042_, _03512_);
  or (_29044_, _29043_, _03504_);
  or (_29045_, _29044_, _29040_);
  nor (_29047_, _29026_, _13066_);
  nor (_29048_, _29047_, _29028_);
  or (_29049_, _29048_, _03505_);
  and (_29050_, _29049_, _03501_);
  and (_29051_, _29050_, _29045_);
  nor (_29052_, _13030_, _10861_);
  nor (_29053_, _29052_, _29026_);
  nor (_29054_, _29053_, _03501_);
  nor (_29055_, _29054_, _07441_);
  not (_29056_, _29055_);
  nor (_29058_, _29056_, _29051_);
  and (_29059_, _29033_, _07441_);
  or (_29060_, _29059_, _05969_);
  nor (_29061_, _29060_, _29058_);
  or (_29062_, _29061_, _29012_);
  and (_29063_, _29062_, _03275_);
  nor (_29064_, _13139_, _10824_);
  nor (_29065_, _29064_, _29009_);
  nor (_29066_, _29065_, _03275_);
  or (_29067_, _29066_, _08861_);
  or (_29069_, _29067_, _29063_);
  and (_29070_, _13154_, _05353_);
  or (_29071_, _29009_, _04591_);
  or (_29072_, _29071_, _29070_);
  and (_29073_, _06358_, _05353_);
  nor (_29074_, _29073_, _29009_);
  and (_29075_, _29074_, _03650_);
  nor (_29076_, _29075_, _03778_);
  and (_29077_, _29076_, _29072_);
  and (_29078_, _29077_, _29069_);
  and (_29080_, _13160_, _05353_);
  nor (_29081_, _29080_, _29009_);
  nor (_29082_, _29081_, _04589_);
  nor (_29083_, _29082_, _29078_);
  nor (_29084_, _29083_, _03655_);
  nor (_29085_, _29009_, _05601_);
  not (_29086_, _29085_);
  nor (_29087_, _29074_, _04596_);
  and (_29088_, _29087_, _29086_);
  nor (_29089_, _29088_, _29084_);
  nor (_29091_, _29089_, _03773_);
  nor (_29092_, _29015_, _04594_);
  and (_29093_, _29092_, _29086_);
  nor (_29094_, _29093_, _03653_);
  not (_29095_, _29094_);
  nor (_29096_, _29095_, _29091_);
  nor (_29097_, _13152_, _10824_);
  or (_29098_, _29009_, _04608_);
  nor (_29099_, _29098_, _29097_);
  or (_29100_, _29099_, _03786_);
  nor (_29102_, _29100_, _29096_);
  nor (_29103_, _13159_, _10824_);
  nor (_29104_, _29103_, _29009_);
  nor (_29105_, _29104_, _04606_);
  or (_29106_, _29105_, _29102_);
  and (_29107_, _29106_, _04260_);
  nor (_29108_, _29021_, _04260_);
  or (_29109_, _29108_, _29107_);
  and (_29110_, _29109_, _03206_);
  nor (_29111_, _29042_, _03206_);
  or (_29113_, _29111_, _29110_);
  and (_29114_, _29113_, _03820_);
  and (_29115_, _13217_, _05353_);
  nor (_29116_, _29115_, _29009_);
  nor (_29117_, _29116_, _03820_);
  or (_29118_, _29117_, _29114_);
  or (_29119_, _29118_, _43231_);
  or (_29120_, _43227_, \oc8051_golden_model_1.TCON [5]);
  and (_29121_, _29120_, _41991_);
  and (_43562_, _29121_, _29119_);
  not (_29123_, \oc8051_golden_model_1.TCON [6]);
  nor (_29124_, _05353_, _29123_);
  and (_29125_, _06531_, _05353_);
  or (_29126_, _29125_, _29124_);
  and (_29127_, _29126_, _05969_);
  and (_29128_, _05353_, \oc8051_golden_model_1.ACC [6]);
  nor (_29129_, _29128_, _29124_);
  nor (_29130_, _29129_, _04500_);
  nor (_29131_, _04499_, _29123_);
  or (_29132_, _29131_, _29130_);
  and (_29134_, _29132_, _04515_);
  nor (_29135_, _13235_, _10824_);
  nor (_29136_, _29135_, _29124_);
  nor (_29137_, _29136_, _04515_);
  or (_29138_, _29137_, _29134_);
  and (_29139_, _29138_, _03516_);
  nor (_29140_, _05997_, _29123_);
  and (_29141_, _13266_, _05997_);
  nor (_29142_, _29141_, _29140_);
  nor (_29143_, _29142_, _03516_);
  or (_29145_, _29143_, _03597_);
  or (_29146_, _29145_, _29139_);
  nor (_29147_, _05442_, _10824_);
  nor (_29148_, _29147_, _29124_);
  nand (_29149_, _29148_, _03597_);
  and (_29150_, _29149_, _29146_);
  and (_29151_, _29150_, _03611_);
  nor (_29152_, _29129_, _03611_);
  or (_29153_, _29152_, _29151_);
  and (_29154_, _29153_, _03512_);
  and (_29156_, _13251_, _05997_);
  nor (_29157_, _29156_, _29140_);
  nor (_29158_, _29157_, _03512_);
  or (_29159_, _29158_, _29154_);
  and (_29160_, _29159_, _03505_);
  nor (_29161_, _29140_, _13281_);
  nor (_29162_, _29161_, _29142_);
  and (_29163_, _29162_, _03504_);
  or (_29164_, _29163_, _29160_);
  and (_29165_, _29164_, _03501_);
  nor (_29167_, _13249_, _10861_);
  nor (_29168_, _29167_, _29140_);
  nor (_29169_, _29168_, _03501_);
  nor (_29170_, _29169_, _07441_);
  not (_29171_, _29170_);
  nor (_29172_, _29171_, _29165_);
  and (_29173_, _29148_, _07441_);
  or (_29174_, _29173_, _05969_);
  nor (_29175_, _29174_, _29172_);
  or (_29176_, _29175_, _29127_);
  and (_29178_, _29176_, _03275_);
  nor (_29179_, _13356_, _10824_);
  nor (_29180_, _29179_, _29124_);
  nor (_29181_, _29180_, _03275_);
  or (_29182_, _29181_, _08861_);
  or (_29183_, _29182_, _29178_);
  and (_29184_, _13245_, _05353_);
  or (_29185_, _29124_, _04591_);
  or (_29186_, _29185_, _29184_);
  and (_29187_, _13363_, _05353_);
  nor (_29189_, _29187_, _29124_);
  and (_29190_, _29189_, _03650_);
  nor (_29191_, _29190_, _03778_);
  and (_29192_, _29191_, _29186_);
  and (_29193_, _29192_, _29183_);
  and (_29194_, _13374_, _05353_);
  nor (_29195_, _29194_, _29124_);
  nor (_29196_, _29195_, _04589_);
  nor (_29197_, _29196_, _29193_);
  nor (_29198_, _29197_, _03655_);
  nor (_29200_, _29124_, _05491_);
  not (_29201_, _29200_);
  nor (_29202_, _29189_, _04596_);
  and (_29203_, _29202_, _29201_);
  nor (_29204_, _29203_, _29198_);
  nor (_29205_, _29204_, _03773_);
  nor (_29206_, _29129_, _04594_);
  and (_29207_, _29206_, _29201_);
  nor (_29208_, _29207_, _03653_);
  not (_29209_, _29208_);
  nor (_29211_, _29209_, _29205_);
  nor (_29212_, _13243_, _10824_);
  or (_29213_, _29124_, _04608_);
  nor (_29214_, _29213_, _29212_);
  or (_29215_, _29214_, _03786_);
  nor (_29216_, _29215_, _29211_);
  nor (_29217_, _13373_, _10824_);
  nor (_29218_, _29217_, _29124_);
  nor (_29219_, _29218_, _04606_);
  or (_29220_, _29219_, _29216_);
  and (_29222_, _29220_, _04260_);
  nor (_29223_, _29136_, _04260_);
  or (_29224_, _29223_, _29222_);
  and (_29225_, _29224_, _03206_);
  nor (_29226_, _29157_, _03206_);
  or (_29227_, _29226_, _29225_);
  and (_29228_, _29227_, _03820_);
  and (_29229_, _13425_, _05353_);
  nor (_29230_, _29229_, _29124_);
  nor (_29231_, _29230_, _03820_);
  or (_29233_, _29231_, _29228_);
  or (_29234_, _29233_, _43231_);
  or (_29235_, _43227_, \oc8051_golden_model_1.TCON [6]);
  and (_29236_, _29235_, _41991_);
  and (_43563_, _29236_, _29234_);
  not (_29237_, \oc8051_golden_model_1.TH0 [0]);
  nor (_29238_, _05304_, _29237_);
  nor (_29239_, _05744_, _10931_);
  nor (_29240_, _29239_, _29238_);
  and (_29241_, _29240_, _17220_);
  and (_29243_, _05304_, _04491_);
  nor (_29244_, _29243_, _29238_);
  and (_29245_, _29244_, _07441_);
  and (_29246_, _05304_, \oc8051_golden_model_1.ACC [0]);
  nor (_29247_, _29246_, _29238_);
  nor (_29248_, _29247_, _03611_);
  nor (_29249_, _29247_, _04500_);
  nor (_29250_, _04499_, _29237_);
  or (_29251_, _29250_, _29249_);
  and (_29252_, _29251_, _04515_);
  nor (_29254_, _29240_, _04515_);
  or (_29255_, _29254_, _29252_);
  and (_29256_, _29255_, _04524_);
  nor (_29257_, _29244_, _04524_);
  nor (_29258_, _29257_, _29256_);
  nor (_29259_, _29258_, _03603_);
  or (_29260_, _29259_, _07441_);
  nor (_29261_, _29260_, _29248_);
  nor (_29262_, _29261_, _29245_);
  nor (_29263_, _29262_, _05969_);
  and (_29265_, _06836_, _05304_);
  nor (_29266_, _29238_, _05970_);
  not (_29267_, _29266_);
  nor (_29268_, _29267_, _29265_);
  nor (_29269_, _29268_, _29263_);
  nor (_29270_, _29269_, _03644_);
  nor (_29271_, _12129_, _10931_);
  or (_29272_, _29238_, _03275_);
  nor (_29273_, _29272_, _29271_);
  or (_29274_, _29273_, _03650_);
  nor (_29276_, _29274_, _29270_);
  and (_29277_, _05304_, _06366_);
  nor (_29278_, _29277_, _29238_);
  nand (_29279_, _29278_, _04591_);
  and (_29280_, _29279_, _08861_);
  nor (_29281_, _29280_, _29276_);
  and (_29282_, _12019_, _05304_);
  nor (_29283_, _29282_, _29238_);
  and (_29284_, _29283_, _03649_);
  nor (_29285_, _29284_, _29281_);
  nor (_29287_, _29285_, _03778_);
  and (_29288_, _12145_, _05304_);
  or (_29289_, _29238_, _04589_);
  nor (_29290_, _29289_, _29288_);
  or (_29291_, _29290_, _03655_);
  nor (_29292_, _29291_, _29287_);
  or (_29293_, _29278_, _04596_);
  nor (_29294_, _29293_, _29239_);
  nor (_29295_, _29294_, _29292_);
  nor (_29296_, _29295_, _03773_);
  and (_29298_, _12144_, _05304_);
  or (_29299_, _29298_, _29238_);
  and (_29300_, _29299_, _03773_);
  or (_29301_, _29300_, _29296_);
  and (_29302_, _29301_, _04608_);
  nor (_29303_, _12017_, _10931_);
  nor (_29304_, _29303_, _29238_);
  nor (_29305_, _29304_, _04608_);
  or (_29306_, _29305_, _29302_);
  and (_29307_, _29306_, _04606_);
  nor (_29309_, _12015_, _10931_);
  nor (_29310_, _29309_, _29238_);
  nor (_29311_, _29310_, _04606_);
  nor (_29312_, _29311_, _17220_);
  not (_29313_, _29312_);
  nor (_29314_, _29313_, _29307_);
  nor (_29315_, _29314_, _29241_);
  or (_29316_, _29315_, _43231_);
  or (_29317_, _43227_, \oc8051_golden_model_1.TH0 [0]);
  and (_29318_, _29317_, _41991_);
  and (_43566_, _29318_, _29316_);
  and (_29320_, _06835_, _05304_);
  not (_29321_, \oc8051_golden_model_1.TH0 [1]);
  nor (_29322_, _05304_, _29321_);
  nor (_29323_, _29322_, _05970_);
  not (_29324_, _29323_);
  nor (_29325_, _29324_, _29320_);
  not (_29326_, _29325_);
  nor (_29327_, _05304_, \oc8051_golden_model_1.TH0 [1]);
  and (_29328_, _05304_, _03320_);
  nor (_29330_, _29328_, _29327_);
  and (_29331_, _29330_, _03603_);
  and (_29332_, _29330_, _04499_);
  nor (_29333_, _04499_, _29321_);
  or (_29334_, _29333_, _29332_);
  and (_29335_, _29334_, _04515_);
  and (_29336_, _12234_, _05304_);
  nor (_29337_, _29336_, _29327_);
  and (_29338_, _29337_, _03599_);
  or (_29339_, _29338_, _29335_);
  and (_29341_, _29339_, _04524_);
  and (_29342_, _05304_, _05898_);
  nor (_29343_, _29342_, _29322_);
  nor (_29344_, _29343_, _04524_);
  nor (_29345_, _29344_, _29341_);
  nor (_29346_, _29345_, _03603_);
  or (_29347_, _29346_, _07441_);
  nor (_29348_, _29347_, _29331_);
  and (_29349_, _29343_, _07441_);
  nor (_29350_, _29349_, _29348_);
  nor (_29352_, _29350_, _05969_);
  nor (_29353_, _29352_, _03644_);
  and (_29354_, _29353_, _29326_);
  not (_29355_, _29327_);
  and (_29356_, _12330_, _05304_);
  nor (_29357_, _29356_, _03275_);
  and (_29358_, _29357_, _29355_);
  nor (_29359_, _29358_, _29354_);
  nor (_29360_, _29359_, _08861_);
  nor (_29361_, _12220_, _10931_);
  nor (_29363_, _29361_, _04591_);
  and (_29364_, _05304_, _04347_);
  nor (_29365_, _29364_, _04582_);
  nor (_29366_, _29365_, _29363_);
  nor (_29367_, _29366_, _29327_);
  nor (_29368_, _29367_, _29360_);
  nor (_29369_, _29368_, _03778_);
  nor (_29370_, _12347_, _10931_);
  nor (_29371_, _29370_, _04589_);
  and (_29372_, _29371_, _29355_);
  nor (_29373_, _29372_, _29369_);
  nor (_29374_, _29373_, _03655_);
  nor (_29375_, _12219_, _10931_);
  nor (_29376_, _29375_, _04596_);
  and (_29377_, _29376_, _29355_);
  nor (_29378_, _29377_, _29374_);
  nor (_29379_, _29378_, _03773_);
  nor (_29380_, _29322_, _05699_);
  nor (_29381_, _29380_, _04594_);
  and (_29382_, _29381_, _29330_);
  nor (_29384_, _29382_, _29379_);
  or (_29385_, _29384_, _18553_);
  and (_29386_, _29364_, _05698_);
  nor (_29387_, _29386_, _04608_);
  and (_29388_, _29387_, _29355_);
  nand (_29389_, _29328_, _05698_);
  nor (_29390_, _29327_, _04606_);
  and (_29391_, _29390_, _29389_);
  or (_29392_, _29391_, _03809_);
  nor (_29393_, _29392_, _29388_);
  and (_29395_, _29393_, _29385_);
  nor (_29396_, _29337_, _04260_);
  nor (_29397_, _29396_, _29395_);
  and (_29398_, _29397_, _03820_);
  nor (_29399_, _29336_, _29322_);
  nor (_29400_, _29399_, _03820_);
  or (_29401_, _29400_, _29398_);
  or (_29402_, _29401_, _43231_);
  or (_29403_, _43227_, \oc8051_golden_model_1.TH0 [1]);
  and (_29404_, _29403_, _41991_);
  and (_43567_, _29404_, _29402_);
  not (_29406_, \oc8051_golden_model_1.TH0 [2]);
  nor (_29407_, _05304_, _29406_);
  nor (_29408_, _12543_, _10931_);
  nor (_29409_, _29408_, _29407_);
  nor (_29410_, _29409_, _04606_);
  and (_29411_, _06839_, _05304_);
  nor (_29412_, _29411_, _29407_);
  or (_29413_, _29412_, _05970_);
  and (_29414_, _05304_, \oc8051_golden_model_1.ACC [2]);
  nor (_29416_, _29414_, _29407_);
  nor (_29417_, _29416_, _03611_);
  nor (_29418_, _29416_, _04500_);
  nor (_29419_, _04499_, _29406_);
  or (_29420_, _29419_, _29418_);
  and (_29421_, _29420_, _04515_);
  nor (_29422_, _12430_, _10931_);
  nor (_29423_, _29422_, _29407_);
  nor (_29424_, _29423_, _04515_);
  or (_29425_, _29424_, _29421_);
  and (_29427_, _29425_, _04524_);
  nor (_29428_, _10931_, _05130_);
  nor (_29429_, _29428_, _29407_);
  nor (_29430_, _29429_, _04524_);
  nor (_29431_, _29430_, _29427_);
  nor (_29432_, _29431_, _03603_);
  or (_29433_, _29432_, _07441_);
  nor (_29434_, _29433_, _29417_);
  and (_29435_, _29429_, _07441_);
  or (_29436_, _29435_, _05969_);
  or (_29438_, _29436_, _29434_);
  and (_29439_, _29438_, _03275_);
  and (_29440_, _29439_, _29413_);
  nor (_29441_, _12524_, _10931_);
  or (_29442_, _29407_, _03275_);
  nor (_29443_, _29442_, _29441_);
  or (_29444_, _29443_, _03650_);
  nor (_29445_, _29444_, _29440_);
  and (_29446_, _05304_, _06414_);
  nor (_29447_, _29446_, _29407_);
  nand (_29449_, _29447_, _04591_);
  and (_29450_, _29449_, _08861_);
  nor (_29451_, _29450_, _29445_);
  and (_29452_, _12538_, _05304_);
  nor (_29453_, _29452_, _29407_);
  and (_29454_, _29453_, _03649_);
  nor (_29455_, _29454_, _29451_);
  nor (_29456_, _29455_, _03778_);
  and (_29457_, _12544_, _05304_);
  or (_29458_, _29407_, _04589_);
  nor (_29460_, _29458_, _29457_);
  or (_29461_, _29460_, _03655_);
  nor (_29462_, _29461_, _29456_);
  nor (_29463_, _29407_, _05793_);
  not (_29464_, _29463_);
  nor (_29465_, _29447_, _04596_);
  and (_29466_, _29465_, _29464_);
  nor (_29467_, _29466_, _29462_);
  nor (_29468_, _29467_, _03773_);
  nor (_29469_, _29416_, _04594_);
  and (_29471_, _29469_, _29464_);
  or (_29472_, _29471_, _29468_);
  and (_29473_, _29472_, _04608_);
  nor (_29474_, _12537_, _10931_);
  nor (_29475_, _29474_, _29407_);
  nor (_29476_, _29475_, _04608_);
  or (_29477_, _29476_, _29473_);
  and (_29478_, _29477_, _04606_);
  nor (_29479_, _29478_, _29410_);
  nor (_29480_, _29479_, _03809_);
  nor (_29482_, _29423_, _04260_);
  or (_29483_, _29482_, _03816_);
  nor (_29484_, _29483_, _29480_);
  and (_29485_, _12600_, _05304_);
  or (_29486_, _29407_, _03820_);
  nor (_29487_, _29486_, _29485_);
  nor (_29488_, _29487_, _29484_);
  or (_29489_, _29488_, _43231_);
  or (_29490_, _43227_, \oc8051_golden_model_1.TH0 [2]);
  and (_29491_, _29490_, _41991_);
  and (_43568_, _29491_, _29489_);
  not (_29492_, \oc8051_golden_model_1.TH0 [3]);
  nor (_29493_, _05304_, _29492_);
  nor (_29494_, _12618_, _10931_);
  nor (_29495_, _29494_, _29493_);
  nor (_29496_, _29495_, _04606_);
  and (_29497_, _05304_, \oc8051_golden_model_1.ACC [3]);
  nor (_29498_, _29497_, _29493_);
  nor (_29499_, _29498_, _04500_);
  nor (_29500_, _04499_, _29492_);
  or (_29503_, _29500_, _29499_);
  and (_29504_, _29503_, _04515_);
  nor (_29505_, _12625_, _10931_);
  nor (_29506_, _29505_, _29493_);
  nor (_29507_, _29506_, _04515_);
  or (_29508_, _29507_, _29504_);
  and (_29509_, _29508_, _04524_);
  nor (_29510_, _10931_, _04944_);
  nor (_29511_, _29510_, _29493_);
  nor (_29512_, _29511_, _04524_);
  nor (_29514_, _29512_, _29509_);
  nor (_29515_, _29514_, _03603_);
  nor (_29516_, _29498_, _03611_);
  nor (_29517_, _29516_, _07441_);
  not (_29518_, _29517_);
  nor (_29519_, _29518_, _29515_);
  and (_29520_, _29511_, _07441_);
  or (_29521_, _29520_, _05969_);
  or (_29522_, _29521_, _29519_);
  and (_29523_, _06838_, _05304_);
  nor (_29525_, _29523_, _29493_);
  or (_29526_, _29525_, _05970_);
  and (_29527_, _29526_, _03275_);
  and (_29528_, _29527_, _29522_);
  nor (_29529_, _12731_, _10931_);
  or (_29530_, _29493_, _03275_);
  nor (_29531_, _29530_, _29529_);
  or (_29532_, _29531_, _03650_);
  nor (_29533_, _29532_, _29528_);
  and (_29534_, _05304_, _06347_);
  nor (_29536_, _29534_, _29493_);
  nand (_29537_, _29536_, _04591_);
  and (_29538_, _29537_, _08861_);
  nor (_29539_, _29538_, _29533_);
  and (_29540_, _12746_, _05304_);
  nor (_29541_, _29540_, _29493_);
  and (_29542_, _29541_, _03649_);
  nor (_29543_, _29542_, _29539_);
  nor (_29544_, _29543_, _03778_);
  and (_29545_, _12619_, _05304_);
  or (_29547_, _29493_, _04589_);
  nor (_29548_, _29547_, _29545_);
  or (_29549_, _29548_, _03655_);
  nor (_29550_, _29549_, _29544_);
  nor (_29551_, _29493_, _05650_);
  not (_29552_, _29551_);
  nor (_29553_, _29536_, _04596_);
  and (_29554_, _29553_, _29552_);
  nor (_29555_, _29554_, _29550_);
  nor (_29556_, _29555_, _03773_);
  nor (_29558_, _29498_, _04594_);
  and (_29559_, _29558_, _29552_);
  nor (_29560_, _29559_, _03653_);
  not (_29561_, _29560_);
  nor (_29562_, _29561_, _29556_);
  nor (_29563_, _12745_, _10931_);
  or (_29564_, _29493_, _04608_);
  nor (_29565_, _29564_, _29563_);
  or (_29566_, _29565_, _03786_);
  nor (_29567_, _29566_, _29562_);
  nor (_29569_, _29567_, _29496_);
  nor (_29570_, _29569_, _03809_);
  nor (_29571_, _29506_, _04260_);
  or (_29572_, _29571_, _03816_);
  nor (_29573_, _29572_, _29570_);
  and (_29574_, _12806_, _05304_);
  or (_29575_, _29493_, _03820_);
  nor (_29576_, _29575_, _29574_);
  nor (_29577_, _29576_, _29573_);
  or (_29578_, _29577_, _43231_);
  or (_29580_, _43227_, \oc8051_golden_model_1.TH0 [3]);
  and (_29581_, _29580_, _41991_);
  and (_43569_, _29581_, _29578_);
  not (_29582_, \oc8051_golden_model_1.TH0 [4]);
  nor (_29583_, _05304_, _29582_);
  nor (_29584_, _12956_, _10931_);
  nor (_29585_, _29584_, _29583_);
  nor (_29586_, _29585_, _04606_);
  and (_29587_, _12957_, _05304_);
  nor (_29588_, _29587_, _29583_);
  nor (_29590_, _29588_, _04589_);
  and (_29591_, _06375_, _05304_);
  nor (_29592_, _29591_, _29583_);
  and (_29593_, _29592_, _03650_);
  and (_29594_, _05304_, \oc8051_golden_model_1.ACC [4]);
  nor (_29595_, _29594_, _29583_);
  nor (_29596_, _29595_, _03611_);
  nor (_29597_, _29595_, _04500_);
  nor (_29598_, _04499_, _29582_);
  or (_29599_, _29598_, _29597_);
  and (_29601_, _29599_, _04515_);
  nor (_29602_, _12820_, _10931_);
  nor (_29603_, _29602_, _29583_);
  nor (_29604_, _29603_, _04515_);
  or (_29605_, _29604_, _29601_);
  and (_29606_, _29605_, _04524_);
  nor (_29607_, _05840_, _10931_);
  nor (_29608_, _29607_, _29583_);
  nor (_29609_, _29608_, _04524_);
  nor (_29610_, _29609_, _29606_);
  nor (_29612_, _29610_, _03603_);
  or (_29613_, _29612_, _07441_);
  nor (_29614_, _29613_, _29596_);
  and (_29615_, _29608_, _07441_);
  nor (_29616_, _29615_, _29614_);
  nor (_29617_, _29616_, _05969_);
  and (_29618_, _06843_, _05304_);
  nor (_29619_, _29583_, _05970_);
  not (_29620_, _29619_);
  nor (_29621_, _29620_, _29618_);
  or (_29623_, _29621_, _03644_);
  nor (_29624_, _29623_, _29617_);
  nor (_29625_, _12936_, _10931_);
  nor (_29626_, _29625_, _29583_);
  nor (_29627_, _29626_, _03275_);
  or (_29628_, _29627_, _03650_);
  nor (_29629_, _29628_, _29624_);
  nor (_29630_, _29629_, _29593_);
  or (_29631_, _29630_, _03649_);
  and (_29632_, _12951_, _05304_);
  or (_29634_, _29632_, _29583_);
  or (_29635_, _29634_, _04591_);
  and (_29636_, _29635_, _04589_);
  and (_29637_, _29636_, _29631_);
  nor (_29638_, _29637_, _29590_);
  nor (_29639_, _29638_, _03655_);
  nor (_29640_, _29583_, _05889_);
  not (_29641_, _29640_);
  nor (_29642_, _29592_, _04596_);
  and (_29643_, _29642_, _29641_);
  nor (_29645_, _29643_, _29639_);
  nor (_29646_, _29645_, _03773_);
  nor (_29647_, _29595_, _04594_);
  and (_29648_, _29647_, _29641_);
  nor (_29649_, _29648_, _03653_);
  not (_29650_, _29649_);
  nor (_29651_, _29650_, _29646_);
  nor (_29652_, _12949_, _10931_);
  or (_29653_, _29583_, _04608_);
  nor (_29654_, _29653_, _29652_);
  or (_29656_, _29654_, _03786_);
  nor (_29657_, _29656_, _29651_);
  nor (_29658_, _29657_, _29586_);
  nor (_29659_, _29658_, _03809_);
  nor (_29660_, _29603_, _04260_);
  or (_29661_, _29660_, _03816_);
  nor (_29662_, _29661_, _29659_);
  and (_29663_, _13013_, _05304_);
  or (_29664_, _29583_, _03820_);
  nor (_29665_, _29664_, _29663_);
  nor (_29667_, _29665_, _29662_);
  or (_29668_, _29667_, _43231_);
  or (_29669_, _43227_, \oc8051_golden_model_1.TH0 [4]);
  and (_29670_, _29669_, _41991_);
  and (_43570_, _29670_, _29668_);
  not (_29671_, \oc8051_golden_model_1.TH0 [5]);
  nor (_29672_, _05304_, _29671_);
  nor (_29673_, _13159_, _10931_);
  nor (_29674_, _29673_, _29672_);
  nor (_29675_, _29674_, _04606_);
  and (_29677_, _13160_, _05304_);
  nor (_29678_, _29677_, _29672_);
  nor (_29679_, _29678_, _04589_);
  and (_29680_, _06842_, _05304_);
  or (_29681_, _29680_, _29672_);
  and (_29682_, _29681_, _05969_);
  and (_29683_, _05304_, \oc8051_golden_model_1.ACC [5]);
  nor (_29684_, _29683_, _29672_);
  nor (_29685_, _29684_, _04500_);
  nor (_29686_, _04499_, _29671_);
  or (_29688_, _29686_, _29685_);
  and (_29689_, _29688_, _04515_);
  nor (_29690_, _13035_, _10931_);
  nor (_29691_, _29690_, _29672_);
  nor (_29692_, _29691_, _04515_);
  or (_29693_, _29692_, _29689_);
  and (_29694_, _29693_, _04524_);
  nor (_29695_, _05552_, _10931_);
  nor (_29696_, _29695_, _29672_);
  nor (_29697_, _29696_, _04524_);
  nor (_29699_, _29697_, _29694_);
  nor (_29700_, _29699_, _03603_);
  nor (_29701_, _29684_, _03611_);
  nor (_29702_, _29701_, _07441_);
  not (_29703_, _29702_);
  nor (_29704_, _29703_, _29700_);
  and (_29705_, _29696_, _07441_);
  or (_29706_, _29705_, _05969_);
  nor (_29707_, _29706_, _29704_);
  or (_29708_, _29707_, _29682_);
  and (_29710_, _29708_, _03275_);
  nor (_29711_, _13139_, _10931_);
  nor (_29712_, _29711_, _29672_);
  nor (_29713_, _29712_, _03275_);
  or (_29714_, _29713_, _08861_);
  or (_29715_, _29714_, _29710_);
  and (_29716_, _13154_, _05304_);
  or (_29717_, _29672_, _04591_);
  or (_29718_, _29717_, _29716_);
  and (_29719_, _06358_, _05304_);
  nor (_29721_, _29719_, _29672_);
  and (_29722_, _29721_, _03650_);
  nor (_29723_, _29722_, _03778_);
  and (_29724_, _29723_, _29718_);
  and (_29725_, _29724_, _29715_);
  nor (_29726_, _29725_, _29679_);
  nor (_29727_, _29726_, _03655_);
  nor (_29728_, _29672_, _05601_);
  not (_29729_, _29728_);
  nor (_29730_, _29721_, _04596_);
  and (_29732_, _29730_, _29729_);
  nor (_29733_, _29732_, _29727_);
  nor (_29734_, _29733_, _03773_);
  nor (_29735_, _29684_, _04594_);
  and (_29736_, _29735_, _29729_);
  or (_29737_, _29736_, _29734_);
  and (_29738_, _29737_, _04608_);
  nor (_29739_, _13152_, _10931_);
  nor (_29740_, _29739_, _29672_);
  nor (_29741_, _29740_, _04608_);
  or (_29743_, _29741_, _29738_);
  and (_29744_, _29743_, _04606_);
  nor (_29745_, _29744_, _29675_);
  nor (_29746_, _29745_, _03809_);
  nor (_29747_, _29691_, _04260_);
  or (_29748_, _29747_, _03816_);
  nor (_29749_, _29748_, _29746_);
  and (_29750_, _13217_, _05304_);
  or (_29751_, _29672_, _03820_);
  nor (_29752_, _29751_, _29750_);
  nor (_29753_, _29752_, _29749_);
  or (_29754_, _29753_, _43231_);
  or (_29755_, _43227_, \oc8051_golden_model_1.TH0 [5]);
  and (_29756_, _29755_, _41991_);
  and (_43571_, _29756_, _29754_);
  not (_29757_, \oc8051_golden_model_1.TH0 [6]);
  nor (_29758_, _05304_, _29757_);
  nor (_29759_, _13373_, _10931_);
  nor (_29760_, _29759_, _29758_);
  nor (_29761_, _29760_, _04606_);
  and (_29764_, _13374_, _05304_);
  nor (_29765_, _29764_, _29758_);
  nor (_29766_, _29765_, _04589_);
  and (_29767_, _06531_, _05304_);
  or (_29768_, _29767_, _29758_);
  and (_29769_, _29768_, _05969_);
  and (_29770_, _05304_, \oc8051_golden_model_1.ACC [6]);
  nor (_29771_, _29770_, _29758_);
  nor (_29772_, _29771_, _03611_);
  nor (_29773_, _29771_, _04500_);
  nor (_29775_, _04499_, _29757_);
  or (_29776_, _29775_, _29773_);
  and (_29777_, _29776_, _04515_);
  nor (_29778_, _13235_, _10931_);
  nor (_29779_, _29778_, _29758_);
  nor (_29780_, _29779_, _04515_);
  or (_29781_, _29780_, _29777_);
  and (_29782_, _29781_, _04524_);
  nor (_29783_, _05442_, _10931_);
  nor (_29784_, _29783_, _29758_);
  nor (_29786_, _29784_, _04524_);
  nor (_29787_, _29786_, _29782_);
  nor (_29788_, _29787_, _03603_);
  or (_29789_, _29788_, _07441_);
  nor (_29790_, _29789_, _29772_);
  and (_29791_, _29784_, _07441_);
  or (_29792_, _29791_, _05969_);
  nor (_29793_, _29792_, _29790_);
  or (_29794_, _29793_, _29769_);
  and (_29795_, _29794_, _03275_);
  nor (_29797_, _13356_, _10931_);
  nor (_29798_, _29797_, _29758_);
  nor (_29799_, _29798_, _03275_);
  or (_29800_, _29799_, _08861_);
  or (_29801_, _29800_, _29795_);
  and (_29802_, _13245_, _05304_);
  or (_29803_, _29758_, _04591_);
  or (_29804_, _29803_, _29802_);
  and (_29805_, _13363_, _05304_);
  nor (_29806_, _29805_, _29758_);
  and (_29808_, _29806_, _03650_);
  nor (_29809_, _29808_, _03778_);
  and (_29810_, _29809_, _29804_);
  and (_29811_, _29810_, _29801_);
  nor (_29812_, _29811_, _29766_);
  nor (_29813_, _29812_, _03655_);
  nor (_29814_, _29758_, _05491_);
  not (_29815_, _29814_);
  nor (_29816_, _29806_, _04596_);
  and (_29817_, _29816_, _29815_);
  nor (_29819_, _29817_, _29813_);
  nor (_29820_, _29819_, _03773_);
  nor (_29821_, _29771_, _04594_);
  and (_29822_, _29821_, _29815_);
  nor (_29823_, _29822_, _03653_);
  not (_29824_, _29823_);
  nor (_29825_, _29824_, _29820_);
  nor (_29826_, _13243_, _10931_);
  or (_29827_, _29758_, _04608_);
  nor (_29828_, _29827_, _29826_);
  or (_29830_, _29828_, _03786_);
  nor (_29831_, _29830_, _29825_);
  nor (_29832_, _29831_, _29761_);
  nor (_29833_, _29832_, _03809_);
  nor (_29834_, _29779_, _04260_);
  or (_29835_, _29834_, _03816_);
  nor (_29836_, _29835_, _29833_);
  and (_29837_, _13425_, _05304_);
  or (_29838_, _29758_, _03820_);
  nor (_29839_, _29838_, _29837_);
  nor (_29841_, _29839_, _29836_);
  or (_29842_, _29841_, _43231_);
  or (_29843_, _43227_, \oc8051_golden_model_1.TH0 [6]);
  and (_29844_, _29843_, _41991_);
  and (_43572_, _29844_, _29842_);
  not (_29845_, \oc8051_golden_model_1.TH1 [0]);
  nor (_29846_, _05356_, _29845_);
  nor (_29847_, _05744_, _11013_);
  nor (_29848_, _29847_, _29846_);
  and (_29849_, _29848_, _17220_);
  and (_29851_, _05356_, \oc8051_golden_model_1.ACC [0]);
  nor (_29852_, _29851_, _29846_);
  nor (_29853_, _29852_, _03611_);
  nor (_29854_, _29853_, _07441_);
  nor (_29855_, _29848_, _04515_);
  nor (_29856_, _04499_, _29845_);
  nor (_29857_, _29852_, _04500_);
  nor (_29858_, _29857_, _29856_);
  nor (_29859_, _29858_, _03599_);
  or (_29860_, _29859_, _03597_);
  nor (_29862_, _29860_, _29855_);
  or (_29863_, _29862_, _03603_);
  and (_29864_, _29863_, _29854_);
  and (_29865_, _05356_, _04491_);
  or (_29866_, _29846_, _26194_);
  nor (_29867_, _29866_, _29865_);
  nor (_29868_, _29867_, _29864_);
  nor (_29869_, _29868_, _05969_);
  and (_29870_, _06836_, _05356_);
  nor (_29871_, _29846_, _05970_);
  not (_29873_, _29871_);
  nor (_29874_, _29873_, _29870_);
  nor (_29875_, _29874_, _29869_);
  nor (_29876_, _29875_, _03644_);
  nor (_29877_, _12129_, _11013_);
  or (_29878_, _29846_, _03275_);
  nor (_29879_, _29878_, _29877_);
  or (_29880_, _29879_, _03650_);
  nor (_29881_, _29880_, _29876_);
  and (_29882_, _05356_, _06366_);
  nor (_29884_, _29882_, _29846_);
  nand (_29885_, _29884_, _04591_);
  and (_29886_, _29885_, _08861_);
  nor (_29887_, _29886_, _29881_);
  and (_29888_, _12019_, _05356_);
  nor (_29889_, _29888_, _29846_);
  and (_29890_, _29889_, _03649_);
  nor (_29891_, _29890_, _29887_);
  nor (_29892_, _29891_, _03778_);
  and (_29893_, _12145_, _05356_);
  or (_29895_, _29846_, _04589_);
  nor (_29896_, _29895_, _29893_);
  or (_29897_, _29896_, _03655_);
  nor (_29898_, _29897_, _29892_);
  or (_29899_, _29884_, _04596_);
  nor (_29900_, _29899_, _29847_);
  nor (_29901_, _29900_, _29898_);
  nor (_29902_, _29901_, _03773_);
  nor (_29903_, _29846_, _05744_);
  or (_29904_, _29903_, _04594_);
  nor (_29906_, _29904_, _29852_);
  or (_29907_, _29906_, _29902_);
  and (_29908_, _29907_, _04608_);
  nor (_29909_, _12017_, _11013_);
  nor (_29910_, _29909_, _29846_);
  nor (_29911_, _29910_, _04608_);
  or (_29912_, _29911_, _29908_);
  and (_29913_, _29912_, _04606_);
  nor (_29914_, _12015_, _11013_);
  nor (_29915_, _29914_, _29846_);
  nor (_29917_, _29915_, _04606_);
  nor (_29918_, _29917_, _17220_);
  not (_29919_, _29918_);
  nor (_29920_, _29919_, _29913_);
  nor (_29921_, _29920_, _29849_);
  or (_29922_, _29921_, _43231_);
  or (_29923_, _43227_, \oc8051_golden_model_1.TH1 [0]);
  and (_29924_, _29923_, _41991_);
  and (_43574_, _29924_, _29922_);
  and (_29925_, _06835_, _05356_);
  not (_29927_, \oc8051_golden_model_1.TH1 [1]);
  nor (_29928_, _05356_, _29927_);
  nor (_29929_, _29928_, _05970_);
  not (_29930_, _29929_);
  nor (_29931_, _29930_, _29925_);
  not (_29932_, _29931_);
  and (_29933_, _05356_, _05898_);
  or (_29934_, _29928_, _26194_);
  nor (_29935_, _29934_, _29933_);
  nor (_29936_, _05356_, \oc8051_golden_model_1.TH1 [1]);
  and (_29938_, _05356_, _03320_);
  nor (_29939_, _29938_, _29936_);
  and (_29940_, _29939_, _03603_);
  nor (_29941_, _29940_, _07441_);
  and (_29942_, _12234_, _05356_);
  nor (_29943_, _29942_, _29936_);
  and (_29944_, _29943_, _03599_);
  and (_29945_, _29939_, _04499_);
  nor (_29946_, _04499_, _29927_);
  nor (_29947_, _29946_, _29945_);
  nor (_29949_, _29947_, _03599_);
  or (_29950_, _29949_, _03597_);
  nor (_29951_, _29950_, _29944_);
  or (_29952_, _29951_, _03603_);
  and (_29953_, _29952_, _29941_);
  nor (_29954_, _29953_, _29935_);
  nor (_29955_, _29954_, _05969_);
  nor (_29956_, _29955_, _03644_);
  and (_29957_, _29956_, _29932_);
  not (_29958_, _29936_);
  and (_29960_, _12330_, _05356_);
  nor (_29961_, _29960_, _03275_);
  and (_29962_, _29961_, _29958_);
  nor (_29963_, _29962_, _29957_);
  nor (_29964_, _29963_, _08861_);
  nor (_29965_, _12220_, _11013_);
  nor (_29966_, _29965_, _04591_);
  and (_29967_, _05356_, _04347_);
  nor (_29968_, _29967_, _04582_);
  nor (_29969_, _29968_, _29966_);
  nor (_29971_, _29969_, _29936_);
  nor (_29972_, _29971_, _29964_);
  nor (_29973_, _29972_, _03778_);
  nor (_29974_, _12347_, _11013_);
  nor (_29975_, _29974_, _04589_);
  and (_29976_, _29975_, _29958_);
  nor (_29977_, _29976_, _29973_);
  nor (_29978_, _29977_, _03655_);
  nor (_29979_, _12219_, _11013_);
  nor (_29980_, _29979_, _04596_);
  and (_29982_, _29980_, _29958_);
  nor (_29983_, _29982_, _29978_);
  nor (_29984_, _29983_, _03773_);
  nor (_29985_, _29928_, _05699_);
  nor (_29986_, _29985_, _04594_);
  and (_29987_, _29986_, _29939_);
  nor (_29988_, _29987_, _29984_);
  or (_29989_, _29988_, _18553_);
  nand (_29990_, _12346_, _05356_);
  and (_29991_, _29990_, _03786_);
  and (_29993_, _29991_, _29958_);
  nor (_29994_, _29993_, _03809_);
  and (_29995_, _29967_, _05698_);
  or (_29996_, _29936_, _04608_);
  or (_29997_, _29996_, _29995_);
  and (_29998_, _29997_, _29994_);
  and (_29999_, _29998_, _29989_);
  nor (_30000_, _29943_, _04260_);
  nor (_30001_, _30000_, _29999_);
  and (_30002_, _30001_, _03820_);
  nor (_30004_, _29942_, _29928_);
  nor (_30005_, _30004_, _03820_);
  or (_30006_, _30005_, _30002_);
  or (_30007_, _30006_, _43231_);
  or (_30008_, _43227_, \oc8051_golden_model_1.TH1 [1]);
  and (_30009_, _30008_, _41991_);
  and (_43575_, _30009_, _30007_);
  not (_30010_, \oc8051_golden_model_1.TH1 [2]);
  nor (_30011_, _05356_, _30010_);
  nor (_30012_, _12543_, _11013_);
  nor (_30014_, _30012_, _30011_);
  nor (_30015_, _30014_, _04606_);
  nor (_30016_, _11013_, _05130_);
  nor (_30017_, _30016_, _30011_);
  and (_30018_, _30017_, _07441_);
  nor (_30019_, _12430_, _11013_);
  nor (_30020_, _30019_, _30011_);
  nor (_30021_, _30020_, _04515_);
  nor (_30022_, _04499_, _30010_);
  and (_30023_, _05356_, \oc8051_golden_model_1.ACC [2]);
  nor (_30025_, _30023_, _30011_);
  nor (_30026_, _30025_, _04500_);
  nor (_30027_, _30026_, _30022_);
  nor (_30028_, _30027_, _03599_);
  or (_30029_, _30028_, _30021_);
  and (_30030_, _30029_, _04524_);
  nor (_30031_, _30017_, _04524_);
  or (_30032_, _30031_, _30030_);
  and (_30033_, _30032_, _03611_);
  nor (_30034_, _30025_, _03611_);
  nor (_30036_, _30034_, _07441_);
  not (_30037_, _30036_);
  nor (_30038_, _30037_, _30033_);
  nor (_30039_, _30038_, _30018_);
  nor (_30040_, _30039_, _05969_);
  and (_30041_, _06839_, _05356_);
  nor (_30042_, _30011_, _05970_);
  not (_30043_, _30042_);
  nor (_30044_, _30043_, _30041_);
  nor (_30045_, _30044_, _30040_);
  nor (_30047_, _30045_, _03644_);
  nor (_30048_, _12524_, _11013_);
  or (_30049_, _30011_, _03275_);
  nor (_30050_, _30049_, _30048_);
  or (_30051_, _30050_, _03650_);
  nor (_30052_, _30051_, _30047_);
  and (_30053_, _05356_, _06414_);
  nor (_30054_, _30053_, _30011_);
  nand (_30055_, _30054_, _04591_);
  and (_30056_, _30055_, _08861_);
  nor (_30057_, _30056_, _30052_);
  and (_30058_, _12538_, _05356_);
  nor (_30059_, _30058_, _30011_);
  and (_30060_, _30059_, _03649_);
  nor (_30061_, _30060_, _30057_);
  nor (_30062_, _30061_, _03778_);
  and (_30063_, _12544_, _05356_);
  or (_30064_, _30011_, _04589_);
  nor (_30065_, _30064_, _30063_);
  or (_30066_, _30065_, _03655_);
  nor (_30069_, _30066_, _30062_);
  nor (_30070_, _30011_, _05793_);
  not (_30071_, _30070_);
  nor (_30072_, _30054_, _04596_);
  and (_30073_, _30072_, _30071_);
  nor (_30074_, _30073_, _30069_);
  nor (_30075_, _30074_, _03773_);
  nor (_30076_, _30025_, _04594_);
  and (_30077_, _30076_, _30071_);
  or (_30078_, _30077_, _30075_);
  and (_30080_, _30078_, _04608_);
  nor (_30081_, _12537_, _11013_);
  nor (_30082_, _30081_, _30011_);
  nor (_30083_, _30082_, _04608_);
  or (_30084_, _30083_, _30080_);
  and (_30085_, _30084_, _04606_);
  nor (_30086_, _30085_, _30015_);
  nor (_30087_, _30086_, _03809_);
  nor (_30088_, _30020_, _04260_);
  or (_30089_, _30088_, _03816_);
  nor (_30090_, _30089_, _30087_);
  and (_30091_, _12600_, _05356_);
  or (_30092_, _30011_, _03820_);
  nor (_30093_, _30092_, _30091_);
  nor (_30094_, _30093_, _30090_);
  or (_30095_, _30094_, _43231_);
  or (_30096_, _43227_, \oc8051_golden_model_1.TH1 [2]);
  and (_30097_, _30096_, _41991_);
  and (_43576_, _30097_, _30095_);
  not (_30098_, \oc8051_golden_model_1.TH1 [3]);
  nor (_30100_, _05356_, _30098_);
  nor (_30101_, _12618_, _11013_);
  nor (_30102_, _30101_, _30100_);
  nor (_30103_, _30102_, _04606_);
  and (_30104_, _05356_, \oc8051_golden_model_1.ACC [3]);
  nor (_30105_, _30104_, _30100_);
  nor (_30106_, _30105_, _04500_);
  nor (_30107_, _04499_, _30098_);
  or (_30108_, _30107_, _30106_);
  and (_30109_, _30108_, _04515_);
  nor (_30111_, _12625_, _11013_);
  nor (_30112_, _30111_, _30100_);
  nor (_30113_, _30112_, _04515_);
  or (_30114_, _30113_, _30109_);
  and (_30115_, _30114_, _04524_);
  nor (_30116_, _11013_, _04944_);
  nor (_30117_, _30116_, _30100_);
  nor (_30118_, _30117_, _04524_);
  nor (_30119_, _30118_, _30115_);
  nor (_30120_, _30119_, _03603_);
  nor (_30122_, _30105_, _03611_);
  nor (_30123_, _30122_, _07441_);
  not (_30124_, _30123_);
  nor (_30125_, _30124_, _30120_);
  and (_30126_, _30117_, _07441_);
  or (_30127_, _30126_, _05969_);
  or (_30128_, _30127_, _30125_);
  and (_30129_, _06838_, _05356_);
  nor (_30130_, _30129_, _30100_);
  or (_30131_, _30130_, _05970_);
  and (_30133_, _30131_, _03275_);
  and (_30134_, _30133_, _30128_);
  nor (_30135_, _12731_, _11013_);
  or (_30136_, _30100_, _03275_);
  nor (_30137_, _30136_, _30135_);
  or (_30138_, _30137_, _03650_);
  nor (_30139_, _30138_, _30134_);
  and (_30140_, _05356_, _06347_);
  nor (_30141_, _30140_, _30100_);
  nand (_30142_, _30141_, _04591_);
  and (_30144_, _30142_, _08861_);
  nor (_30145_, _30144_, _30139_);
  and (_30146_, _12746_, _05356_);
  nor (_30147_, _30146_, _30100_);
  and (_30148_, _30147_, _03649_);
  nor (_30149_, _30148_, _30145_);
  nor (_30150_, _30149_, _03778_);
  and (_30151_, _12619_, _05356_);
  or (_30152_, _30100_, _04589_);
  nor (_30153_, _30152_, _30151_);
  or (_30155_, _30153_, _03655_);
  nor (_30156_, _30155_, _30150_);
  nor (_30157_, _30100_, _05650_);
  not (_30158_, _30157_);
  nor (_30159_, _30141_, _04596_);
  and (_30160_, _30159_, _30158_);
  nor (_30161_, _30160_, _30156_);
  nor (_30162_, _30161_, _03773_);
  nor (_30163_, _30105_, _04594_);
  and (_30164_, _30163_, _30158_);
  or (_30166_, _30164_, _30162_);
  and (_30167_, _30166_, _04608_);
  nor (_30168_, _12745_, _11013_);
  nor (_30169_, _30168_, _30100_);
  nor (_30170_, _30169_, _04608_);
  or (_30171_, _30170_, _30167_);
  and (_30172_, _30171_, _04606_);
  nor (_30173_, _30172_, _30103_);
  nor (_30174_, _30173_, _03809_);
  nor (_30175_, _30112_, _04260_);
  or (_30177_, _30175_, _03816_);
  nor (_30178_, _30177_, _30174_);
  and (_30179_, _12806_, _05356_);
  or (_30180_, _30100_, _03820_);
  nor (_30181_, _30180_, _30179_);
  nor (_30182_, _30181_, _30178_);
  or (_30183_, _30182_, _43231_);
  or (_30184_, _43227_, \oc8051_golden_model_1.TH1 [3]);
  and (_30185_, _30184_, _41991_);
  and (_43577_, _30185_, _30183_);
  not (_30187_, \oc8051_golden_model_1.TH1 [4]);
  nor (_30188_, _05356_, _30187_);
  nor (_30189_, _12956_, _11013_);
  nor (_30190_, _30189_, _30188_);
  nor (_30191_, _30190_, _04606_);
  and (_30192_, _12957_, _05356_);
  nor (_30193_, _30192_, _30188_);
  nor (_30194_, _30193_, _04589_);
  and (_30195_, _06375_, _05356_);
  nor (_30196_, _30195_, _30188_);
  and (_30198_, _30196_, _03650_);
  nor (_30199_, _05840_, _11013_);
  nor (_30200_, _30199_, _30188_);
  and (_30201_, _30200_, _07441_);
  and (_30202_, _05356_, \oc8051_golden_model_1.ACC [4]);
  nor (_30203_, _30202_, _30188_);
  nor (_30204_, _30203_, _04500_);
  nor (_30205_, _04499_, _30187_);
  or (_30206_, _30205_, _30204_);
  and (_30207_, _30206_, _04515_);
  nor (_30209_, _12820_, _11013_);
  nor (_30210_, _30209_, _30188_);
  nor (_30211_, _30210_, _04515_);
  or (_30212_, _30211_, _30207_);
  and (_30213_, _30212_, _04524_);
  nor (_30214_, _30200_, _04524_);
  nor (_30215_, _30214_, _30213_);
  nor (_30216_, _30215_, _03603_);
  nor (_30217_, _30203_, _03611_);
  nor (_30218_, _30217_, _07441_);
  not (_30220_, _30218_);
  nor (_30221_, _30220_, _30216_);
  nor (_30222_, _30221_, _30201_);
  nor (_30223_, _30222_, _05969_);
  and (_30224_, _06843_, _05356_);
  nor (_30225_, _30188_, _05970_);
  not (_30226_, _30225_);
  nor (_30227_, _30226_, _30224_);
  or (_30228_, _30227_, _03644_);
  nor (_30229_, _30228_, _30223_);
  nor (_30231_, _12936_, _11013_);
  nor (_30232_, _30231_, _30188_);
  nor (_30233_, _30232_, _03275_);
  or (_30234_, _30233_, _03650_);
  nor (_30235_, _30234_, _30229_);
  nor (_30236_, _30235_, _30198_);
  or (_30237_, _30236_, _03649_);
  and (_30238_, _12951_, _05356_);
  or (_30239_, _30238_, _30188_);
  or (_30240_, _30239_, _04591_);
  and (_30242_, _30240_, _04589_);
  and (_30243_, _30242_, _30237_);
  nor (_30244_, _30243_, _30194_);
  nor (_30245_, _30244_, _03655_);
  nor (_30246_, _30188_, _05889_);
  not (_30247_, _30246_);
  nor (_30248_, _30196_, _04596_);
  and (_30249_, _30248_, _30247_);
  nor (_30250_, _30249_, _30245_);
  nor (_30251_, _30250_, _03773_);
  nor (_30253_, _30203_, _04594_);
  and (_30254_, _30253_, _30247_);
  nor (_30255_, _30254_, _03653_);
  not (_30256_, _30255_);
  nor (_30257_, _30256_, _30251_);
  nor (_30258_, _12949_, _11013_);
  or (_30259_, _30188_, _04608_);
  nor (_30260_, _30259_, _30258_);
  or (_30261_, _30260_, _03786_);
  nor (_30262_, _30261_, _30257_);
  nor (_30264_, _30262_, _30191_);
  nor (_30265_, _30264_, _03809_);
  nor (_30266_, _30210_, _04260_);
  or (_30267_, _30266_, _03816_);
  nor (_30268_, _30267_, _30265_);
  and (_30269_, _13013_, _05356_);
  or (_30270_, _30188_, _03820_);
  nor (_30271_, _30270_, _30269_);
  nor (_30272_, _30271_, _30268_);
  or (_30273_, _30272_, _43231_);
  or (_30275_, _43227_, \oc8051_golden_model_1.TH1 [4]);
  and (_30276_, _30275_, _41991_);
  and (_43578_, _30276_, _30273_);
  not (_30277_, \oc8051_golden_model_1.TH1 [5]);
  nor (_30278_, _05356_, _30277_);
  nor (_30279_, _13159_, _11013_);
  nor (_30280_, _30279_, _30278_);
  nor (_30281_, _30280_, _04606_);
  and (_30282_, _13160_, _05356_);
  nor (_30283_, _30282_, _30278_);
  nor (_30285_, _30283_, _04589_);
  and (_30286_, _06842_, _05356_);
  or (_30287_, _30286_, _30278_);
  and (_30288_, _30287_, _05969_);
  and (_30289_, _05356_, \oc8051_golden_model_1.ACC [5]);
  nor (_30290_, _30289_, _30278_);
  nor (_30291_, _30290_, _04500_);
  nor (_30292_, _04499_, _30277_);
  or (_30293_, _30292_, _30291_);
  and (_30294_, _30293_, _04515_);
  nor (_30296_, _13035_, _11013_);
  nor (_30297_, _30296_, _30278_);
  nor (_30298_, _30297_, _04515_);
  or (_30299_, _30298_, _30294_);
  and (_30300_, _30299_, _04524_);
  nor (_30301_, _05552_, _11013_);
  nor (_30302_, _30301_, _30278_);
  nor (_30303_, _30302_, _04524_);
  nor (_30304_, _30303_, _30300_);
  nor (_30305_, _30304_, _03603_);
  nor (_30307_, _30290_, _03611_);
  nor (_30308_, _30307_, _07441_);
  not (_30309_, _30308_);
  nor (_30310_, _30309_, _30305_);
  and (_30311_, _30302_, _07441_);
  or (_30312_, _30311_, _05969_);
  nor (_30313_, _30312_, _30310_);
  or (_30314_, _30313_, _30288_);
  and (_30315_, _30314_, _03275_);
  nor (_30316_, _13139_, _11013_);
  nor (_30318_, _30316_, _30278_);
  nor (_30319_, _30318_, _03275_);
  or (_30320_, _30319_, _08861_);
  or (_30321_, _30320_, _30315_);
  and (_30322_, _13154_, _05356_);
  or (_30323_, _30278_, _04591_);
  or (_30324_, _30323_, _30322_);
  and (_30325_, _06358_, _05356_);
  nor (_30326_, _30325_, _30278_);
  and (_30327_, _30326_, _03650_);
  nor (_30329_, _30327_, _03778_);
  and (_30330_, _30329_, _30324_);
  and (_30331_, _30330_, _30321_);
  nor (_30332_, _30331_, _30285_);
  nor (_30333_, _30332_, _03655_);
  nor (_30334_, _30278_, _05601_);
  not (_30335_, _30334_);
  nor (_30336_, _30326_, _04596_);
  and (_30337_, _30336_, _30335_);
  nor (_30338_, _30337_, _30333_);
  nor (_30340_, _30338_, _03773_);
  nor (_30341_, _30290_, _04594_);
  and (_30342_, _30341_, _30335_);
  nor (_30343_, _30342_, _03653_);
  not (_30344_, _30343_);
  nor (_30345_, _30344_, _30340_);
  nor (_30346_, _13152_, _11013_);
  or (_30347_, _30278_, _04608_);
  nor (_30348_, _30347_, _30346_);
  or (_30349_, _30348_, _03786_);
  nor (_30351_, _30349_, _30345_);
  nor (_30352_, _30351_, _30281_);
  nor (_30353_, _30352_, _03809_);
  nor (_30354_, _30297_, _04260_);
  or (_30355_, _30354_, _03816_);
  nor (_30356_, _30355_, _30353_);
  and (_30357_, _13217_, _05356_);
  or (_30358_, _30278_, _03820_);
  nor (_30359_, _30358_, _30357_);
  nor (_30360_, _30359_, _30356_);
  or (_30362_, _30360_, _43231_);
  or (_30363_, _43227_, \oc8051_golden_model_1.TH1 [5]);
  and (_30364_, _30363_, _41991_);
  and (_43581_, _30364_, _30362_);
  not (_30365_, \oc8051_golden_model_1.TH1 [6]);
  nor (_30366_, _05356_, _30365_);
  nor (_30367_, _13373_, _11013_);
  nor (_30368_, _30367_, _30366_);
  nor (_30369_, _30368_, _04606_);
  and (_30370_, _13374_, _05356_);
  nor (_30372_, _30370_, _30366_);
  nor (_30373_, _30372_, _04589_);
  and (_30374_, _06531_, _05356_);
  or (_30375_, _30374_, _30366_);
  and (_30376_, _30375_, _05969_);
  and (_30377_, _05356_, \oc8051_golden_model_1.ACC [6]);
  nor (_30378_, _30377_, _30366_);
  nor (_30379_, _30378_, _04500_);
  nor (_30380_, _04499_, _30365_);
  or (_30381_, _30380_, _30379_);
  and (_30382_, _30381_, _04515_);
  nor (_30383_, _13235_, _11013_);
  nor (_30384_, _30383_, _30366_);
  nor (_30385_, _30384_, _04515_);
  or (_30386_, _30385_, _30382_);
  and (_30387_, _30386_, _04524_);
  nor (_30388_, _05442_, _11013_);
  nor (_30389_, _30388_, _30366_);
  nor (_30390_, _30389_, _04524_);
  nor (_30391_, _30390_, _30387_);
  nor (_30394_, _30391_, _03603_);
  nor (_30395_, _30378_, _03611_);
  nor (_30396_, _30395_, _07441_);
  not (_30397_, _30396_);
  nor (_30398_, _30397_, _30394_);
  and (_30399_, _30389_, _07441_);
  or (_30400_, _30399_, _05969_);
  nor (_30401_, _30400_, _30398_);
  or (_30402_, _30401_, _30376_);
  and (_30403_, _30402_, _03275_);
  nor (_30405_, _13356_, _11013_);
  nor (_30406_, _30405_, _30366_);
  nor (_30407_, _30406_, _03275_);
  or (_30408_, _30407_, _08861_);
  or (_30409_, _30408_, _30403_);
  and (_30410_, _13245_, _05356_);
  or (_30411_, _30366_, _04591_);
  or (_30412_, _30411_, _30410_);
  and (_30413_, _13363_, _05356_);
  nor (_30414_, _30413_, _30366_);
  and (_30416_, _30414_, _03650_);
  nor (_30417_, _30416_, _03778_);
  and (_30418_, _30417_, _30412_);
  and (_30419_, _30418_, _30409_);
  nor (_30420_, _30419_, _30373_);
  nor (_30421_, _30420_, _03655_);
  nor (_30422_, _30366_, _05491_);
  not (_30423_, _30422_);
  nor (_30424_, _30414_, _04596_);
  and (_30425_, _30424_, _30423_);
  nor (_30427_, _30425_, _30421_);
  nor (_30428_, _30427_, _03773_);
  nor (_30429_, _30378_, _04594_);
  and (_30430_, _30429_, _30423_);
  or (_30431_, _30430_, _30428_);
  and (_30432_, _30431_, _04608_);
  nor (_30433_, _13243_, _11013_);
  nor (_30434_, _30433_, _30366_);
  nor (_30435_, _30434_, _04608_);
  or (_30436_, _30435_, _30432_);
  and (_30438_, _30436_, _04606_);
  nor (_30439_, _30438_, _30369_);
  nor (_30440_, _30439_, _03809_);
  nor (_30441_, _30384_, _04260_);
  or (_30442_, _30441_, _03816_);
  nor (_30443_, _30442_, _30440_);
  and (_30444_, _13425_, _05356_);
  or (_30445_, _30366_, _03820_);
  nor (_30446_, _30445_, _30444_);
  nor (_30447_, _30446_, _30443_);
  or (_30449_, _30447_, _43231_);
  or (_30450_, _43227_, \oc8051_golden_model_1.TH1 [6]);
  and (_30451_, _30450_, _41991_);
  and (_43582_, _30451_, _30449_);
  not (_30452_, \oc8051_golden_model_1.TL0 [0]);
  nor (_30453_, _05350_, _30452_);
  nor (_30454_, _05744_, _11095_);
  nor (_30455_, _30454_, _30453_);
  and (_30456_, _30455_, _17220_);
  and (_30458_, _05350_, _04491_);
  nor (_30461_, _30458_, _30453_);
  and (_30463_, _30461_, _07441_);
  and (_30465_, _05350_, \oc8051_golden_model_1.ACC [0]);
  nor (_30467_, _30465_, _30453_);
  nor (_30469_, _30467_, _04500_);
  nor (_30471_, _04499_, _30452_);
  or (_30473_, _30471_, _30469_);
  and (_30475_, _30473_, _04515_);
  nor (_30477_, _30455_, _04515_);
  or (_30479_, _30477_, _30475_);
  and (_30481_, _30479_, _04524_);
  nor (_30482_, _30461_, _04524_);
  nor (_30483_, _30482_, _30481_);
  nor (_30484_, _30483_, _03603_);
  nor (_30485_, _30467_, _03611_);
  nor (_30486_, _30485_, _07441_);
  not (_30487_, _30486_);
  nor (_30488_, _30487_, _30484_);
  nor (_30489_, _30488_, _30463_);
  nor (_30490_, _30489_, _05969_);
  and (_30492_, _06836_, _05350_);
  nor (_30493_, _30453_, _05970_);
  not (_30494_, _30493_);
  nor (_30495_, _30494_, _30492_);
  nor (_30496_, _30495_, _30490_);
  nor (_30497_, _30496_, _03644_);
  nor (_30498_, _12129_, _11095_);
  or (_30499_, _30453_, _03275_);
  nor (_30500_, _30499_, _30498_);
  or (_30501_, _30500_, _03650_);
  nor (_30503_, _30501_, _30497_);
  and (_30504_, _05350_, _06366_);
  nor (_30505_, _30504_, _30453_);
  nor (_30506_, _30505_, _04582_);
  or (_30507_, _30506_, _30503_);
  and (_30508_, _30507_, _04591_);
  and (_30509_, _12019_, _05350_);
  nor (_30510_, _30509_, _30453_);
  nor (_30511_, _30510_, _04591_);
  or (_30512_, _30511_, _30508_);
  nor (_30514_, _30512_, _03778_);
  and (_30515_, _12145_, _05350_);
  or (_30516_, _30453_, _04589_);
  nor (_30517_, _30516_, _30515_);
  or (_30518_, _30517_, _03655_);
  nor (_30519_, _30518_, _30514_);
  or (_30520_, _30505_, _04596_);
  nor (_30521_, _30520_, _30454_);
  nor (_30522_, _30521_, _30519_);
  nor (_30523_, _30522_, _03773_);
  nor (_30525_, _30453_, _05744_);
  or (_30526_, _30525_, _04594_);
  nor (_30527_, _30526_, _30467_);
  or (_30528_, _30527_, _30523_);
  and (_30529_, _30528_, _04608_);
  nor (_30530_, _12017_, _11095_);
  nor (_30531_, _30530_, _30453_);
  nor (_30532_, _30531_, _04608_);
  or (_30533_, _30532_, _30529_);
  and (_30534_, _30533_, _04606_);
  nor (_30536_, _12015_, _11095_);
  nor (_30537_, _30536_, _30453_);
  nor (_30538_, _30537_, _04606_);
  nor (_30539_, _30538_, _17220_);
  not (_30540_, _30539_);
  nor (_30541_, _30540_, _30534_);
  nor (_30542_, _30541_, _30456_);
  or (_30543_, _30542_, _43231_);
  or (_30544_, _43227_, \oc8051_golden_model_1.TL0 [0]);
  and (_30545_, _30544_, _41991_);
  and (_43583_, _30545_, _30543_);
  and (_30547_, _06835_, _05350_);
  not (_30548_, \oc8051_golden_model_1.TL0 [1]);
  nor (_30549_, _05350_, _30548_);
  nor (_30550_, _30549_, _05970_);
  not (_30551_, _30550_);
  nor (_30552_, _30551_, _30547_);
  not (_30553_, _30552_);
  and (_30554_, _05350_, _05898_);
  nor (_30555_, _30554_, _30549_);
  and (_30557_, _30555_, _07441_);
  nor (_30558_, _05350_, \oc8051_golden_model_1.TL0 [1]);
  and (_30559_, _05350_, _03320_);
  nor (_30560_, _30559_, _30558_);
  and (_30561_, _30560_, _03603_);
  and (_30562_, _30560_, _04499_);
  nor (_30563_, _04499_, _30548_);
  or (_30564_, _30563_, _30562_);
  and (_30565_, _30564_, _04515_);
  and (_30566_, _12234_, _05350_);
  nor (_30568_, _30566_, _30558_);
  and (_30569_, _30568_, _03599_);
  or (_30570_, _30569_, _30565_);
  and (_30571_, _30570_, _04524_);
  nor (_30572_, _30555_, _04524_);
  nor (_30573_, _30572_, _30571_);
  nor (_30574_, _30573_, _03603_);
  or (_30575_, _30574_, _07441_);
  nor (_30576_, _30575_, _30561_);
  nor (_30577_, _30576_, _30557_);
  nor (_30579_, _30577_, _05969_);
  nor (_30580_, _30579_, _03644_);
  and (_30581_, _30580_, _30553_);
  not (_30582_, _30558_);
  and (_30583_, _12330_, _05350_);
  nor (_30584_, _30583_, _03275_);
  and (_30585_, _30584_, _30582_);
  nor (_30586_, _30585_, _30581_);
  nor (_30587_, _30586_, _08861_);
  nor (_30588_, _12220_, _11095_);
  nor (_30590_, _30588_, _04591_);
  and (_30591_, _05350_, _04347_);
  nor (_30592_, _30591_, _04582_);
  nor (_30593_, _30592_, _30590_);
  nor (_30594_, _30593_, _30558_);
  nor (_30595_, _30594_, _30587_);
  nor (_30596_, _30595_, _03778_);
  nor (_30597_, _12347_, _11095_);
  nor (_30598_, _30597_, _04589_);
  and (_30599_, _30598_, _30582_);
  nor (_30601_, _30599_, _30596_);
  nor (_30602_, _30601_, _03655_);
  nor (_30603_, _12219_, _11095_);
  nor (_30604_, _30603_, _04596_);
  and (_30605_, _30604_, _30582_);
  nor (_30606_, _30605_, _30602_);
  nor (_30607_, _30606_, _03773_);
  nor (_30608_, _30549_, _05699_);
  nor (_30609_, _30608_, _04594_);
  and (_30610_, _30609_, _30560_);
  nor (_30612_, _30610_, _30607_);
  or (_30613_, _30612_, _18553_);
  and (_30614_, _30559_, _05698_);
  nor (_30615_, _30614_, _04606_);
  and (_30616_, _30615_, _30582_);
  nor (_30617_, _30616_, _03809_);
  and (_30618_, _30591_, _05698_);
  or (_30619_, _30558_, _04608_);
  or (_30620_, _30619_, _30618_);
  and (_30621_, _30620_, _30617_);
  and (_30623_, _30621_, _30613_);
  nor (_30624_, _30568_, _04260_);
  nor (_30625_, _30624_, _30623_);
  and (_30626_, _30625_, _03820_);
  nor (_30627_, _30566_, _30549_);
  nor (_30628_, _30627_, _03820_);
  or (_30629_, _30628_, _30626_);
  or (_30630_, _30629_, _43231_);
  or (_30631_, _43227_, \oc8051_golden_model_1.TL0 [1]);
  and (_30632_, _30631_, _41991_);
  and (_43585_, _30632_, _30630_);
  not (_30634_, \oc8051_golden_model_1.TL0 [2]);
  nor (_30635_, _05350_, _30634_);
  nor (_30636_, _12543_, _11095_);
  nor (_30637_, _30636_, _30635_);
  nor (_30638_, _30637_, _04606_);
  and (_30639_, _06839_, _05350_);
  nor (_30640_, _30639_, _30635_);
  or (_30641_, _30640_, _05970_);
  and (_30642_, _05350_, \oc8051_golden_model_1.ACC [2]);
  nor (_30644_, _30642_, _30635_);
  nor (_30645_, _30644_, _03611_);
  nor (_30646_, _30644_, _04500_);
  nor (_30647_, _04499_, _30634_);
  or (_30648_, _30647_, _30646_);
  and (_30649_, _30648_, _04515_);
  nor (_30650_, _12430_, _11095_);
  nor (_30651_, _30650_, _30635_);
  nor (_30652_, _30651_, _04515_);
  or (_30653_, _30652_, _30649_);
  and (_30655_, _30653_, _04524_);
  nor (_30656_, _11095_, _05130_);
  nor (_30657_, _30656_, _30635_);
  nor (_30658_, _30657_, _04524_);
  nor (_30659_, _30658_, _30655_);
  nor (_30660_, _30659_, _03603_);
  or (_30661_, _30660_, _07441_);
  nor (_30662_, _30661_, _30645_);
  and (_30663_, _30657_, _07441_);
  or (_30664_, _30663_, _05969_);
  or (_30666_, _30664_, _30662_);
  and (_30667_, _30666_, _03275_);
  and (_30668_, _30667_, _30641_);
  nor (_30669_, _12524_, _11095_);
  or (_30670_, _30635_, _03275_);
  nor (_30671_, _30670_, _30669_);
  or (_30672_, _30671_, _03650_);
  nor (_30673_, _30672_, _30668_);
  and (_30674_, _05350_, _06414_);
  nor (_30675_, _30674_, _30635_);
  nor (_30677_, _30675_, _04582_);
  or (_30678_, _30677_, _30673_);
  and (_30679_, _30678_, _04591_);
  and (_30680_, _12538_, _05350_);
  nor (_30681_, _30680_, _30635_);
  nor (_30682_, _30681_, _04591_);
  or (_30683_, _30682_, _30679_);
  nor (_30684_, _30683_, _03778_);
  and (_30685_, _12544_, _05350_);
  or (_30686_, _30635_, _04589_);
  nor (_30688_, _30686_, _30685_);
  or (_30689_, _30688_, _03655_);
  nor (_30690_, _30689_, _30684_);
  nor (_30691_, _30635_, _05793_);
  not (_30692_, _30691_);
  nor (_30693_, _30675_, _04596_);
  and (_30694_, _30693_, _30692_);
  nor (_30695_, _30694_, _30690_);
  nor (_30696_, _30695_, _03773_);
  nor (_30697_, _30644_, _04594_);
  and (_30699_, _30697_, _30692_);
  nor (_30700_, _30699_, _03653_);
  not (_30701_, _30700_);
  nor (_30702_, _30701_, _30696_);
  nor (_30703_, _12537_, _11095_);
  or (_30704_, _30635_, _04608_);
  nor (_30705_, _30704_, _30703_);
  or (_30706_, _30705_, _03786_);
  nor (_30707_, _30706_, _30702_);
  nor (_30708_, _30707_, _30638_);
  nor (_30710_, _30708_, _03809_);
  nor (_30711_, _30651_, _04260_);
  or (_30712_, _30711_, _03816_);
  nor (_30713_, _30712_, _30710_);
  and (_30714_, _12600_, _05350_);
  or (_30715_, _30635_, _03820_);
  nor (_30716_, _30715_, _30714_);
  nor (_30717_, _30716_, _30713_);
  or (_30718_, _30717_, _43231_);
  or (_30719_, _43227_, \oc8051_golden_model_1.TL0 [2]);
  and (_30721_, _30719_, _41991_);
  and (_43586_, _30721_, _30718_);
  not (_30722_, \oc8051_golden_model_1.TL0 [3]);
  nor (_30723_, _05350_, _30722_);
  nor (_30724_, _12618_, _11095_);
  nor (_30725_, _30724_, _30723_);
  nor (_30726_, _30725_, _04606_);
  and (_30727_, _12619_, _05350_);
  nor (_30728_, _30727_, _30723_);
  nor (_30729_, _30728_, _04589_);
  and (_30731_, _06838_, _05350_);
  or (_30732_, _30731_, _30723_);
  and (_30733_, _30732_, _05969_);
  and (_30734_, _05350_, \oc8051_golden_model_1.ACC [3]);
  nor (_30735_, _30734_, _30723_);
  nor (_30736_, _30735_, _03611_);
  nor (_30737_, _30735_, _04500_);
  nor (_30738_, _04499_, _30722_);
  or (_30739_, _30738_, _30737_);
  and (_30740_, _30739_, _04515_);
  nor (_30742_, _12625_, _11095_);
  nor (_30743_, _30742_, _30723_);
  nor (_30744_, _30743_, _04515_);
  or (_30745_, _30744_, _30740_);
  and (_30746_, _30745_, _04524_);
  nor (_30747_, _11095_, _04944_);
  nor (_30748_, _30747_, _30723_);
  nor (_30749_, _30748_, _04524_);
  nor (_30750_, _30749_, _30746_);
  nor (_30751_, _30750_, _03603_);
  or (_30753_, _30751_, _07441_);
  nor (_30754_, _30753_, _30736_);
  and (_30755_, _30748_, _07441_);
  or (_30756_, _30755_, _05969_);
  nor (_30757_, _30756_, _30754_);
  or (_30758_, _30757_, _30733_);
  and (_30759_, _30758_, _03275_);
  nor (_30760_, _12731_, _11095_);
  nor (_30761_, _30760_, _30723_);
  nor (_30762_, _30761_, _03275_);
  or (_30764_, _30762_, _08861_);
  or (_30765_, _30764_, _30759_);
  and (_30766_, _12746_, _05350_);
  or (_30767_, _30723_, _04591_);
  or (_30768_, _30767_, _30766_);
  and (_30769_, _05350_, _06347_);
  nor (_30770_, _30769_, _30723_);
  and (_30771_, _30770_, _03650_);
  nor (_30772_, _30771_, _03778_);
  and (_30773_, _30772_, _30768_);
  and (_30775_, _30773_, _30765_);
  nor (_30776_, _30775_, _30729_);
  nor (_30777_, _30776_, _03655_);
  nor (_30778_, _30723_, _05650_);
  not (_30779_, _30778_);
  nor (_30780_, _30770_, _04596_);
  and (_30781_, _30780_, _30779_);
  nor (_30782_, _30781_, _30777_);
  nor (_30783_, _30782_, _03773_);
  nor (_30784_, _30735_, _04594_);
  and (_30786_, _30784_, _30779_);
  or (_30787_, _30786_, _30783_);
  and (_30788_, _30787_, _04608_);
  nor (_30789_, _12745_, _11095_);
  nor (_30790_, _30789_, _30723_);
  nor (_30791_, _30790_, _04608_);
  or (_30792_, _30791_, _30788_);
  and (_30793_, _30792_, _04606_);
  nor (_30794_, _30793_, _30726_);
  nor (_30795_, _30794_, _03809_);
  nor (_30797_, _30743_, _04260_);
  or (_30798_, _30797_, _03816_);
  nor (_30799_, _30798_, _30795_);
  and (_30800_, _12806_, _05350_);
  or (_30801_, _30723_, _03820_);
  nor (_30802_, _30801_, _30800_);
  nor (_30803_, _30802_, _30799_);
  or (_30804_, _30803_, _43231_);
  or (_30805_, _43227_, \oc8051_golden_model_1.TL0 [3]);
  and (_30806_, _30805_, _41991_);
  and (_43587_, _30806_, _30804_);
  not (_30808_, \oc8051_golden_model_1.TL0 [4]);
  nor (_30809_, _05350_, _30808_);
  nor (_30810_, _12956_, _11095_);
  nor (_30811_, _30810_, _30809_);
  nor (_30812_, _30811_, _04606_);
  and (_30813_, _12957_, _05350_);
  nor (_30814_, _30813_, _30809_);
  nor (_30815_, _30814_, _04589_);
  and (_30816_, _06375_, _05350_);
  nor (_30818_, _30816_, _30809_);
  and (_30819_, _30818_, _03650_);
  nor (_30820_, _05840_, _11095_);
  nor (_30821_, _30820_, _30809_);
  and (_30822_, _30821_, _07441_);
  and (_30823_, _05350_, \oc8051_golden_model_1.ACC [4]);
  nor (_30824_, _30823_, _30809_);
  nor (_30825_, _30824_, _03611_);
  nor (_30826_, _30824_, _04500_);
  nor (_30827_, _04499_, _30808_);
  or (_30828_, _30827_, _30826_);
  and (_30829_, _30828_, _04515_);
  nor (_30830_, _12820_, _11095_);
  nor (_30831_, _30830_, _30809_);
  nor (_30832_, _30831_, _04515_);
  or (_30833_, _30832_, _30829_);
  and (_30834_, _30833_, _04524_);
  nor (_30835_, _30821_, _04524_);
  nor (_30836_, _30835_, _30834_);
  nor (_30837_, _30836_, _03603_);
  or (_30839_, _30837_, _07441_);
  nor (_30840_, _30839_, _30825_);
  nor (_30841_, _30840_, _30822_);
  nor (_30842_, _30841_, _05969_);
  and (_30843_, _06843_, _05350_);
  nor (_30844_, _30809_, _05970_);
  not (_30845_, _30844_);
  nor (_30846_, _30845_, _30843_);
  or (_30847_, _30846_, _03644_);
  nor (_30848_, _30847_, _30842_);
  nor (_30850_, _12936_, _11095_);
  nor (_30851_, _30850_, _30809_);
  nor (_30852_, _30851_, _03275_);
  or (_30853_, _30852_, _03650_);
  nor (_30854_, _30853_, _30848_);
  nor (_30855_, _30854_, _30819_);
  or (_30856_, _30855_, _03649_);
  and (_30857_, _12951_, _05350_);
  or (_30858_, _30857_, _30809_);
  or (_30859_, _30858_, _04591_);
  and (_30861_, _30859_, _04589_);
  and (_30862_, _30861_, _30856_);
  nor (_30863_, _30862_, _30815_);
  nor (_30864_, _30863_, _03655_);
  nor (_30865_, _30809_, _05889_);
  not (_30866_, _30865_);
  nor (_30867_, _30818_, _04596_);
  and (_30868_, _30867_, _30866_);
  nor (_30869_, _30868_, _30864_);
  nor (_30870_, _30869_, _03773_);
  nor (_30871_, _30824_, _04594_);
  and (_30872_, _30871_, _30866_);
  or (_30873_, _30872_, _30870_);
  and (_30874_, _30873_, _04608_);
  nor (_30875_, _12949_, _11095_);
  nor (_30876_, _30875_, _30809_);
  nor (_30877_, _30876_, _04608_);
  or (_30878_, _30877_, _30874_);
  and (_30879_, _30878_, _04606_);
  nor (_30880_, _30879_, _30812_);
  nor (_30883_, _30880_, _03809_);
  nor (_30884_, _30831_, _04260_);
  or (_30885_, _30884_, _03816_);
  nor (_30886_, _30885_, _30883_);
  and (_30887_, _13013_, _05350_);
  or (_30888_, _30809_, _03820_);
  nor (_30889_, _30888_, _30887_);
  nor (_30890_, _30889_, _30886_);
  or (_30891_, _30890_, _43231_);
  or (_30892_, _43227_, \oc8051_golden_model_1.TL0 [4]);
  and (_30894_, _30892_, _41991_);
  and (_43588_, _30894_, _30891_);
  not (_30895_, \oc8051_golden_model_1.TL0 [5]);
  nor (_30896_, _05350_, _30895_);
  nor (_30897_, _13159_, _11095_);
  nor (_30898_, _30897_, _30896_);
  nor (_30899_, _30898_, _04606_);
  and (_30900_, _13160_, _05350_);
  nor (_30901_, _30900_, _30896_);
  nor (_30902_, _30901_, _04589_);
  and (_30904_, _06842_, _05350_);
  or (_30905_, _30904_, _30896_);
  and (_30906_, _30905_, _05969_);
  and (_30907_, _05350_, \oc8051_golden_model_1.ACC [5]);
  nor (_30908_, _30907_, _30896_);
  nor (_30909_, _30908_, _03611_);
  nor (_30910_, _30908_, _04500_);
  nor (_30911_, _04499_, _30895_);
  or (_30912_, _30911_, _30910_);
  and (_30913_, _30912_, _04515_);
  nor (_30915_, _13035_, _11095_);
  nor (_30916_, _30915_, _30896_);
  nor (_30917_, _30916_, _04515_);
  or (_30918_, _30917_, _30913_);
  and (_30919_, _30918_, _04524_);
  nor (_30920_, _05552_, _11095_);
  nor (_30921_, _30920_, _30896_);
  nor (_30922_, _30921_, _04524_);
  nor (_30923_, _30922_, _30919_);
  nor (_30924_, _30923_, _03603_);
  or (_30926_, _30924_, _07441_);
  nor (_30927_, _30926_, _30909_);
  and (_30928_, _30921_, _07441_);
  or (_30929_, _30928_, _05969_);
  nor (_30930_, _30929_, _30927_);
  or (_30931_, _30930_, _30906_);
  and (_30932_, _30931_, _03275_);
  nor (_30933_, _13139_, _11095_);
  nor (_30934_, _30933_, _30896_);
  nor (_30935_, _30934_, _03275_);
  or (_30937_, _30935_, _08861_);
  or (_30938_, _30937_, _30932_);
  and (_30939_, _13154_, _05350_);
  or (_30940_, _30896_, _04591_);
  or (_30941_, _30940_, _30939_);
  and (_30942_, _06358_, _05350_);
  nor (_30943_, _30942_, _30896_);
  and (_30944_, _30943_, _03650_);
  nor (_30945_, _30944_, _03778_);
  and (_30946_, _30945_, _30941_);
  and (_30948_, _30946_, _30938_);
  nor (_30949_, _30948_, _30902_);
  nor (_30950_, _30949_, _03655_);
  nor (_30951_, _30896_, _05601_);
  not (_30952_, _30951_);
  nor (_30953_, _30943_, _04596_);
  and (_30954_, _30953_, _30952_);
  nor (_30955_, _30954_, _30950_);
  nor (_30956_, _30955_, _03773_);
  nor (_30957_, _30908_, _04594_);
  and (_30959_, _30957_, _30952_);
  nor (_30960_, _30959_, _03653_);
  not (_30961_, _30960_);
  nor (_30962_, _30961_, _30956_);
  nor (_30963_, _13152_, _11095_);
  or (_30964_, _30896_, _04608_);
  nor (_30965_, _30964_, _30963_);
  or (_30966_, _30965_, _03786_);
  nor (_30967_, _30966_, _30962_);
  nor (_30968_, _30967_, _30899_);
  nor (_30970_, _30968_, _03809_);
  nor (_30971_, _30916_, _04260_);
  or (_30972_, _30971_, _03816_);
  nor (_30973_, _30972_, _30970_);
  and (_30974_, _13217_, _05350_);
  or (_30975_, _30896_, _03820_);
  nor (_30976_, _30975_, _30974_);
  nor (_30977_, _30976_, _30973_);
  or (_30978_, _30977_, _43231_);
  or (_30979_, _43227_, \oc8051_golden_model_1.TL0 [5]);
  and (_30981_, _30979_, _41991_);
  and (_43589_, _30981_, _30978_);
  not (_30982_, \oc8051_golden_model_1.TL0 [6]);
  nor (_30983_, _05350_, _30982_);
  nor (_30984_, _13373_, _11095_);
  nor (_30985_, _30984_, _30983_);
  nor (_30986_, _30985_, _04606_);
  and (_30987_, _13374_, _05350_);
  nor (_30988_, _30987_, _30983_);
  nor (_30989_, _30988_, _04589_);
  and (_30991_, _06531_, _05350_);
  or (_30992_, _30991_, _30983_);
  and (_30993_, _30992_, _05969_);
  and (_30994_, _05350_, \oc8051_golden_model_1.ACC [6]);
  nor (_30995_, _30994_, _30983_);
  nor (_30996_, _30995_, _03611_);
  nor (_30997_, _30995_, _04500_);
  nor (_30998_, _04499_, _30982_);
  or (_30999_, _30998_, _30997_);
  and (_31000_, _30999_, _04515_);
  nor (_31002_, _13235_, _11095_);
  nor (_31003_, _31002_, _30983_);
  nor (_31004_, _31003_, _04515_);
  or (_31005_, _31004_, _31000_);
  and (_31006_, _31005_, _04524_);
  nor (_31007_, _05442_, _11095_);
  nor (_31008_, _31007_, _30983_);
  nor (_31009_, _31008_, _04524_);
  nor (_31010_, _31009_, _31006_);
  nor (_31011_, _31010_, _03603_);
  or (_31013_, _31011_, _07441_);
  nor (_31014_, _31013_, _30996_);
  and (_31015_, _31008_, _07441_);
  or (_31016_, _31015_, _05969_);
  nor (_31017_, _31016_, _31014_);
  or (_31018_, _31017_, _30993_);
  and (_31019_, _31018_, _03275_);
  nor (_31020_, _13356_, _11095_);
  nor (_31021_, _31020_, _30983_);
  nor (_31022_, _31021_, _03275_);
  or (_31024_, _31022_, _08861_);
  or (_31025_, _31024_, _31019_);
  and (_31026_, _13245_, _05350_);
  or (_31027_, _30983_, _04591_);
  or (_31028_, _31027_, _31026_);
  and (_31029_, _13363_, _05350_);
  nor (_31030_, _31029_, _30983_);
  and (_31031_, _31030_, _03650_);
  nor (_31032_, _31031_, _03778_);
  and (_31033_, _31032_, _31028_);
  and (_31035_, _31033_, _31025_);
  nor (_31036_, _31035_, _30989_);
  nor (_31037_, _31036_, _03655_);
  nor (_31038_, _30983_, _05491_);
  not (_31039_, _31038_);
  nor (_31040_, _31030_, _04596_);
  and (_31041_, _31040_, _31039_);
  nor (_31042_, _31041_, _31037_);
  nor (_31043_, _31042_, _03773_);
  nor (_31044_, _30995_, _04594_);
  and (_31046_, _31044_, _31039_);
  nor (_31047_, _31046_, _03653_);
  not (_31048_, _31047_);
  nor (_31049_, _31048_, _31043_);
  nor (_31050_, _13243_, _11095_);
  or (_31051_, _30983_, _04608_);
  nor (_31052_, _31051_, _31050_);
  or (_31053_, _31052_, _03786_);
  nor (_31054_, _31053_, _31049_);
  nor (_31055_, _31054_, _30986_);
  nor (_31057_, _31055_, _03809_);
  nor (_31058_, _31003_, _04260_);
  or (_31059_, _31058_, _03816_);
  nor (_31060_, _31059_, _31057_);
  and (_31061_, _13425_, _05350_);
  or (_31062_, _30983_, _03820_);
  nor (_31063_, _31062_, _31061_);
  nor (_31064_, _31063_, _31060_);
  or (_31065_, _31064_, _43231_);
  or (_31066_, _43227_, \oc8051_golden_model_1.TL0 [6]);
  and (_31068_, _31066_, _41991_);
  and (_43590_, _31068_, _31065_);
  not (_31069_, \oc8051_golden_model_1.TL1 [0]);
  nor (_31070_, _05309_, _31069_);
  nor (_31071_, _05744_, _11178_);
  nor (_31072_, _31071_, _31070_);
  and (_31073_, _31072_, _17220_);
  and (_31074_, _05309_, _04491_);
  nor (_31075_, _31074_, _31070_);
  and (_31076_, _31075_, _07441_);
  and (_31078_, _05309_, \oc8051_golden_model_1.ACC [0]);
  nor (_31079_, _31078_, _31070_);
  nor (_31080_, _31079_, _03611_);
  nor (_31081_, _31079_, _04500_);
  nor (_31082_, _04499_, _31069_);
  or (_31083_, _31082_, _31081_);
  and (_31084_, _31083_, _04515_);
  nor (_31085_, _31072_, _04515_);
  or (_31086_, _31085_, _31084_);
  and (_31087_, _31086_, _04524_);
  nor (_31089_, _31075_, _04524_);
  nor (_31090_, _31089_, _31087_);
  nor (_31091_, _31090_, _03603_);
  or (_31092_, _31091_, _07441_);
  nor (_31093_, _31092_, _31080_);
  nor (_31094_, _31093_, _31076_);
  nor (_31095_, _31094_, _05969_);
  and (_31096_, _06836_, _05309_);
  nor (_31097_, _31070_, _05970_);
  not (_31098_, _31097_);
  nor (_31099_, _31098_, _31096_);
  nor (_31100_, _31099_, _31095_);
  nor (_31101_, _31100_, _03644_);
  nor (_31102_, _12129_, _11178_);
  or (_31103_, _31070_, _03275_);
  nor (_31104_, _31103_, _31102_);
  or (_31105_, _31104_, _03650_);
  nor (_31106_, _31105_, _31101_);
  and (_31107_, _05309_, _06366_);
  nor (_31108_, _31107_, _31070_);
  nor (_31111_, _31108_, _04582_);
  or (_31112_, _31111_, _31106_);
  and (_31113_, _31112_, _04591_);
  and (_31114_, _12019_, _05309_);
  nor (_31115_, _31114_, _31070_);
  nor (_31116_, _31115_, _04591_);
  or (_31117_, _31116_, _31113_);
  nor (_31118_, _31117_, _03778_);
  and (_31119_, _12145_, _05309_);
  or (_31120_, _31070_, _04589_);
  nor (_31122_, _31120_, _31119_);
  or (_31123_, _31122_, _03655_);
  nor (_31124_, _31123_, _31118_);
  or (_31125_, _31108_, _04596_);
  nor (_31126_, _31125_, _31071_);
  nor (_31127_, _31126_, _31124_);
  nor (_31128_, _31127_, _03773_);
  nor (_31129_, _31070_, _05744_);
  or (_31130_, _31129_, _04594_);
  nor (_31131_, _31130_, _31079_);
  or (_31133_, _31131_, _31128_);
  and (_31134_, _31133_, _04608_);
  nor (_31135_, _12017_, _11178_);
  nor (_31136_, _31135_, _31070_);
  nor (_31137_, _31136_, _04608_);
  or (_31138_, _31137_, _31134_);
  and (_31139_, _31138_, _04606_);
  nor (_31140_, _12015_, _11178_);
  nor (_31141_, _31140_, _31070_);
  nor (_31142_, _31141_, _04606_);
  nor (_31144_, _31142_, _17220_);
  not (_31145_, _31144_);
  nor (_31146_, _31145_, _31139_);
  nor (_31147_, _31146_, _31073_);
  or (_31148_, _31147_, _43231_);
  or (_31149_, _43227_, \oc8051_golden_model_1.TL1 [0]);
  and (_31150_, _31149_, _41991_);
  and (_43592_, _31150_, _31148_);
  and (_31151_, _06835_, _05309_);
  not (_31152_, \oc8051_golden_model_1.TL1 [1]);
  nor (_31154_, _05309_, _31152_);
  nor (_31155_, _31154_, _05970_);
  not (_31156_, _31155_);
  nor (_31157_, _31156_, _31151_);
  not (_31158_, _31157_);
  nor (_31159_, _05309_, \oc8051_golden_model_1.TL1 [1]);
  and (_31160_, _05309_, _03320_);
  nor (_31161_, _31160_, _31159_);
  and (_31162_, _31161_, _03603_);
  and (_31163_, _31161_, _04499_);
  nor (_31165_, _04499_, _31152_);
  or (_31166_, _31165_, _31163_);
  and (_31167_, _31166_, _04515_);
  and (_31168_, _12234_, _05309_);
  nor (_31169_, _31168_, _31159_);
  and (_31170_, _31169_, _03599_);
  or (_31171_, _31170_, _31167_);
  and (_31172_, _31171_, _04524_);
  and (_31173_, _05309_, _05898_);
  nor (_31174_, _31173_, _31154_);
  nor (_31176_, _31174_, _04524_);
  nor (_31177_, _31176_, _31172_);
  nor (_31178_, _31177_, _03603_);
  or (_31179_, _31178_, _07441_);
  nor (_31180_, _31179_, _31162_);
  and (_31181_, _31174_, _07441_);
  nor (_31182_, _31181_, _31180_);
  nor (_31183_, _31182_, _05969_);
  nor (_31184_, _31183_, _03644_);
  and (_31185_, _31184_, _31158_);
  and (_31187_, _12330_, _05309_);
  or (_31188_, _31187_, _03275_);
  nor (_31189_, _31188_, _31159_);
  nor (_31190_, _31189_, _31185_);
  nor (_31191_, _31190_, _08861_);
  nor (_31192_, _12220_, _11178_);
  nor (_31193_, _31192_, _04591_);
  and (_31194_, _05309_, _04347_);
  nor (_31195_, _31194_, _04582_);
  nor (_31196_, _31195_, _31193_);
  nor (_31198_, _31196_, _31159_);
  nor (_31199_, _31198_, _31191_);
  nor (_31200_, _31199_, _03778_);
  nor (_31201_, _12347_, _11178_);
  or (_31202_, _31201_, _04589_);
  nor (_31203_, _31202_, _31159_);
  nor (_31204_, _31203_, _31200_);
  nor (_31205_, _31204_, _03655_);
  nor (_31206_, _12219_, _11178_);
  or (_31207_, _31206_, _04596_);
  nor (_31209_, _31207_, _31159_);
  nor (_31210_, _31209_, _31205_);
  nor (_31211_, _31210_, _03773_);
  nor (_31212_, _31154_, _05699_);
  nor (_31213_, _31212_, _04594_);
  and (_31214_, _31213_, _31161_);
  nor (_31215_, _31214_, _31211_);
  or (_31216_, _31215_, _18553_);
  nor (_31217_, _12218_, _11178_);
  or (_31218_, _31217_, _31154_);
  and (_31220_, _31218_, _03653_);
  not (_31221_, _31220_);
  and (_31222_, _12346_, _05309_);
  or (_31223_, _31222_, _04606_);
  nor (_31224_, _31223_, _31159_);
  nor (_31225_, _31224_, _03809_);
  and (_31226_, _31225_, _31221_);
  and (_31227_, _31226_, _31216_);
  nor (_31228_, _31169_, _04260_);
  nor (_31229_, _31228_, _31227_);
  and (_31231_, _31229_, _03820_);
  nor (_31232_, _31168_, _31154_);
  nor (_31233_, _31232_, _03820_);
  or (_31234_, _31233_, _31231_);
  or (_31235_, _31234_, _43231_);
  or (_31236_, _43227_, \oc8051_golden_model_1.TL1 [1]);
  and (_31237_, _31236_, _41991_);
  and (_43593_, _31237_, _31235_);
  not (_31238_, \oc8051_golden_model_1.TL1 [2]);
  nor (_31239_, _05309_, _31238_);
  nor (_31241_, _12543_, _11178_);
  nor (_31242_, _31241_, _31239_);
  nor (_31243_, _31242_, _04606_);
  nor (_31244_, _11178_, _05130_);
  nor (_31245_, _31244_, _31239_);
  and (_31246_, _31245_, _07441_);
  nor (_31247_, _12430_, _11178_);
  nor (_31248_, _31247_, _31239_);
  nor (_31249_, _31248_, _04515_);
  nor (_31250_, _04499_, _31238_);
  and (_31252_, _05309_, \oc8051_golden_model_1.ACC [2]);
  nor (_31253_, _31252_, _31239_);
  nor (_31254_, _31253_, _04500_);
  nor (_31255_, _31254_, _31250_);
  nor (_31256_, _31255_, _03599_);
  or (_31257_, _31256_, _31249_);
  and (_31258_, _31257_, _04524_);
  nor (_31259_, _31245_, _04524_);
  or (_31260_, _31259_, _31258_);
  and (_31261_, _31260_, _03611_);
  nor (_31263_, _31253_, _03611_);
  nor (_31264_, _31263_, _07441_);
  not (_31265_, _31264_);
  nor (_31266_, _31265_, _31261_);
  nor (_31267_, _31266_, _31246_);
  nor (_31268_, _31267_, _05969_);
  and (_31269_, _06839_, _05309_);
  nor (_31270_, _31239_, _05970_);
  not (_31271_, _31270_);
  nor (_31272_, _31271_, _31269_);
  nor (_31274_, _31272_, _31268_);
  nor (_31275_, _31274_, _03644_);
  nor (_31276_, _12524_, _11178_);
  or (_31277_, _31239_, _03275_);
  nor (_31278_, _31277_, _31276_);
  or (_31279_, _31278_, _03650_);
  nor (_31280_, _31279_, _31275_);
  and (_31281_, _05309_, _06414_);
  nor (_31282_, _31281_, _31239_);
  nor (_31283_, _31282_, _04582_);
  or (_31285_, _31283_, _31280_);
  and (_31286_, _31285_, _04591_);
  and (_31287_, _12538_, _05309_);
  nor (_31288_, _31287_, _31239_);
  nor (_31289_, _31288_, _04591_);
  or (_31290_, _31289_, _31286_);
  nor (_31291_, _31290_, _03778_);
  and (_31292_, _12544_, _05309_);
  or (_31293_, _31239_, _04589_);
  nor (_31294_, _31293_, _31292_);
  or (_31296_, _31294_, _03655_);
  nor (_31297_, _31296_, _31291_);
  nor (_31298_, _31239_, _05793_);
  or (_31299_, _31282_, _04596_);
  nor (_31300_, _31299_, _31298_);
  nor (_31301_, _31300_, _31297_);
  nor (_31302_, _31301_, _03773_);
  or (_31303_, _31298_, _04594_);
  or (_31304_, _31303_, _31253_);
  and (_31305_, _31304_, _04608_);
  not (_31307_, _31305_);
  nor (_31308_, _31307_, _31302_);
  nor (_31309_, _12537_, _11178_);
  or (_31310_, _31239_, _04608_);
  nor (_31311_, _31310_, _31309_);
  or (_31312_, _31311_, _03786_);
  nor (_31313_, _31312_, _31308_);
  nor (_31314_, _31313_, _31243_);
  nor (_31315_, _31314_, _03809_);
  nor (_31316_, _31248_, _04260_);
  or (_31318_, _31316_, _03816_);
  nor (_31319_, _31318_, _31315_);
  and (_31320_, _12600_, _05309_);
  or (_31321_, _31239_, _03820_);
  nor (_31322_, _31321_, _31320_);
  nor (_31323_, _31322_, _31319_);
  or (_31324_, _31323_, _43231_);
  or (_31325_, _43227_, \oc8051_golden_model_1.TL1 [2]);
  and (_31326_, _31325_, _41991_);
  and (_43594_, _31326_, _31324_);
  not (_31328_, \oc8051_golden_model_1.TL1 [3]);
  nor (_31329_, _05309_, _31328_);
  nor (_31330_, _12618_, _11178_);
  nor (_31331_, _31330_, _31329_);
  nor (_31332_, _31331_, _04606_);
  and (_31333_, _12619_, _05309_);
  nor (_31334_, _31333_, _31329_);
  nor (_31335_, _31334_, _04589_);
  and (_31336_, _06838_, _05309_);
  or (_31337_, _31336_, _31329_);
  and (_31339_, _31337_, _05969_);
  and (_31340_, _05309_, \oc8051_golden_model_1.ACC [3]);
  nor (_31341_, _31340_, _31329_);
  nor (_31342_, _31341_, _03611_);
  nor (_31343_, _31341_, _04500_);
  nor (_31344_, _04499_, _31328_);
  or (_31345_, _31344_, _31343_);
  and (_31346_, _31345_, _04515_);
  nor (_31347_, _12625_, _11178_);
  nor (_31348_, _31347_, _31329_);
  nor (_31350_, _31348_, _04515_);
  or (_31351_, _31350_, _31346_);
  and (_31352_, _31351_, _04524_);
  nor (_31353_, _11178_, _04944_);
  nor (_31354_, _31353_, _31329_);
  nor (_31355_, _31354_, _04524_);
  nor (_31356_, _31355_, _31352_);
  nor (_31357_, _31356_, _03603_);
  or (_31358_, _31357_, _07441_);
  nor (_31359_, _31358_, _31342_);
  and (_31361_, _31354_, _07441_);
  or (_31362_, _31361_, _05969_);
  nor (_31363_, _31362_, _31359_);
  or (_31364_, _31363_, _31339_);
  and (_31365_, _31364_, _03275_);
  nor (_31366_, _12731_, _11178_);
  nor (_31367_, _31366_, _31329_);
  nor (_31368_, _31367_, _03275_);
  or (_31369_, _31368_, _08861_);
  or (_31370_, _31369_, _31365_);
  and (_31372_, _12746_, _05309_);
  or (_31373_, _31329_, _04591_);
  or (_31374_, _31373_, _31372_);
  and (_31375_, _05309_, _06347_);
  nor (_31376_, _31375_, _31329_);
  and (_31377_, _31376_, _03650_);
  nor (_31378_, _31377_, _03778_);
  and (_31379_, _31378_, _31374_);
  and (_31380_, _31379_, _31370_);
  nor (_31381_, _31380_, _31335_);
  nor (_31383_, _31381_, _03655_);
  nor (_31384_, _31329_, _05650_);
  not (_31385_, _31384_);
  nor (_31386_, _31376_, _04596_);
  and (_31387_, _31386_, _31385_);
  nor (_31388_, _31387_, _31383_);
  nor (_31389_, _31388_, _03773_);
  nor (_31390_, _31341_, _04594_);
  and (_31391_, _31390_, _31385_);
  nor (_31392_, _31391_, _03653_);
  not (_31394_, _31392_);
  nor (_31395_, _31394_, _31389_);
  nor (_31396_, _12745_, _11178_);
  or (_31397_, _31329_, _04608_);
  nor (_31398_, _31397_, _31396_);
  or (_31399_, _31398_, _03786_);
  nor (_31400_, _31399_, _31395_);
  nor (_31401_, _31400_, _31332_);
  nor (_31402_, _31401_, _03809_);
  nor (_31403_, _31348_, _04260_);
  or (_31405_, _31403_, _03816_);
  nor (_31406_, _31405_, _31402_);
  and (_31407_, _12806_, _05309_);
  or (_31408_, _31329_, _03820_);
  nor (_31409_, _31408_, _31407_);
  nor (_31410_, _31409_, _31406_);
  or (_31411_, _31410_, _43231_);
  or (_31412_, _43227_, \oc8051_golden_model_1.TL1 [3]);
  and (_31413_, _31412_, _41991_);
  and (_43595_, _31413_, _31411_);
  not (_31415_, \oc8051_golden_model_1.TL1 [4]);
  nor (_31416_, _05309_, _31415_);
  nor (_31417_, _12956_, _11178_);
  nor (_31418_, _31417_, _31416_);
  nor (_31419_, _31418_, _04606_);
  and (_31420_, _12957_, _05309_);
  nor (_31421_, _31420_, _31416_);
  nor (_31422_, _31421_, _04589_);
  and (_31423_, _06375_, _05309_);
  nor (_31424_, _31423_, _31416_);
  and (_31426_, _31424_, _03650_);
  nor (_31427_, _05840_, _11178_);
  nor (_31428_, _31427_, _31416_);
  and (_31429_, _31428_, _07441_);
  and (_31430_, _05309_, \oc8051_golden_model_1.ACC [4]);
  nor (_31431_, _31430_, _31416_);
  nor (_31432_, _31431_, _03611_);
  nor (_31433_, _31431_, _04500_);
  nor (_31434_, _04499_, _31415_);
  or (_31435_, _31434_, _31433_);
  and (_31437_, _31435_, _04515_);
  nor (_31438_, _12820_, _11178_);
  nor (_31439_, _31438_, _31416_);
  nor (_31440_, _31439_, _04515_);
  or (_31441_, _31440_, _31437_);
  and (_31442_, _31441_, _04524_);
  nor (_31443_, _31428_, _04524_);
  nor (_31444_, _31443_, _31442_);
  nor (_31445_, _31444_, _03603_);
  or (_31446_, _31445_, _07441_);
  nor (_31448_, _31446_, _31432_);
  nor (_31449_, _31448_, _31429_);
  nor (_31450_, _31449_, _05969_);
  and (_31451_, _06843_, _05309_);
  nor (_31452_, _31416_, _05970_);
  not (_31453_, _31452_);
  nor (_31454_, _31453_, _31451_);
  or (_31455_, _31454_, _03644_);
  nor (_31456_, _31455_, _31450_);
  nor (_31457_, _12936_, _11178_);
  nor (_31459_, _31457_, _31416_);
  nor (_31460_, _31459_, _03275_);
  or (_31461_, _31460_, _03650_);
  nor (_31462_, _31461_, _31456_);
  nor (_31463_, _31462_, _31426_);
  or (_31464_, _31463_, _03649_);
  and (_31465_, _12951_, _05309_);
  or (_31466_, _31465_, _31416_);
  or (_31467_, _31466_, _04591_);
  and (_31468_, _31467_, _04589_);
  and (_31470_, _31468_, _31464_);
  nor (_31471_, _31470_, _31422_);
  nor (_31472_, _31471_, _03655_);
  nor (_31473_, _31416_, _05889_);
  not (_31474_, _31473_);
  nor (_31475_, _31424_, _04596_);
  and (_31476_, _31475_, _31474_);
  nor (_31477_, _31476_, _31472_);
  nor (_31478_, _31477_, _03773_);
  nor (_31479_, _31431_, _04594_);
  and (_31481_, _31479_, _31474_);
  nor (_31482_, _31481_, _03653_);
  not (_31483_, _31482_);
  nor (_31484_, _31483_, _31478_);
  nor (_31485_, _12949_, _11178_);
  or (_31486_, _31416_, _04608_);
  nor (_31487_, _31486_, _31485_);
  or (_31488_, _31487_, _03786_);
  nor (_31489_, _31488_, _31484_);
  nor (_31490_, _31489_, _31419_);
  nor (_31492_, _31490_, _03809_);
  nor (_31493_, _31439_, _04260_);
  or (_31494_, _31493_, _03816_);
  nor (_31495_, _31494_, _31492_);
  and (_31496_, _13013_, _05309_);
  or (_31497_, _31416_, _03820_);
  nor (_31498_, _31497_, _31496_);
  nor (_31499_, _31498_, _31495_);
  or (_31500_, _31499_, _43231_);
  or (_31501_, _43227_, \oc8051_golden_model_1.TL1 [4]);
  and (_31503_, _31501_, _41991_);
  and (_43596_, _31503_, _31500_);
  not (_31504_, \oc8051_golden_model_1.TL1 [5]);
  nor (_31505_, _05309_, _31504_);
  nor (_31506_, _13159_, _11178_);
  nor (_31507_, _31506_, _31505_);
  nor (_31508_, _31507_, _04606_);
  and (_31509_, _13160_, _05309_);
  nor (_31510_, _31509_, _31505_);
  nor (_31511_, _31510_, _04589_);
  and (_31513_, _06842_, _05309_);
  or (_31514_, _31513_, _31505_);
  and (_31515_, _31514_, _05969_);
  and (_31516_, _05309_, \oc8051_golden_model_1.ACC [5]);
  nor (_31517_, _31516_, _31505_);
  nor (_31518_, _31517_, _03611_);
  nor (_31519_, _31517_, _04500_);
  nor (_31520_, _04499_, _31504_);
  or (_31521_, _31520_, _31519_);
  and (_31522_, _31521_, _04515_);
  nor (_31524_, _13035_, _11178_);
  nor (_31525_, _31524_, _31505_);
  nor (_31526_, _31525_, _04515_);
  or (_31527_, _31526_, _31522_);
  and (_31528_, _31527_, _04524_);
  nor (_31529_, _05552_, _11178_);
  nor (_31530_, _31529_, _31505_);
  nor (_31531_, _31530_, _04524_);
  nor (_31532_, _31531_, _31528_);
  nor (_31533_, _31532_, _03603_);
  or (_31535_, _31533_, _07441_);
  nor (_31536_, _31535_, _31518_);
  and (_31537_, _31530_, _07441_);
  or (_31538_, _31537_, _05969_);
  nor (_31539_, _31538_, _31536_);
  or (_31540_, _31539_, _31515_);
  and (_31541_, _31540_, _03275_);
  nor (_31542_, _13139_, _11178_);
  nor (_31543_, _31542_, _31505_);
  nor (_31544_, _31543_, _03275_);
  or (_31545_, _31544_, _08861_);
  or (_31546_, _31545_, _31541_);
  and (_31547_, _13154_, _05309_);
  or (_31548_, _31505_, _04591_);
  or (_31549_, _31548_, _31547_);
  and (_31550_, _06358_, _05309_);
  nor (_31551_, _31550_, _31505_);
  and (_31552_, _31551_, _03650_);
  nor (_31553_, _31552_, _03778_);
  and (_31554_, _31553_, _31549_);
  and (_31556_, _31554_, _31546_);
  nor (_31557_, _31556_, _31511_);
  nor (_31558_, _31557_, _03655_);
  nor (_31559_, _31505_, _05601_);
  not (_31560_, _31559_);
  nor (_31561_, _31551_, _04596_);
  and (_31562_, _31561_, _31560_);
  nor (_31563_, _31562_, _31558_);
  nor (_31564_, _31563_, _03773_);
  nor (_31565_, _31517_, _04594_);
  and (_31567_, _31565_, _31560_);
  nor (_31568_, _31567_, _03653_);
  not (_31569_, _31568_);
  nor (_31570_, _31569_, _31564_);
  nor (_31571_, _13152_, _11178_);
  or (_31572_, _31505_, _04608_);
  nor (_31573_, _31572_, _31571_);
  or (_31574_, _31573_, _03786_);
  nor (_31575_, _31574_, _31570_);
  nor (_31576_, _31575_, _31508_);
  nor (_31578_, _31576_, _03809_);
  nor (_31579_, _31525_, _04260_);
  or (_31580_, _31579_, _03816_);
  nor (_31581_, _31580_, _31578_);
  and (_31582_, _13217_, _05309_);
  or (_31583_, _31505_, _03820_);
  nor (_31584_, _31583_, _31582_);
  nor (_31585_, _31584_, _31581_);
  or (_31586_, _31585_, _43231_);
  or (_31587_, _43227_, \oc8051_golden_model_1.TL1 [5]);
  and (_31589_, _31587_, _41991_);
  and (_43597_, _31589_, _31586_);
  not (_31590_, \oc8051_golden_model_1.TL1 [6]);
  nor (_31591_, _05309_, _31590_);
  nor (_31592_, _13373_, _11178_);
  nor (_31593_, _31592_, _31591_);
  nor (_31594_, _31593_, _04606_);
  and (_31595_, _13374_, _05309_);
  nor (_31596_, _31595_, _31591_);
  nor (_31597_, _31596_, _04589_);
  and (_31599_, _06531_, _05309_);
  or (_31600_, _31599_, _31591_);
  and (_31601_, _31600_, _05969_);
  and (_31602_, _05309_, \oc8051_golden_model_1.ACC [6]);
  nor (_31603_, _31602_, _31591_);
  nor (_31604_, _31603_, _03611_);
  nor (_31605_, _31603_, _04500_);
  nor (_31606_, _04499_, _31590_);
  or (_31607_, _31606_, _31605_);
  and (_31608_, _31607_, _04515_);
  nor (_31610_, _13235_, _11178_);
  nor (_31611_, _31610_, _31591_);
  nor (_31612_, _31611_, _04515_);
  or (_31613_, _31612_, _31608_);
  and (_31614_, _31613_, _04524_);
  nor (_31615_, _05442_, _11178_);
  nor (_31616_, _31615_, _31591_);
  nor (_31617_, _31616_, _04524_);
  nor (_31618_, _31617_, _31614_);
  nor (_31619_, _31618_, _03603_);
  or (_31621_, _31619_, _07441_);
  nor (_31622_, _31621_, _31604_);
  and (_31623_, _31616_, _07441_);
  or (_31624_, _31623_, _05969_);
  nor (_31625_, _31624_, _31622_);
  or (_31626_, _31625_, _31601_);
  and (_31627_, _31626_, _03275_);
  nor (_31628_, _13356_, _11178_);
  nor (_31629_, _31628_, _31591_);
  nor (_31630_, _31629_, _03275_);
  or (_31632_, _31630_, _08861_);
  or (_31633_, _31632_, _31627_);
  and (_31634_, _13245_, _05309_);
  or (_31635_, _31591_, _04591_);
  or (_31636_, _31635_, _31634_);
  and (_31637_, _13363_, _05309_);
  nor (_31638_, _31637_, _31591_);
  and (_31639_, _31638_, _03650_);
  nor (_31640_, _31639_, _03778_);
  and (_31641_, _31640_, _31636_);
  and (_31643_, _31641_, _31633_);
  nor (_31644_, _31643_, _31597_);
  nor (_31645_, _31644_, _03655_);
  nor (_31646_, _31591_, _05491_);
  not (_31647_, _31646_);
  nor (_31648_, _31638_, _04596_);
  and (_31649_, _31648_, _31647_);
  nor (_31650_, _31649_, _31645_);
  nor (_31651_, _31650_, _03773_);
  nor (_31652_, _31603_, _04594_);
  and (_31654_, _31652_, _31647_);
  or (_31655_, _31654_, _31651_);
  and (_31656_, _31655_, _04608_);
  nor (_31657_, _13243_, _11178_);
  nor (_31658_, _31657_, _31591_);
  nor (_31659_, _31658_, _04608_);
  or (_31660_, _31659_, _31656_);
  and (_31661_, _31660_, _04606_);
  nor (_31662_, _31661_, _31594_);
  nor (_31663_, _31662_, _03809_);
  nor (_31665_, _31611_, _04260_);
  or (_31666_, _31665_, _03816_);
  nor (_31667_, _31666_, _31663_);
  and (_31668_, _13425_, _05309_);
  or (_31669_, _31591_, _03820_);
  nor (_31670_, _31669_, _31668_);
  nor (_31671_, _31670_, _31667_);
  or (_31672_, _31671_, _43231_);
  or (_31673_, _43227_, \oc8051_golden_model_1.TL1 [6]);
  and (_31674_, _31673_, _41991_);
  and (_43598_, _31674_, _31672_);
  not (_31675_, \oc8051_golden_model_1.TMOD [0]);
  nor (_31676_, _05343_, _31675_);
  nor (_31677_, _05744_, _11261_);
  nor (_31678_, _31677_, _31676_);
  and (_31679_, _31678_, _17220_);
  and (_31680_, _05343_, \oc8051_golden_model_1.ACC [0]);
  nor (_31681_, _31680_, _31676_);
  nor (_31682_, _31681_, _03611_);
  nor (_31683_, _31682_, _07441_);
  nor (_31686_, _31678_, _04515_);
  nor (_31687_, _04499_, _31675_);
  nor (_31688_, _31681_, _04500_);
  nor (_31689_, _31688_, _31687_);
  nor (_31690_, _31689_, _03599_);
  or (_31691_, _31690_, _03597_);
  nor (_31692_, _31691_, _31686_);
  or (_31693_, _31692_, _03603_);
  and (_31694_, _31693_, _31683_);
  and (_31695_, _05343_, _04491_);
  or (_31697_, _31676_, _26194_);
  nor (_31698_, _31697_, _31695_);
  nor (_31699_, _31698_, _31694_);
  nor (_31700_, _31699_, _05969_);
  and (_31701_, _06836_, _05343_);
  nor (_31702_, _31676_, _05970_);
  not (_31703_, _31702_);
  nor (_31704_, _31703_, _31701_);
  nor (_31705_, _31704_, _31700_);
  nor (_31706_, _31705_, _03644_);
  nor (_31708_, _12129_, _11261_);
  or (_31709_, _31676_, _03275_);
  nor (_31710_, _31709_, _31708_);
  or (_31711_, _31710_, _03650_);
  nor (_31712_, _31711_, _31706_);
  and (_31713_, _05343_, _06366_);
  nor (_31714_, _31713_, _31676_);
  nor (_31715_, _31714_, _04582_);
  or (_31716_, _31715_, _31712_);
  and (_31717_, _31716_, _04591_);
  and (_31719_, _12019_, _05343_);
  nor (_31720_, _31719_, _31676_);
  nor (_31721_, _31720_, _04591_);
  or (_31722_, _31721_, _31717_);
  nor (_31723_, _31722_, _03778_);
  and (_31724_, _12145_, _05343_);
  or (_31725_, _31676_, _04589_);
  nor (_31726_, _31725_, _31724_);
  or (_31727_, _31726_, _03655_);
  nor (_31728_, _31727_, _31723_);
  or (_31730_, _31714_, _04596_);
  nor (_31731_, _31730_, _31677_);
  nor (_31732_, _31731_, _31728_);
  nor (_31733_, _31732_, _03773_);
  and (_31734_, _12144_, _05343_);
  or (_31735_, _31734_, _31676_);
  and (_31736_, _31735_, _03773_);
  or (_31737_, _31736_, _31733_);
  and (_31738_, _31737_, _04608_);
  nor (_31739_, _12017_, _11261_);
  nor (_31741_, _31739_, _31676_);
  nor (_31742_, _31741_, _04608_);
  or (_31743_, _31742_, _31738_);
  and (_31744_, _31743_, _04606_);
  nor (_31745_, _12015_, _11261_);
  nor (_31746_, _31745_, _31676_);
  nor (_31747_, _31746_, _04606_);
  nor (_31748_, _31747_, _17220_);
  not (_31749_, _31748_);
  nor (_31750_, _31749_, _31744_);
  nor (_31752_, _31750_, _31679_);
  or (_31753_, _31752_, _43231_);
  or (_31754_, _43227_, \oc8051_golden_model_1.TMOD [0]);
  and (_31755_, _31754_, _41991_);
  and (_43600_, _31755_, _31753_);
  and (_31756_, _06835_, _05343_);
  not (_31757_, \oc8051_golden_model_1.TMOD [1]);
  nor (_31758_, _05343_, _31757_);
  nor (_31759_, _31758_, _05970_);
  not (_31760_, _31759_);
  nor (_31762_, _31760_, _31756_);
  not (_31763_, _31762_);
  and (_31764_, _05343_, _05898_);
  nor (_31765_, _31764_, _31758_);
  and (_31766_, _31765_, _07441_);
  nor (_31767_, _05343_, \oc8051_golden_model_1.TMOD [1]);
  and (_31768_, _05343_, _03320_);
  nor (_31769_, _31768_, _31767_);
  and (_31770_, _31769_, _04499_);
  nor (_31771_, _04499_, _31757_);
  or (_31773_, _31771_, _31770_);
  and (_31774_, _31773_, _04515_);
  and (_31775_, _12234_, _05343_);
  nor (_31776_, _31775_, _31767_);
  and (_31777_, _31776_, _03599_);
  or (_31778_, _31777_, _31774_);
  and (_31779_, _31778_, _04524_);
  nor (_31780_, _31765_, _04524_);
  nor (_31781_, _31780_, _31779_);
  nor (_31782_, _31781_, _03603_);
  and (_31784_, _31769_, _03603_);
  nor (_31785_, _31784_, _07441_);
  not (_31786_, _31785_);
  nor (_31787_, _31786_, _31782_);
  nor (_31788_, _31787_, _31766_);
  nor (_31789_, _31788_, _05969_);
  nor (_31790_, _31789_, _03644_);
  and (_31791_, _31790_, _31763_);
  not (_31792_, _31767_);
  and (_31793_, _12330_, _05343_);
  nor (_31795_, _31793_, _03275_);
  and (_31796_, _31795_, _31792_);
  nor (_31797_, _31796_, _31791_);
  nor (_31798_, _31797_, _08861_);
  nor (_31799_, _12220_, _11261_);
  nor (_31800_, _31799_, _04591_);
  and (_31801_, _05343_, _04347_);
  nor (_31802_, _31801_, _04582_);
  or (_31803_, _31802_, _31800_);
  and (_31804_, _31803_, _31792_);
  nor (_31806_, _31804_, _31798_);
  nor (_31807_, _31806_, _03778_);
  nor (_31808_, _12347_, _11261_);
  nor (_31809_, _31808_, _04589_);
  and (_31810_, _31809_, _31792_);
  nor (_31811_, _31810_, _31807_);
  nor (_31812_, _31811_, _03655_);
  nor (_31813_, _12219_, _11261_);
  nor (_31814_, _31813_, _04596_);
  and (_31815_, _31814_, _31792_);
  nor (_31817_, _31815_, _31812_);
  nor (_31818_, _31817_, _03773_);
  nor (_31819_, _31758_, _05699_);
  nor (_31820_, _31819_, _04594_);
  and (_31821_, _31820_, _31769_);
  nor (_31822_, _31821_, _31818_);
  or (_31823_, _31822_, _18553_);
  and (_31824_, _31801_, _05698_);
  nor (_31825_, _31824_, _04608_);
  and (_31826_, _31825_, _31792_);
  nand (_31828_, _31768_, _05698_);
  nor (_31829_, _31767_, _04606_);
  and (_31830_, _31829_, _31828_);
  or (_31831_, _31830_, _03809_);
  nor (_31832_, _31831_, _31826_);
  and (_31833_, _31832_, _31823_);
  nor (_31834_, _31776_, _04260_);
  nor (_31835_, _31834_, _31833_);
  and (_31836_, _31835_, _03820_);
  nor (_31837_, _31775_, _31758_);
  nor (_31839_, _31837_, _03820_);
  or (_31840_, _31839_, _31836_);
  or (_31841_, _31840_, _43231_);
  or (_31842_, _43227_, \oc8051_golden_model_1.TMOD [1]);
  and (_31843_, _31842_, _41991_);
  and (_43601_, _31843_, _31841_);
  not (_31844_, \oc8051_golden_model_1.TMOD [2]);
  nor (_31845_, _05343_, _31844_);
  nor (_31846_, _12543_, _11261_);
  nor (_31847_, _31846_, _31845_);
  nor (_31849_, _31847_, _04606_);
  nor (_31850_, _11261_, _05130_);
  nor (_31851_, _31850_, _31845_);
  and (_31852_, _31851_, _07441_);
  nor (_31853_, _12430_, _11261_);
  nor (_31854_, _31853_, _31845_);
  nor (_31855_, _31854_, _04515_);
  nor (_31856_, _04499_, _31844_);
  and (_31857_, _05343_, \oc8051_golden_model_1.ACC [2]);
  nor (_31858_, _31857_, _31845_);
  nor (_31860_, _31858_, _04500_);
  nor (_31861_, _31860_, _31856_);
  nor (_31862_, _31861_, _03599_);
  or (_31863_, _31862_, _31855_);
  and (_31864_, _31863_, _04524_);
  nor (_31865_, _31851_, _04524_);
  or (_31866_, _31865_, _31864_);
  and (_31867_, _31866_, _03611_);
  nor (_31868_, _31858_, _03611_);
  nor (_31869_, _31868_, _07441_);
  not (_31871_, _31869_);
  nor (_31872_, _31871_, _31867_);
  nor (_31873_, _31872_, _31852_);
  nor (_31874_, _31873_, _05969_);
  and (_31875_, _06839_, _05343_);
  nor (_31876_, _31845_, _05970_);
  not (_31877_, _31876_);
  nor (_31878_, _31877_, _31875_);
  nor (_31879_, _31878_, _31874_);
  nor (_31880_, _31879_, _03644_);
  nor (_31882_, _12524_, _11261_);
  or (_31883_, _31845_, _03275_);
  nor (_31884_, _31883_, _31882_);
  or (_31885_, _31884_, _03650_);
  nor (_31886_, _31885_, _31880_);
  and (_31887_, _05343_, _06414_);
  nor (_31888_, _31887_, _31845_);
  nor (_31889_, _31888_, _04582_);
  or (_31890_, _31889_, _31886_);
  and (_31891_, _31890_, _04591_);
  and (_31893_, _12538_, _05343_);
  nor (_31894_, _31893_, _31845_);
  nor (_31895_, _31894_, _04591_);
  or (_31896_, _31895_, _31891_);
  nor (_31897_, _31896_, _03778_);
  and (_31898_, _12544_, _05343_);
  or (_31899_, _31845_, _04589_);
  nor (_31900_, _31899_, _31898_);
  or (_31901_, _31900_, _03655_);
  nor (_31902_, _31901_, _31897_);
  nor (_31904_, _31845_, _05793_);
  or (_31905_, _31888_, _04596_);
  nor (_31906_, _31905_, _31904_);
  nor (_31907_, _31906_, _31902_);
  nor (_31908_, _31907_, _03773_);
  or (_31909_, _31904_, _04594_);
  or (_31910_, _31909_, _31858_);
  and (_31911_, _31910_, _04608_);
  not (_31912_, _31911_);
  nor (_31913_, _31912_, _31908_);
  nor (_31915_, _12537_, _11261_);
  or (_31916_, _31845_, _04608_);
  nor (_31917_, _31916_, _31915_);
  or (_31918_, _31917_, _03786_);
  nor (_31919_, _31918_, _31913_);
  nor (_31920_, _31919_, _31849_);
  nor (_31921_, _31920_, _03809_);
  nor (_31922_, _31854_, _04260_);
  or (_31923_, _31922_, _03816_);
  nor (_31924_, _31923_, _31921_);
  and (_31926_, _12600_, _05343_);
  or (_31927_, _31845_, _03820_);
  nor (_31928_, _31927_, _31926_);
  nor (_31929_, _31928_, _31924_);
  or (_31930_, _31929_, _43231_);
  or (_31931_, _43227_, \oc8051_golden_model_1.TMOD [2]);
  and (_31932_, _31931_, _41991_);
  and (_43602_, _31932_, _31930_);
  not (_31933_, \oc8051_golden_model_1.TMOD [3]);
  nor (_31934_, _05343_, _31933_);
  nor (_31936_, _12618_, _11261_);
  nor (_31937_, _31936_, _31934_);
  nor (_31938_, _31937_, _04606_);
  and (_31939_, _06838_, _05343_);
  nor (_31940_, _31939_, _31934_);
  or (_31941_, _31940_, _05970_);
  and (_31942_, _05343_, \oc8051_golden_model_1.ACC [3]);
  nor (_31943_, _31942_, _31934_);
  nor (_31944_, _31943_, _04500_);
  nor (_31945_, _04499_, _31933_);
  or (_31947_, _31945_, _31944_);
  and (_31948_, _31947_, _04515_);
  nor (_31949_, _12625_, _11261_);
  nor (_31950_, _31949_, _31934_);
  nor (_31951_, _31950_, _04515_);
  or (_31952_, _31951_, _31948_);
  and (_31953_, _31952_, _04524_);
  nor (_31954_, _11261_, _04944_);
  nor (_31955_, _31954_, _31934_);
  nor (_31956_, _31955_, _04524_);
  nor (_31958_, _31956_, _31953_);
  nor (_31959_, _31958_, _03603_);
  nor (_31960_, _31943_, _03611_);
  nor (_31961_, _31960_, _07441_);
  not (_31962_, _31961_);
  nor (_31963_, _31962_, _31959_);
  and (_31964_, _31955_, _07441_);
  or (_31965_, _31964_, _05969_);
  or (_31966_, _31965_, _31963_);
  and (_31967_, _31966_, _03275_);
  and (_31969_, _31967_, _31941_);
  nor (_31970_, _12731_, _11261_);
  or (_31971_, _31934_, _03275_);
  nor (_31972_, _31971_, _31970_);
  or (_31973_, _31972_, _03650_);
  nor (_31974_, _31973_, _31969_);
  and (_31975_, _05343_, _06347_);
  nor (_31976_, _31975_, _31934_);
  nor (_31977_, _31976_, _04582_);
  or (_31978_, _31977_, _31974_);
  and (_31980_, _31978_, _04591_);
  and (_31981_, _12746_, _05343_);
  nor (_31982_, _31981_, _31934_);
  nor (_31983_, _31982_, _04591_);
  or (_31984_, _31983_, _31980_);
  nor (_31985_, _31984_, _03778_);
  and (_31986_, _12619_, _05343_);
  or (_31987_, _31934_, _04589_);
  nor (_31988_, _31987_, _31986_);
  or (_31989_, _31988_, _03655_);
  nor (_31991_, _31989_, _31985_);
  nor (_31992_, _31934_, _05650_);
  or (_31993_, _31976_, _04596_);
  nor (_31994_, _31993_, _31992_);
  nor (_31995_, _31994_, _31991_);
  nor (_31996_, _31995_, _03773_);
  or (_31997_, _31992_, _04594_);
  nor (_31998_, _31997_, _31943_);
  or (_31999_, _31998_, _31996_);
  and (_32000_, _31999_, _04608_);
  nor (_32002_, _12745_, _11261_);
  nor (_32003_, _32002_, _31934_);
  nor (_32004_, _32003_, _04608_);
  or (_32005_, _32004_, _32000_);
  and (_32006_, _32005_, _04606_);
  nor (_32007_, _32006_, _31938_);
  nor (_32008_, _32007_, _03809_);
  nor (_32009_, _31950_, _04260_);
  or (_32010_, _32009_, _03816_);
  nor (_32011_, _32010_, _32008_);
  and (_32013_, _12806_, _05343_);
  or (_32014_, _31934_, _03820_);
  nor (_32015_, _32014_, _32013_);
  nor (_32016_, _32015_, _32011_);
  or (_32017_, _32016_, _43231_);
  or (_32018_, _43227_, \oc8051_golden_model_1.TMOD [3]);
  and (_32019_, _32018_, _41991_);
  and (_43604_, _32019_, _32017_);
  not (_32020_, \oc8051_golden_model_1.TMOD [4]);
  nor (_32021_, _05343_, _32020_);
  nor (_32023_, _12956_, _11261_);
  nor (_32024_, _32023_, _32021_);
  nor (_32025_, _32024_, _04606_);
  and (_32026_, _12957_, _05343_);
  nor (_32027_, _32026_, _32021_);
  nor (_32028_, _32027_, _04589_);
  and (_32029_, _06375_, _05343_);
  nor (_32030_, _32029_, _32021_);
  and (_32031_, _32030_, _03650_);
  and (_32032_, _05343_, \oc8051_golden_model_1.ACC [4]);
  nor (_32034_, _32032_, _32021_);
  nor (_32035_, _32034_, _03611_);
  nor (_32036_, _32034_, _04500_);
  nor (_32037_, _04499_, _32020_);
  or (_32038_, _32037_, _32036_);
  and (_32039_, _32038_, _04515_);
  nor (_32040_, _12820_, _11261_);
  nor (_32041_, _32040_, _32021_);
  nor (_32042_, _32041_, _04515_);
  or (_32043_, _32042_, _32039_);
  and (_32045_, _32043_, _04524_);
  nor (_32046_, _05840_, _11261_);
  nor (_32047_, _32046_, _32021_);
  nor (_32048_, _32047_, _04524_);
  nor (_32049_, _32048_, _32045_);
  nor (_32050_, _32049_, _03603_);
  or (_32051_, _32050_, _07441_);
  nor (_32052_, _32051_, _32035_);
  and (_32053_, _32047_, _07441_);
  nor (_32054_, _32053_, _32052_);
  nor (_32056_, _32054_, _05969_);
  and (_32057_, _06843_, _05343_);
  nor (_32058_, _32021_, _05970_);
  not (_32059_, _32058_);
  nor (_32060_, _32059_, _32057_);
  or (_32061_, _32060_, _03644_);
  nor (_32062_, _32061_, _32056_);
  nor (_32063_, _12936_, _11261_);
  nor (_32064_, _32063_, _32021_);
  nor (_32065_, _32064_, _03275_);
  or (_32067_, _32065_, _03650_);
  nor (_32068_, _32067_, _32062_);
  nor (_32069_, _32068_, _32031_);
  or (_32070_, _32069_, _03649_);
  and (_32071_, _12951_, _05343_);
  or (_32072_, _32071_, _32021_);
  or (_32073_, _32072_, _04591_);
  and (_32074_, _32073_, _04589_);
  and (_32075_, _32074_, _32070_);
  nor (_32076_, _32075_, _32028_);
  nor (_32078_, _32076_, _03655_);
  nor (_32079_, _32021_, _05889_);
  not (_32080_, _32079_);
  nor (_32081_, _32030_, _04596_);
  and (_32082_, _32081_, _32080_);
  nor (_32083_, _32082_, _32078_);
  nor (_32084_, _32083_, _03773_);
  nor (_32085_, _32034_, _04594_);
  and (_32086_, _32085_, _32080_);
  nor (_32087_, _32086_, _03653_);
  not (_32089_, _32087_);
  nor (_32090_, _32089_, _32084_);
  nor (_32091_, _12949_, _11261_);
  or (_32092_, _32021_, _04608_);
  nor (_32093_, _32092_, _32091_);
  or (_32094_, _32093_, _03786_);
  nor (_32095_, _32094_, _32090_);
  nor (_32096_, _32095_, _32025_);
  nor (_32097_, _32096_, _03809_);
  nor (_32098_, _32041_, _04260_);
  or (_32100_, _32098_, _03816_);
  nor (_32101_, _32100_, _32097_);
  and (_32102_, _13013_, _05343_);
  or (_32103_, _32021_, _03820_);
  nor (_32104_, _32103_, _32102_);
  nor (_32105_, _32104_, _32101_);
  or (_32106_, _32105_, _43231_);
  or (_32107_, _43227_, \oc8051_golden_model_1.TMOD [4]);
  and (_32108_, _32107_, _41991_);
  and (_43605_, _32108_, _32106_);
  not (_32110_, \oc8051_golden_model_1.TMOD [5]);
  nor (_32111_, _05343_, _32110_);
  nor (_32112_, _13159_, _11261_);
  nor (_32113_, _32112_, _32111_);
  nor (_32114_, _32113_, _04606_);
  and (_32115_, _13160_, _05343_);
  nor (_32116_, _32115_, _32111_);
  nor (_32117_, _32116_, _04589_);
  and (_32118_, _06842_, _05343_);
  or (_32119_, _32118_, _32111_);
  and (_32121_, _32119_, _05969_);
  and (_32122_, _05343_, \oc8051_golden_model_1.ACC [5]);
  nor (_32123_, _32122_, _32111_);
  nor (_32124_, _32123_, _03611_);
  nor (_32125_, _32123_, _04500_);
  nor (_32126_, _04499_, _32110_);
  or (_32127_, _32126_, _32125_);
  and (_32128_, _32127_, _04515_);
  nor (_32129_, _13035_, _11261_);
  nor (_32130_, _32129_, _32111_);
  nor (_32132_, _32130_, _04515_);
  or (_32133_, _32132_, _32128_);
  and (_32134_, _32133_, _04524_);
  nor (_32135_, _05552_, _11261_);
  nor (_32136_, _32135_, _32111_);
  nor (_32137_, _32136_, _04524_);
  nor (_32138_, _32137_, _32134_);
  nor (_32139_, _32138_, _03603_);
  or (_32140_, _32139_, _07441_);
  nor (_32141_, _32140_, _32124_);
  and (_32143_, _32136_, _07441_);
  or (_32144_, _32143_, _05969_);
  nor (_32145_, _32144_, _32141_);
  or (_32146_, _32145_, _32121_);
  and (_32147_, _32146_, _03275_);
  nor (_32148_, _13139_, _11261_);
  nor (_32149_, _32148_, _32111_);
  nor (_32150_, _32149_, _03275_);
  or (_32151_, _32150_, _08861_);
  or (_32152_, _32151_, _32147_);
  and (_32154_, _13154_, _05343_);
  or (_32155_, _32111_, _04591_);
  or (_32156_, _32155_, _32154_);
  and (_32157_, _06358_, _05343_);
  nor (_32158_, _32157_, _32111_);
  and (_32159_, _32158_, _03650_);
  nor (_32160_, _32159_, _03778_);
  and (_32161_, _32160_, _32156_);
  and (_32162_, _32161_, _32152_);
  nor (_32163_, _32162_, _32117_);
  nor (_32165_, _32163_, _03655_);
  nor (_32166_, _32111_, _05601_);
  not (_32167_, _32166_);
  nor (_32168_, _32158_, _04596_);
  and (_32169_, _32168_, _32167_);
  nor (_32170_, _32169_, _32165_);
  nor (_32171_, _32170_, _03773_);
  nor (_32172_, _32123_, _04594_);
  and (_32173_, _32172_, _32167_);
  or (_32174_, _32173_, _32171_);
  and (_32176_, _32174_, _04608_);
  nor (_32177_, _13152_, _11261_);
  nor (_32178_, _32177_, _32111_);
  nor (_32179_, _32178_, _04608_);
  or (_32180_, _32179_, _32176_);
  and (_32181_, _32180_, _04606_);
  nor (_32182_, _32181_, _32114_);
  nor (_32183_, _32182_, _03809_);
  nor (_32184_, _32130_, _04260_);
  or (_32185_, _32184_, _03816_);
  nor (_32187_, _32185_, _32183_);
  and (_32188_, _13217_, _05343_);
  or (_32189_, _32111_, _03820_);
  nor (_32190_, _32189_, _32188_);
  nor (_32191_, _32190_, _32187_);
  or (_32192_, _32191_, _43231_);
  or (_32193_, _43227_, \oc8051_golden_model_1.TMOD [5]);
  and (_32194_, _32193_, _41991_);
  and (_43606_, _32194_, _32192_);
  not (_32195_, \oc8051_golden_model_1.TMOD [6]);
  nor (_32197_, _05343_, _32195_);
  nor (_32198_, _13373_, _11261_);
  nor (_32199_, _32198_, _32197_);
  nor (_32200_, _32199_, _04606_);
  and (_32201_, _13374_, _05343_);
  nor (_32202_, _32201_, _32197_);
  nor (_32203_, _32202_, _04589_);
  and (_32204_, _06531_, _05343_);
  or (_32205_, _32204_, _32197_);
  and (_32206_, _32205_, _05969_);
  and (_32208_, _05343_, \oc8051_golden_model_1.ACC [6]);
  nor (_32209_, _32208_, _32197_);
  nor (_32210_, _32209_, _04500_);
  nor (_32211_, _04499_, _32195_);
  or (_32212_, _32211_, _32210_);
  and (_32213_, _32212_, _04515_);
  nor (_32214_, _13235_, _11261_);
  nor (_32215_, _32214_, _32197_);
  nor (_32216_, _32215_, _04515_);
  or (_32217_, _32216_, _32213_);
  and (_32219_, _32217_, _04524_);
  nor (_32220_, _05442_, _11261_);
  nor (_32221_, _32220_, _32197_);
  nor (_32222_, _32221_, _04524_);
  nor (_32223_, _32222_, _32219_);
  nor (_32224_, _32223_, _03603_);
  nor (_32225_, _32209_, _03611_);
  nor (_32226_, _32225_, _07441_);
  not (_32227_, _32226_);
  nor (_32228_, _32227_, _32224_);
  and (_32230_, _32221_, _07441_);
  or (_32231_, _32230_, _05969_);
  nor (_32232_, _32231_, _32228_);
  or (_32233_, _32232_, _32206_);
  and (_32234_, _32233_, _03275_);
  nor (_32235_, _13356_, _11261_);
  nor (_32236_, _32235_, _32197_);
  nor (_32237_, _32236_, _03275_);
  or (_32238_, _32237_, _08861_);
  or (_32239_, _32238_, _32234_);
  and (_32241_, _13245_, _05343_);
  or (_32242_, _32197_, _04591_);
  or (_32243_, _32242_, _32241_);
  and (_32244_, _13363_, _05343_);
  nor (_32245_, _32244_, _32197_);
  and (_32246_, _32245_, _03650_);
  nor (_32247_, _32246_, _03778_);
  and (_32248_, _32247_, _32243_);
  and (_32249_, _32248_, _32239_);
  nor (_32250_, _32249_, _32203_);
  nor (_32252_, _32250_, _03655_);
  nor (_32253_, _32197_, _05491_);
  not (_32254_, _32253_);
  nor (_32255_, _32245_, _04596_);
  and (_32256_, _32255_, _32254_);
  nor (_32257_, _32256_, _32252_);
  nor (_32258_, _32257_, _03773_);
  nor (_32259_, _32209_, _04594_);
  and (_32260_, _32259_, _32254_);
  or (_32261_, _32260_, _32258_);
  and (_32262_, _32261_, _04608_);
  nor (_32263_, _13243_, _11261_);
  nor (_32264_, _32263_, _32197_);
  nor (_32265_, _32264_, _04608_);
  or (_32266_, _32265_, _32262_);
  and (_32267_, _32266_, _04606_);
  nor (_32268_, _32267_, _32200_);
  nor (_32269_, _32268_, _03809_);
  nor (_32270_, _32215_, _04260_);
  or (_32271_, _32270_, _03816_);
  nor (_32273_, _32271_, _32269_);
  and (_32274_, _13425_, _05343_);
  or (_32275_, _32197_, _03820_);
  nor (_32276_, _32275_, _32274_);
  nor (_32277_, _32276_, _32273_);
  or (_32278_, _32277_, _43231_);
  or (_32279_, _43227_, \oc8051_golden_model_1.TMOD [6]);
  and (_32280_, _32279_, _41991_);
  and (_43607_, _32280_, _32278_);
  and (_32281_, _11984_, _04172_);
  and (_32283_, _11967_, _11974_);
  nor (_32284_, _32283_, _02938_);
  and (_32285_, _11945_, _11952_);
  nor (_32286_, _32285_, _02938_);
  not (_32287_, _03246_);
  and (_32288_, _11353_, _08770_);
  nor (_32289_, _32288_, _02938_);
  and (_32290_, _08375_, \oc8051_golden_model_1.PC [0]);
  nor (_32291_, _08375_, \oc8051_golden_model_1.PC [0]);
  or (_32292_, _32291_, _32290_);
  or (_32294_, _32292_, _11894_);
  not (_32295_, _03236_);
  and (_32296_, _11361_, _04608_);
  nor (_32297_, _32296_, _02938_);
  not (_32298_, _03238_);
  and (_32299_, _11370_, _04596_);
  nor (_32300_, _32299_, _02938_);
  not (_32301_, _03231_);
  and (_32302_, _11841_, _04591_);
  nor (_32303_, _32302_, _02938_);
  and (_32304_, _03650_, _02938_);
  nor (_32305_, _04172_, _03265_);
  nor (_32306_, _04172_, _03260_);
  nor (_32307_, _11540_, _02938_);
  not (_32308_, _04063_);
  and (_32309_, _11531_, _32308_);
  nor (_32310_, _32309_, _02938_);
  and (_32311_, _32309_, _02938_);
  nor (_32312_, _32311_, _32310_);
  nand (_32313_, _32312_, _04868_);
  or (_32316_, _04172_, _04868_);
  and (_32317_, _32316_, _11540_);
  and (_32318_, _32317_, _32313_);
  nor (_32319_, _32318_, _32307_);
  nor (_32320_, _32319_, _12226_);
  and (_32321_, _11554_, \oc8051_golden_model_1.PC [0]);
  and (_32322_, _04042_, _02938_);
  nor (_32323_, _32322_, _11618_);
  and (_32324_, _32323_, _11556_);
  or (_32325_, _32324_, _32321_);
  nor (_32327_, _32325_, _06054_);
  nor (_32328_, _32327_, _32320_);
  nor (_32329_, _32328_, _04509_);
  and (_32330_, _04509_, \oc8051_golden_model_1.PC [0]);
  nor (_32331_, _32330_, _32329_);
  and (_32332_, _32331_, _04515_);
  and (_32333_, _11397_, \oc8051_golden_model_1.PC [0]);
  not (_32334_, _32333_);
  and (_32335_, _04172_, \oc8051_golden_model_1.PC [0]);
  nor (_32336_, _32335_, _11472_);
  not (_32338_, _32336_);
  and (_32339_, _32338_, _11526_);
  nor (_32340_, _32339_, _04515_);
  and (_32341_, _32340_, _32334_);
  nor (_32342_, _32341_, _11392_);
  not (_32343_, _32342_);
  nor (_32344_, _32343_, _32332_);
  nor (_32345_, _11391_, _02938_);
  nor (_32346_, _32345_, _04857_);
  not (_32347_, _32346_);
  nor (_32349_, _32347_, _32344_);
  nor (_32350_, _04172_, _03257_);
  and (_32351_, _11692_, _11684_);
  not (_32352_, _32351_);
  nor (_32353_, _32352_, _32350_);
  not (_32354_, _32353_);
  nor (_32355_, _32354_, _32349_);
  nor (_32356_, _32351_, _02938_);
  nor (_32357_, _32356_, _11696_);
  not (_32358_, _32357_);
  nor (_32360_, _32358_, _32355_);
  or (_32361_, _32360_, _11706_);
  nor (_32362_, _32361_, _32306_);
  and (_32363_, _10037_, _02938_);
  nor (_32364_, _32338_, _10037_);
  or (_32365_, _32364_, _09988_);
  nor (_32366_, _32365_, _32363_);
  or (_32367_, _32366_, _10041_);
  nor (_32368_, _32367_, _32362_);
  or (_32369_, _32336_, _10089_);
  nand (_32371_, _10089_, \oc8051_golden_model_1.PC [0]);
  and (_32372_, _32371_, _10041_);
  and (_32373_, _32372_, _32369_);
  or (_32374_, _32373_, _32368_);
  and (_32375_, _32374_, _04046_);
  and (_32376_, _09946_, _02938_);
  nor (_32377_, _32338_, _09946_);
  nor (_32378_, _32377_, _32376_);
  nor (_32379_, _32378_, _04046_);
  nor (_32380_, _32379_, _32375_);
  nor (_32382_, _32380_, _03676_);
  and (_32383_, _10133_, _02938_);
  nor (_32384_, _32338_, _10133_);
  or (_32385_, _32384_, _32383_);
  and (_32386_, _32385_, _03676_);
  or (_32387_, _32386_, _32382_);
  and (_32388_, _32387_, _11389_);
  and (_32389_, _10096_, _02938_);
  or (_32390_, _32389_, _32388_);
  and (_32391_, _32390_, _03253_);
  nor (_32393_, _04172_, _03253_);
  nor (_32394_, _32393_, _11387_);
  not (_32395_, _32394_);
  nor (_32396_, _32395_, _32391_);
  not (_32397_, _03265_);
  nor (_32398_, _11386_, _02938_);
  nor (_32399_, _32398_, _32397_);
  not (_32400_, _32399_);
  nor (_32401_, _32400_, _32396_);
  and (_32402_, _11381_, _03285_);
  not (_32404_, _32402_);
  or (_32405_, _32404_, _32401_);
  nor (_32406_, _32405_, _32305_);
  nor (_32407_, _32402_, _02938_);
  nor (_32408_, _32407_, _03497_);
  not (_32409_, _32408_);
  nor (_32410_, _32409_, _32406_);
  nor (_32411_, _04172_, _03278_);
  nor (_32412_, _03656_, _03644_);
  and (_32413_, _32412_, _11767_);
  not (_32415_, _32413_);
  nor (_32416_, _32415_, _32411_);
  not (_32417_, _32416_);
  nor (_32418_, _32417_, _32410_);
  nor (_32419_, _32413_, _02938_);
  nor (_32420_, _32419_, _03220_);
  not (_32421_, _32420_);
  nor (_32422_, _32421_, _32418_);
  nor (_32423_, _04172_, _03221_);
  or (_32424_, _32423_, _11372_);
  or (_32426_, _32424_, _32422_);
  or (_32427_, _32323_, _11373_);
  and (_32428_, _32427_, _32426_);
  and (_32429_, _32428_, _04582_);
  or (_32430_, _32429_, _32304_);
  and (_32431_, _32430_, _11785_);
  and (_32432_, _11784_, _03388_);
  or (_32433_, _32432_, _32431_);
  and (_32434_, _32433_, _27673_);
  nor (_32435_, _04172_, _27673_);
  or (_32437_, _32435_, _32434_);
  and (_32438_, _32437_, _11827_);
  not (_32439_, _32302_);
  and (_32440_, _08820_, \oc8051_golden_model_1.PC [0]);
  and (_32441_, _32323_, _11832_);
  or (_32442_, _32441_, _32440_);
  and (_32443_, _32442_, _11826_);
  nor (_32444_, _32443_, _32439_);
  not (_32445_, _32444_);
  nor (_32446_, _32445_, _32438_);
  nor (_32448_, _32446_, _32303_);
  and (_32449_, _32448_, _32301_);
  nor (_32450_, _04172_, _32301_);
  or (_32451_, _32450_, _32449_);
  and (_32452_, _32451_, _11857_);
  not (_32453_, _32299_);
  nor (_32454_, _32323_, _11832_);
  nor (_32455_, _08820_, \oc8051_golden_model_1.PC [0]);
  nor (_32456_, _32455_, _11857_);
  not (_32457_, _32456_);
  nor (_32459_, _32457_, _32454_);
  nor (_32460_, _32459_, _32453_);
  not (_32461_, _32460_);
  nor (_32462_, _32461_, _32452_);
  nor (_32463_, _32462_, _32300_);
  and (_32464_, _32463_, _32298_);
  nor (_32465_, _04172_, _32298_);
  or (_32466_, _32465_, _32464_);
  and (_32467_, _32466_, _11364_);
  not (_32468_, _32296_);
  and (_32470_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and (_32471_, _32323_, _07911_);
  or (_32472_, _32471_, _32470_);
  and (_32473_, _32472_, _11363_);
  nor (_32474_, _32473_, _32468_);
  not (_32475_, _32474_);
  nor (_32476_, _32475_, _32467_);
  nor (_32477_, _32476_, _32297_);
  and (_32478_, _32477_, _32295_);
  nor (_32479_, _04172_, _32295_);
  or (_32481_, _32479_, _32478_);
  and (_32482_, _32481_, _11894_);
  and (_32483_, _11355_, _08601_);
  not (_32484_, _32483_);
  nor (_32485_, _32484_, _32482_);
  and (_32486_, _32485_, _32294_);
  nor (_32487_, _32483_, _02938_);
  nor (_32488_, _32487_, _03792_);
  not (_32489_, _32488_);
  nor (_32490_, _32489_, _32486_);
  and (_32492_, _06836_, _03792_);
  or (_32493_, _32492_, _32490_);
  and (_32494_, _32493_, _06475_);
  nor (_32495_, _04172_, _06475_);
  or (_32496_, _32495_, _32494_);
  and (_32497_, _32496_, _03796_);
  and (_32498_, _32338_, _09914_);
  nor (_32499_, _09914_, _02938_);
  or (_32500_, _32499_, _03796_);
  or (_32501_, _32500_, _32498_);
  and (_32503_, _32501_, _32288_);
  not (_32504_, _32503_);
  nor (_32505_, _32504_, _32497_);
  nor (_32506_, _32505_, _32289_);
  and (_32507_, _32506_, _03522_);
  and (_32508_, _06836_, _03521_);
  or (_32509_, _32508_, _32507_);
  and (_32510_, _32509_, _32287_);
  nor (_32511_, _04172_, _32287_);
  nor (_32512_, _32511_, _32510_);
  nor (_32514_, _32512_, _03519_);
  not (_32515_, _32285_);
  and (_32516_, _09914_, \oc8051_golden_model_1.PC [0]);
  nor (_32517_, _32336_, _09914_);
  nor (_32518_, _32517_, _32516_);
  and (_32519_, _32518_, _03519_);
  nor (_32520_, _32519_, _32515_);
  not (_32521_, _32520_);
  nor (_32522_, _32521_, _32514_);
  nor (_32523_, _32522_, _32286_);
  nor (_32525_, _32523_, _05047_);
  and (_32526_, _05047_, _04172_);
  nor (_32527_, _32526_, _03205_);
  not (_32528_, _32527_);
  nor (_32529_, _32528_, _32525_);
  not (_32530_, _32283_);
  and (_32531_, _32518_, _03205_);
  nor (_32532_, _32531_, _32530_);
  not (_32533_, _32532_);
  nor (_32534_, _32533_, _32529_);
  nor (_32536_, _32534_, _32284_);
  nor (_32537_, _32536_, _11984_);
  or (_32538_, _32537_, _11982_);
  nor (_32539_, _32538_, _32281_);
  and (_32540_, _11982_, _02938_);
  nor (_32541_, _32540_, _32539_);
  nand (_32542_, _32541_, _43227_);
  or (_32543_, _43227_, \oc8051_golden_model_1.PC [0]);
  and (_32544_, _32543_, _41991_);
  and (_43608_, _32544_, _32542_);
  and (_32546_, _03816_, _02911_);
  and (_32547_, _03809_, _02911_);
  or (_32548_, _11353_, _11470_);
  nor (_32549_, _06886_, _04220_);
  nand (_32550_, _32549_, _03321_);
  or (_32551_, _11361_, _11470_);
  and (_32552_, _04563_, _03237_);
  nand (_32553_, _32552_, _03321_);
  or (_32554_, _11841_, _11470_);
  or (_32555_, _11381_, _11470_);
  nand (_32557_, _10096_, _03321_);
  nor (_32558_, _03681_, _03678_);
  not (_32559_, _32558_);
  nor (_32560_, _11474_, _11472_);
  nor (_32561_, _32560_, _11475_);
  or (_32562_, _32561_, _10037_);
  nand (_32563_, _10037_, _11470_);
  and (_32564_, _32563_, _32562_);
  or (_32565_, _32564_, _09988_);
  or (_32566_, _11692_, _11470_);
  and (_32568_, _04509_, _11470_);
  nor (_32569_, _11620_, _11618_);
  nor (_32570_, _32569_, _11621_);
  and (_32571_, _32570_, _11556_);
  and (_32572_, _11554_, _02911_);
  or (_32573_, _32572_, _32571_);
  or (_32574_, _32573_, _06054_);
  or (_32575_, _11540_, _11470_);
  nor (_32576_, _04347_, _04868_);
  not (_32577_, _11540_);
  nand (_32579_, _04063_, _03321_);
  nor (_32580_, _11531_, _02938_);
  nor (_32581_, _32580_, _04499_);
  and (_32582_, _32581_, \oc8051_golden_model_1.PC [1]);
  nor (_32583_, _32581_, \oc8051_golden_model_1.PC [1]);
  or (_32584_, _32583_, _32582_);
  or (_32585_, _32584_, _04063_);
  and (_32586_, _32585_, _32579_);
  and (_32587_, _32586_, _04868_);
  or (_32588_, _32587_, _32577_);
  or (_32590_, _32588_, _32576_);
  and (_32591_, _32590_, _32575_);
  or (_32592_, _32591_, _12226_);
  and (_32593_, _32592_, _06068_);
  and (_32594_, _32593_, _32574_);
  or (_32595_, _32594_, _32568_);
  and (_32596_, _32595_, _04515_);
  and (_32597_, _11397_, _03321_);
  and (_32598_, _32561_, _11526_);
  or (_32599_, _32598_, _32597_);
  and (_32601_, _32599_, _03599_);
  or (_32602_, _32601_, _11392_);
  or (_32603_, _32602_, _32596_);
  or (_32604_, _11391_, _11470_);
  and (_32605_, _32604_, _03516_);
  and (_32606_, _32605_, _32603_);
  and (_32607_, _03515_, _02911_);
  or (_32608_, _32607_, _04857_);
  or (_32609_, _32608_, _32606_);
  nand (_32610_, _04347_, _04857_);
  and (_32611_, _32610_, _04524_);
  and (_32612_, _32611_, _32609_);
  nand (_32613_, _03597_, _02911_);
  nand (_32614_, _32613_, _11684_);
  or (_32615_, _32614_, _32612_);
  or (_32616_, _11684_, _11470_);
  and (_32617_, _32616_, _03611_);
  and (_32618_, _32617_, _32615_);
  nand (_32619_, _03603_, _02911_);
  nand (_32620_, _32619_, _11692_);
  or (_32623_, _32620_, _32618_);
  and (_32624_, _32623_, _32566_);
  or (_32625_, _32624_, _03511_);
  nand (_32626_, _03511_, \oc8051_golden_model_1.PC [1]);
  and (_32627_, _32626_, _03260_);
  and (_32628_, _32627_, _32625_);
  nor (_32629_, _04347_, _03260_);
  or (_32630_, _32629_, _32628_);
  and (_32631_, _32630_, _04650_);
  nand (_32632_, _03510_, _02911_);
  nand (_32634_, _32632_, _09988_);
  or (_32635_, _32634_, _32631_);
  and (_32636_, _32635_, _32565_);
  or (_32637_, _32636_, _32559_);
  and (_32638_, _10089_, _03321_);
  and (_32639_, _32561_, _11713_);
  or (_32640_, _32639_, _32558_);
  or (_32641_, _32640_, _32638_);
  and (_32642_, _32641_, _04046_);
  and (_32643_, _32642_, _32637_);
  and (_32645_, _32561_, _11719_);
  and (_32646_, _09946_, _03321_);
  or (_32647_, _32646_, _32645_);
  and (_32648_, _32647_, _03615_);
  or (_32649_, _32648_, _32643_);
  and (_32650_, _32649_, _09916_);
  nand (_32651_, _10133_, _11470_);
  or (_32652_, _32561_, _10133_);
  and (_32653_, _32652_, _03676_);
  and (_32654_, _32653_, _32651_);
  or (_32656_, _32654_, _10096_);
  or (_32657_, _32656_, _32650_);
  and (_32658_, _32657_, _32557_);
  or (_32659_, _32658_, _03504_);
  nand (_32660_, _03504_, \oc8051_golden_model_1.PC [1]);
  and (_32661_, _32660_, _03253_);
  and (_32662_, _32661_, _32659_);
  nor (_32663_, _04347_, _03253_);
  not (_32664_, _05073_);
  and (_32665_, _23569_, _32664_);
  and (_32667_, _32665_, _23572_);
  not (_32668_, _32667_);
  or (_32669_, _32668_, _32663_);
  or (_32670_, _32669_, _32662_);
  or (_32671_, _32667_, _02911_);
  and (_32672_, _32671_, _11384_);
  and (_32673_, _32672_, _32670_);
  nand (_32674_, _11383_, _11470_);
  nand (_32675_, _32674_, _11385_);
  or (_32676_, _32675_, _32673_);
  or (_32678_, _11385_, _11470_);
  and (_32679_, _32678_, _09729_);
  and (_32680_, _32679_, _32676_);
  and (_32681_, _03630_, _02911_);
  or (_32682_, _32681_, _32397_);
  or (_32683_, _32682_, _32680_);
  nand (_32684_, _04347_, _32397_);
  and (_32685_, _32684_, _09728_);
  and (_32686_, _32685_, _32683_);
  nand (_32687_, _03629_, _02911_);
  nand (_32689_, _32687_, _11381_);
  or (_32690_, _32689_, _32686_);
  and (_32691_, _32690_, _32555_);
  or (_32692_, _32691_, _11380_);
  or (_32693_, _11379_, _02911_);
  and (_32694_, _32693_, _03285_);
  and (_32695_, _32694_, _32692_);
  nor (_32696_, _03321_, _03285_);
  or (_32697_, _32696_, _03500_);
  or (_32698_, _32697_, _32695_);
  nand (_32700_, _03500_, \oc8051_golden_model_1.PC [1]);
  and (_32701_, _32700_, _32698_);
  or (_32702_, _32701_, _03497_);
  nand (_32703_, _04347_, _03497_);
  and (_32704_, _32703_, _08865_);
  and (_32705_, _32704_, _32702_);
  nand (_32706_, _03656_, _03321_);
  nand (_32707_, _32706_, _11759_);
  or (_32708_, _32707_, _32705_);
  or (_32709_, _11759_, _02911_);
  and (_32711_, _32709_, _03275_);
  and (_32712_, _32711_, _32708_);
  or (_32713_, _11470_, _03275_);
  nand (_32714_, _32713_, _11767_);
  or (_32715_, _32714_, _32712_);
  not (_32716_, _03562_);
  or (_32717_, _11767_, _11470_);
  and (_32718_, _32717_, _32716_);
  and (_32719_, _32718_, _32715_);
  and (_32720_, _03562_, _02911_);
  or (_32722_, _32720_, _03220_);
  or (_32723_, _32722_, _32719_);
  nand (_32724_, _04347_, _03220_);
  and (_32725_, _32724_, _11373_);
  and (_32726_, _32725_, _32723_);
  and (_32727_, _32570_, _11372_);
  or (_32728_, _32727_, _06246_);
  or (_32729_, _32728_, _32726_);
  nor (_32730_, _03650_, \oc8051_golden_model_1.PC [1]);
  or (_32731_, _32730_, _05967_);
  and (_32733_, _32731_, _32729_);
  and (_32734_, _03650_, _03321_);
  or (_32735_, _32734_, _08445_);
  or (_32736_, _32735_, _32733_);
  nand (_32737_, _08445_, \oc8051_golden_model_1.PC [1]);
  and (_32738_, _32737_, _32736_);
  or (_32739_, _32738_, _11784_);
  or (_32740_, _11785_, _03373_);
  and (_32741_, _32740_, _04181_);
  and (_32742_, _32741_, _32739_);
  and (_32744_, _03561_, _02911_);
  or (_32745_, _32744_, _03227_);
  or (_32746_, _32745_, _32742_);
  nand (_32747_, _04347_, _03227_);
  and (_32748_, _32747_, _11827_);
  and (_32749_, _32748_, _32746_);
  or (_32750_, _32570_, _08820_);
  nand (_32751_, _08820_, \oc8051_golden_model_1.PC [1]);
  and (_32752_, _32751_, _11826_);
  and (_32753_, _32752_, _32750_);
  or (_32755_, _32753_, _11845_);
  or (_32756_, _32755_, _32749_);
  and (_32757_, _32756_, _32554_);
  or (_32758_, _32757_, _11844_);
  or (_32759_, _11843_, _02911_);
  and (_32760_, _32759_, _04591_);
  and (_32761_, _32760_, _32758_);
  and (_32762_, _03649_, _03321_);
  or (_32763_, _32762_, _03778_);
  or (_32764_, _32763_, _32761_);
  nand (_32766_, _03778_, \oc8051_golden_model_1.PC [1]);
  and (_32767_, _32766_, _32764_);
  or (_32768_, _32767_, _03231_);
  nand (_32769_, _04347_, _03231_);
  and (_32770_, _32769_, _11857_);
  and (_32771_, _32770_, _32768_);
  or (_32772_, _32570_, _11832_);
  or (_32773_, _08820_, _02911_);
  and (_32774_, _32773_, _11856_);
  and (_32775_, _32774_, _32772_);
  or (_32777_, _32775_, _32552_);
  or (_32778_, _32777_, _32771_);
  and (_32779_, _32778_, _32553_);
  and (_32780_, _04839_, _08044_);
  nor (_32781_, _32780_, _04194_);
  or (_32782_, _32781_, _32779_);
  and (_32783_, _32781_, _03321_);
  nor (_32784_, _32783_, _04199_);
  and (_32785_, _32784_, _32782_);
  nand (_32786_, _04199_, _11470_);
  nand (_32788_, _32786_, _11367_);
  or (_32789_, _32788_, _32785_);
  or (_32790_, _11367_, _02911_);
  and (_32791_, _32790_, _04596_);
  and (_32792_, _32791_, _32789_);
  and (_32793_, _03655_, _03321_);
  or (_32794_, _32793_, _03773_);
  or (_32795_, _32794_, _32792_);
  nand (_32796_, _03773_, \oc8051_golden_model_1.PC [1]);
  and (_32797_, _32796_, _32795_);
  or (_32799_, _32797_, _03238_);
  nand (_32800_, _04347_, _03238_);
  and (_32801_, _32800_, _11364_);
  and (_32802_, _32801_, _32799_);
  or (_32803_, _32570_, \oc8051_golden_model_1.PSW [7]);
  nand (_32804_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_32805_, _32804_, _11363_);
  and (_32806_, _32805_, _32803_);
  or (_32807_, _32806_, _11877_);
  or (_32808_, _32807_, _32802_);
  and (_32810_, _32808_, _32551_);
  or (_32811_, _32810_, _11358_);
  or (_32812_, _11357_, _02911_);
  and (_32813_, _32812_, _04608_);
  and (_32814_, _32813_, _32811_);
  and (_32815_, _03653_, _03321_);
  or (_32816_, _32815_, _03786_);
  or (_32817_, _32816_, _32814_);
  nand (_32818_, _03786_, \oc8051_golden_model_1.PC [1]);
  and (_32819_, _32818_, _32817_);
  or (_32821_, _32819_, _03236_);
  nand (_32822_, _04347_, _03236_);
  and (_32823_, _32822_, _11894_);
  and (_32824_, _32823_, _32821_);
  or (_32825_, _32570_, _07911_);
  or (_32826_, \oc8051_golden_model_1.PSW [7], _02911_);
  and (_32827_, _32826_, _11893_);
  and (_32828_, _32827_, _32825_);
  or (_32829_, _32828_, _32549_);
  or (_32830_, _32829_, _32824_);
  and (_32832_, _32830_, _32550_);
  and (_32833_, _03567_, _03283_);
  or (_32834_, _32833_, _03680_);
  and (_32835_, _32834_, _03247_);
  or (_32836_, _32835_, _32832_);
  and (_32837_, _32835_, _03321_);
  nor (_32838_, _32837_, _04217_);
  and (_32839_, _32838_, _32836_);
  nand (_32840_, _04217_, _11470_);
  nand (_32841_, _32840_, _08570_);
  or (_32843_, _32841_, _32839_);
  or (_32844_, _08570_, _02911_);
  and (_32845_, _32844_, _08601_);
  and (_32846_, _32845_, _32843_);
  and (_32847_, _08600_, _11470_);
  or (_32848_, _32847_, _03792_);
  or (_32849_, _32848_, _32846_);
  or (_32850_, _06835_, _10680_);
  and (_32851_, _32850_, _32849_);
  or (_32852_, _32851_, _03248_);
  nand (_32854_, _04347_, _03248_);
  and (_32855_, _32854_, _03796_);
  and (_32856_, _32855_, _32852_);
  or (_32857_, _32561_, _11920_);
  or (_32858_, _09914_, _03321_);
  and (_32859_, _32858_, _03652_);
  and (_32860_, _32859_, _32857_);
  or (_32861_, _32860_, _11919_);
  or (_32862_, _32861_, _32856_);
  and (_32863_, _32862_, _32548_);
  or (_32865_, _32863_, _08722_);
  or (_32866_, _08721_, _02911_);
  and (_32867_, _32866_, _08770_);
  and (_32868_, _32867_, _32865_);
  and (_32869_, _08769_, _11470_);
  or (_32870_, _32869_, _03521_);
  or (_32871_, _32870_, _32868_);
  or (_32872_, _06835_, _03522_);
  and (_32873_, _32872_, _32871_);
  or (_32874_, _32873_, _03246_);
  nand (_32876_, _04347_, _03246_);
  and (_32877_, _32876_, _03520_);
  and (_32878_, _32877_, _32874_);
  or (_32879_, _32561_, _09914_);
  nand (_32880_, _09914_, _11470_);
  and (_32881_, _32880_, _32879_);
  and (_32882_, _32881_, _03519_);
  or (_32883_, _32882_, _06481_);
  or (_32884_, _32883_, _32878_);
  nand (_32885_, _06481_, _03321_);
  and (_32887_, _32885_, _32884_);
  or (_32888_, _32887_, _04827_);
  nand (_32889_, _04827_, _03321_);
  and (_32890_, _32889_, _04260_);
  and (_32891_, _32890_, _32888_);
  or (_32892_, _32891_, _32547_);
  and (_32893_, _32892_, _11952_);
  nor (_32894_, _11952_, _03321_);
  or (_32895_, _32894_, _05047_);
  or (_32896_, _32895_, _32893_);
  nand (_32898_, _05047_, _04347_);
  and (_32899_, _32898_, _03206_);
  and (_32900_, _32899_, _32896_);
  or (_32901_, _06886_, _04838_);
  nand (_32902_, _32881_, _03205_);
  nand (_32903_, _32902_, _32901_);
  or (_32904_, _32903_, _32900_);
  nor (_32905_, _04642_, _04266_);
  or (_32906_, _32901_, _11470_);
  and (_32907_, _32906_, _32905_);
  and (_32909_, _32907_, _32904_);
  nor (_32910_, _32905_, _03321_);
  or (_32911_, _32910_, _04271_);
  or (_32912_, _32911_, _32909_);
  and (_32913_, _04271_, _03321_);
  nor (_32914_, _32913_, _03816_);
  and (_32915_, _32914_, _32912_);
  or (_32916_, _32915_, _32546_);
  and (_32917_, _32916_, _11974_);
  nor (_32918_, _11974_, _03321_);
  or (_32920_, _32918_, _11984_);
  or (_32921_, _32920_, _32917_);
  nand (_32922_, _11984_, _04347_);
  and (_32923_, _32922_, _11990_);
  and (_32924_, _32923_, _32921_);
  and (_32925_, _11982_, _11470_);
  or (_32926_, _32925_, _32924_);
  or (_32927_, _32926_, _43231_);
  or (_32928_, _43227_, \oc8051_golden_model_1.PC [1]);
  and (_32929_, _32928_, _41991_);
  and (_43611_, _32929_, _32927_);
  and (_32931_, _03816_, _03356_);
  and (_32932_, _03809_, _03356_);
  nor (_32933_, _11353_, _03318_);
  nor (_32934_, _11355_, _03318_);
  nor (_32935_, _11361_, _03318_);
  nor (_32936_, _11370_, _03318_);
  nor (_32937_, _11841_, _03318_);
  and (_32938_, _03500_, _03362_);
  nor (_32939_, _11381_, _03318_);
  nor (_32941_, _32667_, _03356_);
  not (_32942_, _03318_);
  and (_32943_, _10096_, _32942_);
  and (_32944_, _11467_, _09946_);
  and (_32945_, _11479_, _11476_);
  nor (_32946_, _32945_, _11480_);
  not (_32947_, _32946_);
  nor (_32948_, _32947_, _09946_);
  nor (_32949_, _32948_, _32944_);
  or (_32950_, _32949_, _04046_);
  and (_32952_, _11467_, _10089_);
  nor (_32953_, _32947_, _10089_);
  nor (_32954_, _32953_, _32952_);
  nand (_32955_, _32954_, _10041_);
  or (_32956_, _32947_, _11397_);
  or (_32957_, _11468_, _11526_);
  and (_32958_, _32957_, _03599_);
  and (_32959_, _32958_, _32956_);
  and (_32960_, _11554_, _03362_);
  and (_32961_, _11625_, _11622_);
  nor (_32962_, _32961_, _11626_);
  not (_32963_, _32962_);
  and (_32964_, _32963_, _11556_);
  or (_32965_, _32964_, _06054_);
  or (_32966_, _32965_, _32960_);
  and (_32967_, _03947_, _03943_);
  nand (_32968_, _03946_, _03362_);
  and (_32969_, _11531_, \oc8051_golden_model_1.PC [2]);
  or (_32970_, _32969_, _04499_);
  and (_32971_, _32970_, _11537_);
  nor (_32974_, _11531_, _32942_);
  or (_32975_, _32974_, _32971_);
  and (_32976_, _32975_, _32968_);
  and (_32977_, _11540_, _04868_);
  nand (_32978_, _11536_, _03318_);
  nand (_32979_, _32978_, _32977_);
  nor (_32980_, _32979_, _32976_);
  nor (_32981_, _11540_, _03318_);
  or (_32982_, _32981_, _12226_);
  or (_32983_, _32982_, _32980_);
  or (_32985_, _32983_, _32967_);
  and (_32986_, _32985_, _32966_);
  or (_32987_, _32986_, _04509_);
  nand (_32988_, _04509_, _03318_);
  and (_32989_, _32988_, _04515_);
  and (_32990_, _32989_, _32987_);
  or (_32991_, _32990_, _32959_);
  nand (_32992_, _32991_, _11391_);
  nor (_32993_, _11391_, _03318_);
  nor (_32994_, _32993_, _03515_);
  nand (_32996_, _32994_, _32992_);
  and (_32997_, _03515_, _03356_);
  nor (_32998_, _32997_, _04857_);
  nand (_32999_, _32998_, _32996_);
  and (_33000_, _03943_, _04857_);
  nor (_33001_, _33000_, _03597_);
  nand (_33002_, _33001_, _32999_);
  not (_33003_, _11684_);
  and (_33004_, _03597_, _03356_);
  nor (_33005_, _33004_, _33003_);
  nand (_33007_, _33005_, _33002_);
  nor (_33008_, _11684_, _03318_);
  nor (_33009_, _33008_, _03603_);
  nand (_33010_, _33009_, _33007_);
  and (_33011_, _03603_, _03356_);
  nor (_33012_, _33011_, _11694_);
  nand (_33013_, _33012_, _33010_);
  nor (_33014_, _11692_, _03318_);
  nor (_33015_, _33014_, _03511_);
  nand (_33016_, _33015_, _33013_);
  and (_33017_, _03511_, _03356_);
  nor (_33018_, _33017_, _11696_);
  nand (_33019_, _33018_, _33016_);
  and (_33020_, _03943_, _11696_);
  nor (_33021_, _33020_, _03510_);
  nand (_33022_, _33021_, _33019_);
  and (_33023_, _03510_, _03356_);
  nor (_33024_, _33023_, _11706_);
  and (_33025_, _33024_, _33022_);
  and (_33026_, _11467_, _10037_);
  nor (_33028_, _32947_, _10037_);
  or (_33029_, _33028_, _33026_);
  nor (_33030_, _33029_, _09988_);
  or (_33031_, _33030_, _33025_);
  nand (_33032_, _33031_, _10042_);
  nand (_33033_, _33032_, _32955_);
  or (_33034_, _33033_, _03615_);
  and (_33035_, _33034_, _32950_);
  or (_33036_, _33035_, _03676_);
  nand (_33037_, _11468_, _10133_);
  or (_33039_, _32946_, _10133_);
  and (_33040_, _33039_, _03676_);
  and (_33041_, _33040_, _33037_);
  nor (_33042_, _33041_, _10096_);
  and (_33043_, _33042_, _33036_);
  or (_33044_, _33043_, _32943_);
  nand (_33045_, _33044_, _03505_);
  and (_33046_, _03504_, _03362_);
  nor (_33047_, _33046_, _04998_);
  nand (_33048_, _33047_, _33045_);
  nor (_33050_, _03943_, _03253_);
  nor (_33051_, _33050_, _32668_);
  and (_33052_, _33051_, _33048_);
  or (_33053_, _33052_, _32941_);
  nand (_33054_, _33053_, _11386_);
  nor (_33055_, _11386_, _03318_);
  nor (_33056_, _33055_, _03630_);
  nand (_33057_, _33056_, _33054_);
  and (_33058_, _03630_, _03356_);
  nor (_33059_, _33058_, _32397_);
  nand (_33061_, _33059_, _33057_);
  and (_33062_, _03943_, _32397_);
  nor (_33063_, _33062_, _03629_);
  nand (_33064_, _33063_, _33061_);
  not (_33065_, _11381_);
  and (_33066_, _03629_, _03356_);
  nor (_33067_, _33066_, _33065_);
  and (_33068_, _33067_, _33064_);
  or (_33069_, _33068_, _32939_);
  nand (_33070_, _33069_, _11379_);
  nor (_33072_, _11379_, _03356_);
  nor (_33073_, _33072_, _03371_);
  nand (_33074_, _33073_, _33070_);
  nor (_33075_, _32942_, _03285_);
  nor (_33076_, _33075_, _03500_);
  and (_33077_, _33076_, _33074_);
  or (_33078_, _33077_, _32938_);
  nand (_33079_, _33078_, _03278_);
  and (_33080_, _03943_, _03497_);
  nor (_33081_, _33080_, _03656_);
  nand (_33083_, _33081_, _33079_);
  and (_33084_, _11467_, _03656_);
  not (_33085_, _33084_);
  and (_33086_, _33085_, _11759_);
  nand (_33087_, _33086_, _33083_);
  nor (_33088_, _11759_, _03356_);
  nor (_33089_, _33088_, _03644_);
  nand (_33090_, _33089_, _33087_);
  nor (_33091_, _11468_, _03275_);
  nor (_33092_, _33091_, _11770_);
  nand (_33094_, _33092_, _33090_);
  nor (_33095_, _11767_, _03318_);
  nor (_33096_, _33095_, _03562_);
  and (_33097_, _33096_, _33094_);
  and (_33098_, _03562_, _03356_);
  or (_33099_, _33098_, _03220_);
  nor (_33100_, _33099_, _33097_);
  and (_33101_, _03943_, _03220_);
  or (_33102_, _33101_, _33100_);
  nand (_33103_, _33102_, _11373_);
  nor (_33105_, _32962_, _11373_);
  not (_33106_, _04844_);
  and (_33107_, _03584_, _03226_);
  nor (_33108_, _33107_, _04849_);
  and (_33109_, _33108_, _33106_);
  not (_33110_, _33109_);
  nor (_33111_, _33110_, _33105_);
  nand (_33112_, _33111_, _33103_);
  nor (_33113_, _33109_, _03362_);
  and (_33114_, _03568_, _03226_);
  not (_33116_, _33114_);
  and (_33117_, _04815_, _33116_);
  not (_33118_, _33117_);
  nor (_33119_, _33118_, _33113_);
  nand (_33120_, _33119_, _33112_);
  nor (_33121_, _33117_, _03356_);
  nor (_33122_, _33121_, _03650_);
  and (_33123_, _33122_, _33120_);
  and (_33124_, _11467_, _03650_);
  or (_33125_, _33124_, _08445_);
  nor (_33127_, _33125_, _33123_);
  and (_33128_, _08445_, _03362_);
  or (_33129_, _33128_, _33127_);
  nand (_33130_, _33129_, _11785_);
  and (_33131_, _11784_, _03348_);
  nor (_33132_, _33131_, _03561_);
  nand (_33133_, _33132_, _33130_);
  and (_33134_, _03561_, _03356_);
  nor (_33135_, _33134_, _03227_);
  nand (_33136_, _33135_, _33133_);
  and (_33138_, _03943_, _03227_);
  nor (_33139_, _33138_, _11826_);
  nand (_33140_, _33139_, _33136_);
  and (_33141_, _08820_, _03356_);
  and (_33142_, _32962_, _11832_);
  or (_33143_, _33142_, _33141_);
  and (_33144_, _33143_, _11826_);
  nor (_33145_, _33144_, _11845_);
  and (_33146_, _33145_, _33140_);
  or (_33147_, _33146_, _32937_);
  nand (_33149_, _33147_, _11843_);
  nor (_33150_, _11843_, _03356_);
  nor (_33151_, _33150_, _03649_);
  and (_33152_, _33151_, _33149_);
  and (_33153_, _11467_, _03649_);
  or (_33154_, _33153_, _03778_);
  nor (_33155_, _33154_, _33152_);
  and (_33156_, _03778_, _03362_);
  or (_33157_, _33156_, _33155_);
  nand (_33158_, _33157_, _32301_);
  and (_33160_, _03943_, _03231_);
  nor (_33161_, _33160_, _11856_);
  nand (_33162_, _33161_, _33158_);
  nor (_33163_, _32962_, _11832_);
  nor (_33164_, _08820_, _03356_);
  nor (_33165_, _33164_, _11857_);
  not (_33166_, _33165_);
  nor (_33167_, _33166_, _33163_);
  nor (_33168_, _33167_, _11865_);
  and (_33169_, _33168_, _33162_);
  or (_33171_, _33169_, _32936_);
  nand (_33172_, _33171_, _11367_);
  nor (_33173_, _11367_, _03356_);
  nor (_33174_, _33173_, _03655_);
  and (_33175_, _33174_, _33172_);
  and (_33176_, _11467_, _03655_);
  or (_33177_, _33176_, _03773_);
  nor (_33178_, _33177_, _33175_);
  and (_33179_, _03773_, _03362_);
  or (_33180_, _33179_, _33178_);
  nand (_33182_, _33180_, _32298_);
  and (_33183_, _03943_, _03238_);
  nor (_33184_, _33183_, _11363_);
  nand (_33185_, _33184_, _33182_);
  and (_33186_, _03356_, \oc8051_golden_model_1.PSW [7]);
  and (_33187_, _32962_, _07911_);
  or (_33188_, _33187_, _33186_);
  and (_33189_, _33188_, _11363_);
  nor (_33190_, _33189_, _11877_);
  and (_33191_, _33190_, _33185_);
  or (_33193_, _33191_, _32935_);
  nand (_33194_, _33193_, _11357_);
  nor (_33195_, _11357_, _03356_);
  nor (_33196_, _33195_, _03653_);
  and (_33197_, _33196_, _33194_);
  and (_33198_, _11467_, _03653_);
  or (_33199_, _33198_, _03786_);
  nor (_33200_, _33199_, _33197_);
  and (_33201_, _03786_, _03362_);
  or (_33202_, _33201_, _33200_);
  nand (_33204_, _33202_, _32295_);
  and (_33205_, _03943_, _03236_);
  nor (_33206_, _33205_, _11893_);
  nand (_33207_, _33206_, _33204_);
  nor (_33208_, _32962_, _07911_);
  nor (_33209_, _03356_, \oc8051_golden_model_1.PSW [7]);
  nor (_33210_, _33209_, _11894_);
  not (_33211_, _33210_);
  nor (_33212_, _33211_, _33208_);
  nor (_33213_, _33212_, _11898_);
  and (_33215_, _33213_, _33207_);
  or (_33216_, _33215_, _32934_);
  nand (_33217_, _33216_, _08570_);
  nor (_33218_, _08570_, _03356_);
  nor (_33219_, _33218_, _08600_);
  nand (_33220_, _33219_, _33217_);
  and (_33221_, _08600_, _03318_);
  nor (_33222_, _33221_, _03792_);
  and (_33223_, _33222_, _33220_);
  and (_33224_, _06714_, _03792_);
  or (_33226_, _33224_, _33223_);
  nand (_33227_, _33226_, _06475_);
  and (_33228_, _03943_, _03248_);
  nor (_33229_, _33228_, _03652_);
  nand (_33230_, _33229_, _33227_);
  nor (_33231_, _11467_, _09914_);
  and (_33232_, _32947_, _09914_);
  or (_33233_, _33232_, _03796_);
  nor (_33234_, _33233_, _33231_);
  nor (_33235_, _33234_, _11919_);
  and (_33237_, _33235_, _33230_);
  or (_33238_, _33237_, _32933_);
  nand (_33239_, _33238_, _08721_);
  nor (_33240_, _08721_, _03356_);
  nor (_33241_, _33240_, _08769_);
  nand (_33242_, _33241_, _33239_);
  and (_33243_, _08769_, _03318_);
  nor (_33244_, _33243_, _03521_);
  and (_33245_, _33244_, _33242_);
  and (_33246_, _06714_, _03521_);
  or (_33248_, _33246_, _33245_);
  nand (_33249_, _33248_, _32287_);
  and (_33250_, _03943_, _03246_);
  nor (_33251_, _33250_, _03519_);
  nand (_33252_, _33251_, _33249_);
  nor (_33253_, _32946_, _09914_);
  and (_33254_, _11468_, _09914_);
  nor (_33255_, _33254_, _33253_);
  and (_33256_, _33255_, _03519_);
  nor (_33257_, _33256_, _11946_);
  nand (_33259_, _33257_, _33252_);
  nor (_33260_, _11945_, _03318_);
  nor (_33261_, _33260_, _03809_);
  and (_33262_, _33261_, _33259_);
  or (_33263_, _33262_, _32932_);
  nand (_33264_, _33263_, _11952_);
  nor (_33265_, _11952_, _32942_);
  nor (_33266_, _33265_, _05047_);
  nand (_33267_, _33266_, _33264_);
  and (_33268_, _05047_, _03943_);
  nor (_33270_, _33268_, _03205_);
  nand (_33271_, _33270_, _33267_);
  and (_33272_, _33255_, _03205_);
  nor (_33273_, _33272_, _11968_);
  nand (_33274_, _33273_, _33271_);
  nor (_33275_, _11967_, _03318_);
  nor (_33276_, _33275_, _03816_);
  and (_33277_, _33276_, _33274_);
  or (_33278_, _33277_, _32931_);
  nand (_33279_, _33278_, _11974_);
  nor (_33281_, _11974_, _32942_);
  nor (_33282_, _33281_, _11984_);
  nand (_33283_, _33282_, _33279_);
  and (_33284_, _11984_, _03943_);
  nor (_33285_, _33284_, _11982_);
  and (_33286_, _33285_, _33283_);
  and (_33287_, _11982_, _03318_);
  or (_33288_, _33287_, _33286_);
  or (_33289_, _33288_, _43231_);
  or (_33290_, _43227_, \oc8051_golden_model_1.PC [2]);
  and (_33292_, _33290_, _41991_);
  and (_43612_, _33292_, _33289_);
  and (_33293_, _03816_, _03210_);
  and (_33294_, _03809_, _03210_);
  nor (_33295_, _11353_, _03701_);
  nor (_33296_, _11355_, _03701_);
  nor (_33297_, _11361_, _03701_);
  nor (_33298_, _11370_, _03701_);
  nor (_33299_, _11841_, _03701_);
  and (_33300_, _08445_, _03211_);
  and (_33302_, _03500_, _03211_);
  nor (_33303_, _11381_, _03701_);
  nor (_33304_, _32667_, _03210_);
  and (_33305_, _10096_, _03309_);
  and (_33306_, _03947_, _03766_);
  nor (_33307_, _11540_, _03701_);
  nand (_33308_, _03946_, _03211_);
  and (_33309_, _11531_, \oc8051_golden_model_1.PC [3]);
  or (_33310_, _33309_, _04499_);
  and (_33311_, _33310_, _11537_);
  nor (_33313_, _11531_, _03309_);
  or (_33314_, _33313_, _33311_);
  and (_33315_, _33314_, _33308_);
  nand (_33316_, _11536_, _03701_);
  nand (_33317_, _33316_, _32977_);
  nor (_33318_, _33317_, _33315_);
  or (_33319_, _33318_, _33307_);
  nor (_33320_, _33319_, _33306_);
  nor (_33321_, _33320_, _12226_);
  or (_33322_, _11615_, _11614_);
  and (_33324_, _33322_, _11627_);
  nor (_33325_, _33322_, _11627_);
  nor (_33326_, _33325_, _33324_);
  nand (_33327_, _33326_, _11556_);
  or (_33328_, _11556_, _03211_);
  and (_33329_, _33328_, _12226_);
  and (_33330_, _33329_, _33327_);
  or (_33331_, _33330_, _33321_);
  nand (_33332_, _33331_, _06068_);
  and (_33333_, _04509_, _03309_);
  nor (_33334_, _33333_, _03599_);
  nand (_33335_, _33334_, _33332_);
  or (_33336_, _11465_, _11464_);
  and (_33337_, _33336_, _11481_);
  nor (_33338_, _33336_, _11481_);
  nor (_33339_, _33338_, _33337_);
  or (_33340_, _33339_, _11397_);
  and (_33341_, _33340_, _03599_);
  or (_33342_, _11462_, _11526_);
  nand (_33343_, _33342_, _33341_);
  and (_33346_, _33343_, _11391_);
  nand (_33347_, _33346_, _33335_);
  nor (_33348_, _11391_, _03701_);
  nor (_33349_, _33348_, _03515_);
  nand (_33350_, _33349_, _33347_);
  and (_33351_, _03515_, _03210_);
  nor (_33352_, _33351_, _04857_);
  nand (_33353_, _33352_, _33350_);
  and (_33354_, _03766_, _04857_);
  nor (_33355_, _33354_, _03597_);
  nand (_33357_, _33355_, _33353_);
  and (_33358_, _03597_, _03210_);
  nor (_33359_, _33358_, _33003_);
  nand (_33360_, _33359_, _33357_);
  nor (_33361_, _11684_, _03701_);
  nor (_33362_, _33361_, _03603_);
  nand (_33363_, _33362_, _33360_);
  and (_33364_, _03603_, _03210_);
  nor (_33365_, _33364_, _11694_);
  nand (_33366_, _33365_, _33363_);
  nor (_33368_, _11692_, _03701_);
  nor (_33369_, _33368_, _03511_);
  nand (_33370_, _33369_, _33366_);
  and (_33371_, _03511_, _03210_);
  nor (_33372_, _33371_, _11696_);
  nand (_33373_, _33372_, _33370_);
  and (_33374_, _03766_, _11696_);
  nor (_33375_, _33374_, _03510_);
  nand (_33376_, _33375_, _33373_);
  and (_33377_, _03510_, _03210_);
  nor (_33379_, _33377_, _11706_);
  nand (_33380_, _33379_, _33376_);
  and (_33381_, _11462_, _10037_);
  not (_33382_, _33339_);
  nor (_33383_, _33382_, _10037_);
  or (_33384_, _33383_, _33381_);
  nor (_33385_, _33384_, _09988_);
  nor (_33386_, _33385_, _10041_);
  nand (_33387_, _33386_, _33380_);
  or (_33388_, _33339_, _10089_);
  nand (_33390_, _11463_, _10089_);
  and (_33391_, _33390_, _10041_);
  nand (_33392_, _33391_, _33388_);
  and (_33393_, _33392_, _04046_);
  nand (_33394_, _33393_, _33387_);
  nor (_33395_, _33382_, _09946_);
  not (_33396_, _33395_);
  and (_33397_, _11462_, _09946_);
  nor (_33398_, _33397_, _04046_);
  and (_33399_, _33398_, _33396_);
  nor (_33401_, _33399_, _03676_);
  nand (_33402_, _33401_, _33394_);
  and (_33403_, _11463_, _10133_);
  nor (_33404_, _33339_, _10133_);
  or (_33405_, _33404_, _09916_);
  nor (_33406_, _33405_, _33403_);
  nor (_33407_, _33406_, _10096_);
  and (_33408_, _33407_, _33402_);
  or (_33409_, _33408_, _33305_);
  nand (_33410_, _33409_, _03505_);
  and (_33412_, _03504_, _03211_);
  nor (_33413_, _33412_, _04998_);
  nand (_33414_, _33413_, _33410_);
  nor (_33415_, _03766_, _03253_);
  nor (_33416_, _33415_, _32668_);
  and (_33417_, _33416_, _33414_);
  or (_33418_, _33417_, _33304_);
  nand (_33419_, _33418_, _11386_);
  nor (_33420_, _11386_, _03701_);
  nor (_33421_, _33420_, _03630_);
  nand (_33423_, _33421_, _33419_);
  and (_33424_, _03630_, _03210_);
  nor (_33425_, _33424_, _32397_);
  nand (_33426_, _33425_, _33423_);
  and (_33427_, _03766_, _32397_);
  nor (_33428_, _33427_, _03629_);
  nand (_33429_, _33428_, _33426_);
  and (_33430_, _03629_, _03210_);
  nor (_33431_, _33430_, _33065_);
  and (_33432_, _33431_, _33429_);
  or (_33434_, _33432_, _33303_);
  nand (_33435_, _33434_, _11379_);
  nor (_33436_, _11379_, _03210_);
  nor (_33437_, _33436_, _03371_);
  nand (_33438_, _33437_, _33435_);
  nor (_33439_, _03285_, _03309_);
  nor (_33440_, _33439_, _03500_);
  and (_33441_, _33440_, _33438_);
  or (_33442_, _33441_, _33302_);
  nand (_33443_, _33442_, _03278_);
  and (_33445_, _03766_, _03497_);
  nor (_33446_, _33445_, _03656_);
  nand (_33447_, _33446_, _33443_);
  and (_33448_, _11462_, _03656_);
  not (_33449_, _33448_);
  and (_33450_, _33449_, _11759_);
  nand (_33451_, _33450_, _33447_);
  nor (_33452_, _11759_, _03210_);
  nor (_33453_, _33452_, _03644_);
  nand (_33454_, _33453_, _33451_);
  nor (_33456_, _11463_, _03275_);
  nor (_33457_, _33456_, _11770_);
  nand (_33458_, _33457_, _33454_);
  nor (_33459_, _11767_, _03701_);
  nor (_33460_, _33459_, _03562_);
  nand (_33461_, _33460_, _33458_);
  and (_33462_, _03562_, _03210_);
  nor (_33463_, _33462_, _03220_);
  nand (_33464_, _33463_, _33461_);
  and (_33465_, _03766_, _03220_);
  nor (_33467_, _33465_, _11372_);
  nand (_33468_, _33467_, _33464_);
  and (_33469_, _33326_, _11372_);
  nor (_33470_, _33469_, _06246_);
  nand (_33471_, _33470_, _33468_);
  nor (_33472_, _05966_, _03210_);
  nor (_33473_, _33472_, _03650_);
  nand (_33474_, _33473_, _33471_);
  and (_33475_, _11462_, _03650_);
  nor (_33476_, _33475_, _08445_);
  and (_33478_, _33476_, _33474_);
  or (_33479_, _33478_, _33300_);
  nand (_33480_, _33479_, _11785_);
  nor (_33481_, _11785_, _03304_);
  nor (_33482_, _33481_, _03561_);
  nand (_33483_, _33482_, _33480_);
  and (_33484_, _03561_, _03210_);
  nor (_33485_, _33484_, _03227_);
  nand (_33486_, _33485_, _33483_);
  and (_33487_, _03766_, _03227_);
  nor (_33489_, _33487_, _11826_);
  nand (_33490_, _33489_, _33486_);
  and (_33491_, _08820_, _03210_);
  and (_33492_, _33326_, _11832_);
  or (_33493_, _33492_, _33491_);
  and (_33494_, _33493_, _11826_);
  nor (_33495_, _33494_, _11845_);
  and (_33496_, _33495_, _33490_);
  or (_33497_, _33496_, _33299_);
  nand (_33498_, _33497_, _11843_);
  nor (_33500_, _11843_, _03210_);
  nor (_33501_, _33500_, _03649_);
  and (_33502_, _33501_, _33498_);
  and (_33503_, _11462_, _03649_);
  or (_33504_, _33503_, _03778_);
  nor (_33505_, _33504_, _33502_);
  and (_33506_, _03778_, _03211_);
  or (_33507_, _33506_, _33505_);
  nand (_33508_, _33507_, _32301_);
  and (_33509_, _03766_, _03231_);
  nor (_33511_, _33509_, _11856_);
  nand (_33512_, _33511_, _33508_);
  nor (_33513_, _33326_, _11832_);
  nor (_33514_, _08820_, _03210_);
  nor (_33515_, _33514_, _11857_);
  not (_33516_, _33515_);
  nor (_33517_, _33516_, _33513_);
  nor (_33518_, _33517_, _11865_);
  and (_33519_, _33518_, _33512_);
  or (_33520_, _33519_, _33298_);
  nand (_33522_, _33520_, _11367_);
  nor (_33523_, _11367_, _03210_);
  nor (_33524_, _33523_, _03655_);
  and (_33525_, _33524_, _33522_);
  and (_33526_, _11462_, _03655_);
  or (_33527_, _33526_, _03773_);
  nor (_33528_, _33527_, _33525_);
  and (_33529_, _03773_, _03211_);
  or (_33530_, _33529_, _33528_);
  nand (_33531_, _33530_, _32298_);
  and (_33533_, _03766_, _03238_);
  nor (_33534_, _33533_, _11363_);
  nand (_33535_, _33534_, _33531_);
  and (_33536_, _03210_, \oc8051_golden_model_1.PSW [7]);
  and (_33537_, _33326_, _07911_);
  or (_33538_, _33537_, _33536_);
  and (_33539_, _33538_, _11363_);
  nor (_33540_, _33539_, _11877_);
  and (_33541_, _33540_, _33535_);
  or (_33542_, _33541_, _33297_);
  nand (_33544_, _33542_, _11357_);
  nor (_33545_, _11357_, _03210_);
  nor (_33546_, _33545_, _03653_);
  and (_33547_, _33546_, _33544_);
  and (_33548_, _11462_, _03653_);
  or (_33549_, _33548_, _03786_);
  nor (_33550_, _33549_, _33547_);
  and (_33551_, _03786_, _03211_);
  or (_33552_, _33551_, _33550_);
  nand (_33553_, _33552_, _32295_);
  and (_33555_, _03766_, _03236_);
  nor (_33556_, _33555_, _11893_);
  nand (_33557_, _33556_, _33553_);
  nor (_33558_, _33326_, _07911_);
  nor (_33559_, _03210_, \oc8051_golden_model_1.PSW [7]);
  nor (_33560_, _33559_, _11894_);
  not (_33561_, _33560_);
  nor (_33562_, _33561_, _33558_);
  nor (_33563_, _33562_, _11898_);
  and (_33564_, _33563_, _33557_);
  or (_33566_, _33564_, _33296_);
  nand (_33567_, _33566_, _08570_);
  nor (_33568_, _08570_, _03210_);
  nor (_33569_, _33568_, _08600_);
  and (_33570_, _33569_, _33567_);
  and (_33571_, _08600_, _03701_);
  or (_33572_, _33571_, _03792_);
  nor (_33573_, _33572_, _33570_);
  and (_33574_, _06668_, _03792_);
  or (_33575_, _33574_, _33573_);
  nand (_33577_, _33575_, _06475_);
  and (_33578_, _03766_, _03248_);
  nor (_33579_, _33578_, _03652_);
  nand (_33580_, _33579_, _33577_);
  and (_33581_, _33382_, _09914_);
  nor (_33582_, _11462_, _09914_);
  or (_33583_, _33582_, _03796_);
  or (_33584_, _33583_, _33581_);
  and (_33585_, _33584_, _11353_);
  and (_33586_, _33585_, _33580_);
  or (_33588_, _33586_, _33295_);
  nand (_33589_, _33588_, _08721_);
  nor (_33590_, _08721_, _03210_);
  nor (_33591_, _33590_, _08769_);
  nand (_33592_, _33591_, _33589_);
  and (_33593_, _08769_, _03701_);
  nor (_33594_, _33593_, _03521_);
  and (_33595_, _33594_, _33592_);
  and (_33596_, _06668_, _03521_);
  or (_33597_, _33596_, _33595_);
  nand (_33599_, _33597_, _32287_);
  and (_33600_, _03766_, _03246_);
  nor (_33601_, _33600_, _03519_);
  nand (_33602_, _33601_, _33599_);
  nor (_33603_, _33339_, _09914_);
  and (_33604_, _11463_, _09914_);
  nor (_33605_, _33604_, _33603_);
  and (_33606_, _33605_, _03519_);
  nor (_33607_, _33606_, _11946_);
  nand (_33608_, _33607_, _33602_);
  nor (_33610_, _11945_, _03701_);
  nor (_33611_, _33610_, _03809_);
  and (_33612_, _33611_, _33608_);
  or (_33613_, _33612_, _33294_);
  nand (_33614_, _33613_, _11952_);
  nor (_33615_, _11952_, _03309_);
  nor (_33616_, _33615_, _05047_);
  nand (_33617_, _33616_, _33614_);
  and (_33618_, _05047_, _03766_);
  nor (_33619_, _33618_, _03205_);
  nand (_33621_, _33619_, _33617_);
  and (_33622_, _33605_, _03205_);
  nor (_33623_, _33622_, _11968_);
  nand (_33624_, _33623_, _33621_);
  nor (_33625_, _11967_, _03701_);
  nor (_33626_, _33625_, _03816_);
  and (_33627_, _33626_, _33624_);
  or (_33628_, _33627_, _33293_);
  nand (_33629_, _33628_, _11974_);
  nor (_33630_, _11974_, _03309_);
  nor (_33632_, _33630_, _11984_);
  nand (_33633_, _33632_, _33629_);
  and (_33634_, _11984_, _03766_);
  nor (_33635_, _33634_, _11982_);
  and (_33636_, _33635_, _33633_);
  and (_33637_, _11982_, _03701_);
  or (_33638_, _33637_, _33636_);
  or (_33639_, _33638_, _43231_);
  or (_33640_, _43227_, \oc8051_golden_model_1.PC [3]);
  and (_33641_, _33640_, _41991_);
  and (_43613_, _33641_, _33639_);
  and (_33643_, _06344_, _05047_);
  and (_33644_, _06344_, _32397_);
  nor (_33645_, _32667_, _11611_);
  not (_33646_, \oc8051_golden_model_1.PC [4]);
  nor (_33647_, _02925_, _33646_);
  and (_33648_, _02925_, _33646_);
  nor (_33649_, _33648_, _33647_);
  not (_33650_, _33649_);
  and (_33651_, _33650_, _10096_);
  and (_33653_, _11612_, _03511_);
  nor (_33654_, _33649_, _11684_);
  and (_33655_, _06344_, _03947_);
  nor (_33656_, _33649_, _11531_);
  and (_33657_, _11531_, _33646_);
  or (_33658_, _33657_, _33656_);
  and (_33659_, _33658_, _04500_);
  and (_33660_, _11612_, _04499_);
  or (_33661_, _33660_, _04063_);
  or (_33662_, _33661_, _33659_);
  nand (_33664_, _33649_, _11536_);
  and (_33665_, _33664_, _04868_);
  and (_33666_, _33665_, _33662_);
  or (_33667_, _33666_, _32577_);
  or (_33668_, _33667_, _33655_);
  or (_33669_, _33650_, _11540_);
  and (_33670_, _33669_, _06054_);
  and (_33671_, _33670_, _33668_);
  and (_33672_, _11632_, _11629_);
  or (_33673_, _33672_, _11633_);
  or (_33675_, _33673_, _11554_);
  or (_33676_, _11612_, _11556_);
  and (_33677_, _33676_, _33675_);
  and (_33678_, _33677_, _12226_);
  or (_33679_, _33678_, _33671_);
  and (_33680_, _33679_, _06068_);
  and (_33681_, _33650_, _04509_);
  or (_33682_, _33681_, _03599_);
  or (_33683_, _33682_, _33680_);
  and (_33684_, _11486_, _11483_);
  or (_33686_, _33684_, _11487_);
  and (_33687_, _33686_, _11526_);
  or (_33688_, _33687_, _04515_);
  and (_33689_, _11459_, _11397_);
  or (_33690_, _33689_, _33688_);
  and (_33691_, _33690_, _33683_);
  or (_33692_, _33691_, _11392_);
  or (_33693_, _33650_, _11391_);
  and (_33694_, _33693_, _03516_);
  and (_33695_, _33694_, _33692_);
  and (_33697_, _11612_, _03515_);
  or (_33698_, _33697_, _04857_);
  or (_33699_, _33698_, _33695_);
  or (_33700_, _06344_, _03257_);
  and (_33701_, _33700_, _04524_);
  and (_33702_, _33701_, _33699_);
  and (_33703_, _11612_, _03597_);
  or (_33704_, _33703_, _33702_);
  and (_33705_, _33704_, _11684_);
  or (_33706_, _33705_, _33654_);
  and (_33708_, _33706_, _03611_);
  nand (_33709_, _11612_, _03603_);
  nand (_33710_, _33709_, _11692_);
  or (_33711_, _33710_, _33708_);
  or (_33712_, _33650_, _11692_);
  and (_33713_, _33712_, _03512_);
  and (_33714_, _33713_, _33711_);
  or (_33715_, _33714_, _33653_);
  and (_33716_, _33715_, _03260_);
  and (_33717_, _06344_, _11696_);
  or (_33719_, _33717_, _03510_);
  or (_33720_, _33719_, _33716_);
  nand (_33721_, _11611_, _03510_);
  and (_33722_, _33721_, _09988_);
  and (_33723_, _33722_, _33720_);
  or (_33724_, _33686_, _10037_);
  nand (_33725_, _11458_, _10037_);
  and (_33726_, _33725_, _11706_);
  and (_33727_, _33726_, _33724_);
  or (_33728_, _33727_, _33723_);
  and (_33730_, _33728_, _10042_);
  nand (_33731_, _11458_, _10089_);
  or (_33732_, _33686_, _10089_);
  and (_33733_, _33732_, _33731_);
  and (_33734_, _33733_, _10041_);
  or (_33735_, _33734_, _33730_);
  and (_33736_, _33735_, _04046_);
  nand (_33737_, _11458_, _09946_);
  or (_33738_, _33686_, _09946_);
  and (_33739_, _33738_, _03615_);
  and (_33740_, _33739_, _33737_);
  or (_33741_, _33740_, _03676_);
  or (_33742_, _33741_, _33736_);
  not (_33743_, _10133_);
  and (_33744_, _33686_, _33743_);
  and (_33745_, _11459_, _10133_);
  or (_33746_, _33745_, _09916_);
  or (_33747_, _33746_, _33744_);
  and (_33748_, _33747_, _11389_);
  and (_33749_, _33748_, _33742_);
  or (_33751_, _33749_, _33651_);
  and (_33752_, _33751_, _03505_);
  and (_33753_, _11612_, _03504_);
  or (_33754_, _33753_, _04998_);
  or (_33755_, _33754_, _33752_);
  or (_33756_, _06344_, _03253_);
  and (_33757_, _33756_, _32667_);
  and (_33758_, _33757_, _33755_);
  or (_33759_, _33758_, _33645_);
  and (_33760_, _33759_, _11386_);
  nor (_33762_, _33649_, _11386_);
  or (_33763_, _33762_, _03630_);
  or (_33764_, _33763_, _33760_);
  nand (_33765_, _11611_, _03630_);
  and (_33766_, _33765_, _03265_);
  and (_33767_, _33766_, _33764_);
  or (_33768_, _33767_, _33644_);
  and (_33769_, _33768_, _09728_);
  nand (_33770_, _11612_, _03629_);
  nand (_33771_, _33770_, _11381_);
  or (_33773_, _33771_, _33769_);
  or (_33774_, _33650_, _11381_);
  and (_33775_, _33774_, _11379_);
  and (_33776_, _33775_, _33773_);
  nor (_33777_, _11611_, _11379_);
  or (_33778_, _33777_, _03371_);
  or (_33779_, _33778_, _33776_);
  or (_33780_, _33650_, _03285_);
  and (_33781_, _33780_, _03501_);
  and (_33782_, _33781_, _33779_);
  and (_33784_, _11612_, _03500_);
  or (_33785_, _33784_, _33782_);
  and (_33786_, _33785_, _03278_);
  and (_33787_, _06344_, _03497_);
  or (_33788_, _33787_, _03656_);
  or (_33789_, _33788_, _33786_);
  nand (_33790_, _11458_, _03656_);
  and (_33791_, _33790_, _11759_);
  and (_33792_, _33791_, _33789_);
  nor (_33793_, _11611_, _11759_);
  or (_33795_, _33793_, _03644_);
  or (_33796_, _33795_, _33792_);
  or (_33797_, _11459_, _03275_);
  and (_33798_, _33797_, _11767_);
  and (_33799_, _33798_, _33796_);
  nor (_33800_, _33649_, _11767_);
  or (_33801_, _33800_, _03562_);
  or (_33802_, _33801_, _33799_);
  nand (_33803_, _11611_, _03562_);
  and (_33804_, _33803_, _03221_);
  and (_33806_, _33804_, _33802_);
  and (_33807_, _06344_, _03220_);
  or (_33808_, _33807_, _11372_);
  or (_33809_, _33808_, _33806_);
  or (_33810_, _33673_, _11373_);
  and (_33811_, _33810_, _05966_);
  and (_33812_, _33811_, _33809_);
  nor (_33813_, _11611_, _05966_);
  or (_33814_, _33813_, _03650_);
  or (_33815_, _33814_, _33812_);
  nand (_33817_, _11458_, _03650_);
  and (_33818_, _33817_, _08446_);
  and (_33819_, _33818_, _33815_);
  and (_33820_, _11612_, _08445_);
  or (_33821_, _33820_, _11784_);
  or (_33822_, _33821_, _33819_);
  and (_33823_, _11803_, _11800_);
  nor (_33824_, _33823_, _11804_);
  nand (_33825_, _33824_, _11784_);
  and (_33826_, _33825_, _04181_);
  and (_33828_, _33826_, _33822_);
  and (_33829_, _11612_, _03561_);
  or (_33830_, _33829_, _33828_);
  and (_33831_, _33830_, _27673_);
  and (_33832_, _06344_, _03227_);
  or (_33833_, _33832_, _11826_);
  or (_33834_, _33833_, _33831_);
  and (_33835_, _33673_, _11832_);
  nand (_33836_, _11612_, _08820_);
  nand (_33837_, _33836_, _11826_);
  or (_33839_, _33837_, _33835_);
  and (_33840_, _33839_, _33834_);
  or (_33841_, _33840_, _11845_);
  or (_33842_, _33650_, _11841_);
  and (_33843_, _33842_, _11843_);
  and (_33844_, _33843_, _33841_);
  nor (_33845_, _11611_, _11843_);
  or (_33846_, _33845_, _03649_);
  or (_33847_, _33846_, _33844_);
  nand (_33848_, _11458_, _03649_);
  and (_33850_, _33848_, _04589_);
  and (_33851_, _33850_, _33847_);
  and (_33852_, _11612_, _03778_);
  or (_33853_, _33852_, _33851_);
  and (_33854_, _33853_, _32301_);
  and (_33855_, _06344_, _03231_);
  or (_33856_, _33855_, _11856_);
  or (_33857_, _33856_, _33854_);
  and (_33858_, _33673_, _08820_);
  or (_33859_, _11611_, _08820_);
  nand (_33860_, _33859_, _11856_);
  or (_33861_, _33860_, _33858_);
  and (_33862_, _33861_, _33857_);
  or (_33863_, _33862_, _11865_);
  or (_33864_, _33650_, _11370_);
  and (_33865_, _33864_, _11367_);
  and (_33866_, _33865_, _33863_);
  nor (_33867_, _11367_, _11611_);
  or (_33868_, _33867_, _03655_);
  or (_33869_, _33868_, _33866_);
  nand (_33872_, _11458_, _03655_);
  and (_33873_, _33872_, _04594_);
  and (_33874_, _33873_, _33869_);
  and (_33875_, _11612_, _03773_);
  or (_33876_, _33875_, _33874_);
  and (_33877_, _33876_, _32298_);
  and (_33878_, _06344_, _03238_);
  or (_33879_, _33878_, _11363_);
  or (_33880_, _33879_, _33877_);
  and (_33881_, _33673_, _07911_);
  or (_33883_, _11611_, _07911_);
  nand (_33884_, _33883_, _11363_);
  or (_33885_, _33884_, _33881_);
  and (_33886_, _33885_, _33880_);
  or (_33887_, _33886_, _11877_);
  or (_33888_, _33650_, _11361_);
  and (_33889_, _33888_, _11357_);
  and (_33890_, _33889_, _33887_);
  nor (_33891_, _11611_, _11357_);
  or (_33892_, _33891_, _03653_);
  or (_33894_, _33892_, _33890_);
  nand (_33895_, _11458_, _03653_);
  and (_33896_, _33895_, _04606_);
  and (_33897_, _33896_, _33894_);
  and (_33898_, _11612_, _03786_);
  or (_33899_, _33898_, _33897_);
  and (_33900_, _33899_, _32295_);
  and (_33901_, _06344_, _03236_);
  or (_33902_, _33901_, _11893_);
  or (_33903_, _33902_, _33900_);
  and (_33905_, _33673_, \oc8051_golden_model_1.PSW [7]);
  or (_33906_, _11611_, \oc8051_golden_model_1.PSW [7]);
  nand (_33907_, _33906_, _11893_);
  or (_33908_, _33907_, _33905_);
  and (_33909_, _33908_, _33903_);
  or (_33910_, _33909_, _11898_);
  or (_33911_, _33650_, _11355_);
  and (_33912_, _33911_, _08570_);
  and (_33913_, _33912_, _33910_);
  nor (_33914_, _11611_, _08570_);
  or (_33916_, _33914_, _08600_);
  or (_33917_, _33916_, _33913_);
  nand (_33918_, _33649_, _08600_);
  and (_33919_, _33918_, _10680_);
  and (_33920_, _33919_, _33917_);
  and (_33921_, _06806_, _03792_);
  or (_33922_, _33921_, _33920_);
  and (_33923_, _33922_, _06475_);
  and (_33924_, _06344_, _03248_);
  or (_33925_, _33924_, _03652_);
  or (_33927_, _33925_, _33923_);
  or (_33928_, _11459_, _09914_);
  or (_33929_, _33686_, _11920_);
  and (_33930_, _33929_, _33928_);
  or (_33931_, _33930_, _03796_);
  and (_33932_, _33931_, _33927_);
  or (_33933_, _33932_, _11919_);
  or (_33934_, _33650_, _11353_);
  and (_33935_, _33934_, _08721_);
  and (_33936_, _33935_, _33933_);
  nor (_33938_, _11611_, _08721_);
  or (_33939_, _33938_, _08769_);
  or (_33940_, _33939_, _33936_);
  nand (_33941_, _33649_, _08769_);
  and (_33942_, _33941_, _03522_);
  and (_33943_, _33942_, _33940_);
  and (_33944_, _06806_, _03521_);
  or (_33945_, _33944_, _03246_);
  or (_33946_, _33945_, _33943_);
  or (_33947_, _06344_, _32287_);
  and (_33949_, _33947_, _03520_);
  and (_33950_, _33949_, _33946_);
  nand (_33951_, _11458_, _09914_);
  or (_33952_, _33686_, _09914_);
  and (_33953_, _33952_, _33951_);
  and (_33954_, _33953_, _03519_);
  or (_33955_, _33954_, _11946_);
  or (_33956_, _33955_, _33950_);
  or (_33957_, _33650_, _11945_);
  and (_33958_, _33957_, _04260_);
  and (_33960_, _33958_, _33956_);
  nand (_33961_, _11612_, _03809_);
  nand (_33962_, _33961_, _11952_);
  or (_33963_, _33962_, _33960_);
  or (_33964_, _33650_, _11952_);
  and (_33965_, _33964_, _04625_);
  and (_33966_, _33965_, _33963_);
  or (_33967_, _33966_, _33643_);
  and (_33968_, _33967_, _03206_);
  and (_33969_, _33953_, _03205_);
  or (_33971_, _33969_, _11968_);
  nor (_33972_, _33971_, _33968_);
  nor (_33973_, _33650_, _11967_);
  nor (_33974_, _33973_, _03816_);
  not (_33975_, _33974_);
  nor (_33976_, _33975_, _33972_);
  not (_33977_, _11974_);
  and (_33978_, _11612_, _03816_);
  nor (_33979_, _33978_, _33977_);
  not (_33980_, _33979_);
  or (_33982_, _33980_, _33976_);
  nor (_33983_, _33650_, _11974_);
  nor (_33984_, _33983_, _11984_);
  nand (_33985_, _33984_, _33982_);
  and (_33986_, _11984_, _06344_);
  nor (_33987_, _33986_, _11982_);
  and (_33988_, _33987_, _33985_);
  and (_33989_, _33649_, _11982_);
  or (_33990_, _33989_, _33988_);
  or (_33991_, _33990_, _43231_);
  or (_33993_, _43227_, \oc8051_golden_model_1.PC [4]);
  and (_33994_, _33993_, _41991_);
  and (_43614_, _33994_, _33991_);
  and (_33995_, _11606_, _03816_);
  and (_33996_, _11606_, _03809_);
  nor (_33997_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_33998_, _11606_, _02938_);
  nor (_33999_, _33998_, _33997_);
  nor (_34000_, _33999_, _11353_);
  and (_34001_, _06761_, _03792_);
  nor (_34003_, _33999_, _11355_);
  nor (_34004_, _33999_, _11361_);
  nor (_34005_, _33999_, _11370_);
  nor (_34006_, _33999_, _11841_);
  nor (_34007_, _32667_, _11606_);
  not (_34008_, _33999_);
  and (_34009_, _34008_, _10096_);
  and (_34010_, _06313_, _03947_);
  nor (_34011_, _33999_, _11540_);
  not (_34012_, _32977_);
  nor (_34014_, _33999_, _32309_);
  and (_34015_, _11607_, _03946_);
  nor (_34016_, _04499_, \oc8051_golden_model_1.PC [5]);
  and (_34017_, _34016_, _11531_);
  nor (_34018_, _34017_, _34015_);
  nor (_34019_, _34018_, _11536_);
  nor (_34020_, _34019_, _34014_);
  nor (_34021_, _34020_, _34012_);
  or (_34022_, _34021_, _34011_);
  nor (_34023_, _34022_, _34010_);
  nor (_34025_, _34023_, _12226_);
  or (_34026_, _11609_, _11608_);
  not (_34027_, _34026_);
  nor (_34028_, _34027_, _11634_);
  and (_34029_, _34027_, _11634_);
  nor (_34030_, _34029_, _34028_);
  nor (_34031_, _34030_, _11554_);
  or (_34032_, _11607_, _11556_);
  nand (_34033_, _34032_, _12226_);
  nor (_34034_, _34033_, _34031_);
  or (_34036_, _34034_, _34025_);
  nand (_34037_, _34036_, _06068_);
  and (_34038_, _34008_, _04509_);
  nor (_34039_, _34038_, _03599_);
  nand (_34040_, _34039_, _34037_);
  or (_34041_, _11456_, _11455_);
  not (_34042_, _34041_);
  nor (_34043_, _34042_, _11488_);
  and (_34044_, _34042_, _11488_);
  nor (_34045_, _34044_, _34043_);
  not (_34047_, _34045_);
  or (_34048_, _34047_, _11397_);
  nand (_34049_, _34048_, _03599_);
  and (_34050_, _11454_, _11397_);
  or (_34051_, _34050_, _34049_);
  and (_34052_, _34051_, _11391_);
  nand (_34053_, _34052_, _34040_);
  nor (_34054_, _33999_, _11391_);
  nor (_34055_, _34054_, _03515_);
  nand (_34056_, _34055_, _34053_);
  and (_34058_, _11606_, _03515_);
  nor (_34059_, _34058_, _04857_);
  nand (_34060_, _34059_, _34056_);
  and (_34061_, _06313_, _04857_);
  nor (_34062_, _34061_, _03597_);
  nand (_34063_, _34062_, _34060_);
  and (_34064_, _11606_, _03597_);
  nor (_34065_, _34064_, _33003_);
  nand (_34066_, _34065_, _34063_);
  nor (_34067_, _33999_, _11684_);
  nor (_34069_, _34067_, _03603_);
  nand (_34070_, _34069_, _34066_);
  and (_34071_, _11606_, _03603_);
  nor (_34072_, _34071_, _11694_);
  nand (_34073_, _34072_, _34070_);
  nor (_34074_, _33999_, _11692_);
  nor (_34075_, _34074_, _03511_);
  nand (_34076_, _34075_, _34073_);
  and (_34077_, _11606_, _03511_);
  nor (_34078_, _34077_, _11696_);
  nand (_34080_, _34078_, _34076_);
  and (_34081_, _06313_, _11696_);
  nor (_34082_, _34081_, _03510_);
  nand (_34083_, _34082_, _34080_);
  and (_34084_, _11606_, _03510_);
  nor (_34085_, _34084_, _11706_);
  nand (_34086_, _34085_, _34083_);
  and (_34087_, _11453_, _10037_);
  nor (_34088_, _34045_, _10037_);
  or (_34089_, _34088_, _34087_);
  nor (_34091_, _34089_, _09988_);
  nor (_34092_, _34091_, _10041_);
  nand (_34093_, _34092_, _34086_);
  or (_34094_, _34047_, _10089_);
  nand (_34095_, _11454_, _10089_);
  and (_34096_, _34095_, _10041_);
  nand (_34097_, _34096_, _34094_);
  and (_34098_, _34097_, _04046_);
  nand (_34099_, _34098_, _34093_);
  nor (_34100_, _34045_, _09946_);
  not (_34102_, _34100_);
  and (_34103_, _11453_, _09946_);
  nor (_34104_, _34103_, _04046_);
  and (_34105_, _34104_, _34102_);
  nor (_34106_, _34105_, _03676_);
  nand (_34107_, _34106_, _34099_);
  and (_34108_, _11454_, _10133_);
  and (_34109_, _34045_, _33743_);
  or (_34110_, _34109_, _09916_);
  or (_34111_, _34110_, _34108_);
  and (_34113_, _34111_, _11389_);
  and (_34114_, _34113_, _34107_);
  or (_34115_, _34114_, _34009_);
  nand (_34116_, _34115_, _03505_);
  and (_34117_, _11607_, _03504_);
  nor (_34118_, _34117_, _04998_);
  nand (_34119_, _34118_, _34116_);
  nor (_34120_, _06313_, _03253_);
  nor (_34121_, _34120_, _32668_);
  and (_34122_, _34121_, _34119_);
  or (_34124_, _34122_, _34007_);
  nand (_34125_, _34124_, _11386_);
  nor (_34126_, _33999_, _11386_);
  nor (_34127_, _34126_, _03630_);
  nand (_34128_, _34127_, _34125_);
  and (_34129_, _11606_, _03630_);
  nor (_34130_, _34129_, _32397_);
  nand (_34131_, _34130_, _34128_);
  and (_34132_, _06313_, _32397_);
  nor (_34133_, _34132_, _03629_);
  nand (_34134_, _34133_, _34131_);
  and (_34135_, _11606_, _03629_);
  nor (_34136_, _34135_, _33065_);
  and (_34137_, _34136_, _34134_);
  nor (_34138_, _33999_, _11381_);
  or (_34139_, _34138_, _34137_);
  nand (_34140_, _34139_, _11379_);
  nor (_34141_, _11606_, _11379_);
  nor (_34142_, _34141_, _03371_);
  and (_34143_, _34142_, _34140_);
  nor (_34146_, _34008_, _03285_);
  or (_34147_, _34146_, _03500_);
  nor (_34148_, _34147_, _34143_);
  and (_34149_, _11607_, _03500_);
  or (_34150_, _34149_, _34148_);
  nand (_34151_, _34150_, _03278_);
  and (_34152_, _06313_, _03497_);
  nor (_34153_, _34152_, _03656_);
  nand (_34154_, _34153_, _34151_);
  and (_34155_, _11453_, _03656_);
  not (_34157_, _34155_);
  and (_34158_, _34157_, _11759_);
  nand (_34159_, _34158_, _34154_);
  nor (_34160_, _11606_, _11759_);
  nor (_34161_, _34160_, _03644_);
  nand (_34162_, _34161_, _34159_);
  nor (_34163_, _11454_, _03275_);
  nor (_34164_, _34163_, _11770_);
  nand (_34165_, _34164_, _34162_);
  nor (_34166_, _33999_, _11767_);
  nor (_34168_, _34166_, _03562_);
  and (_34169_, _34168_, _34165_);
  and (_34170_, _11606_, _03562_);
  or (_34171_, _34170_, _03220_);
  or (_34172_, _34171_, _34169_);
  and (_34173_, _06313_, _03220_);
  nor (_34174_, _34173_, _11372_);
  nand (_34175_, _34174_, _34172_);
  nor (_34176_, _34030_, _11373_);
  nor (_34177_, _34176_, _06246_);
  nand (_34179_, _34177_, _34175_);
  nor (_34180_, _11606_, _05966_);
  nor (_34181_, _34180_, _03650_);
  nand (_34182_, _34181_, _34179_);
  and (_34183_, _11453_, _03650_);
  nor (_34184_, _34183_, _08445_);
  nand (_34185_, _34184_, _34182_);
  and (_34186_, _11607_, _08445_);
  nor (_34187_, _34186_, _11784_);
  nand (_34188_, _34187_, _34185_);
  and (_34190_, _11805_, _11798_);
  nor (_34191_, _34190_, _11806_);
  and (_34192_, _34191_, _11784_);
  nor (_34193_, _34192_, _03561_);
  and (_34194_, _34193_, _34188_);
  and (_34195_, _11607_, _03561_);
  or (_34196_, _34195_, _34194_);
  nand (_34197_, _34196_, _27673_);
  and (_34198_, _06313_, _03227_);
  nor (_34199_, _34198_, _11826_);
  nand (_34201_, _34199_, _34197_);
  and (_34202_, _11606_, _08820_);
  nor (_34203_, _34030_, _08820_);
  or (_34204_, _34203_, _34202_);
  and (_34205_, _34204_, _11826_);
  nor (_34206_, _34205_, _11845_);
  and (_34207_, _34206_, _34201_);
  or (_34208_, _34207_, _34006_);
  nand (_34209_, _34208_, _11843_);
  nor (_34210_, _11606_, _11843_);
  nor (_34212_, _34210_, _03649_);
  and (_34213_, _34212_, _34209_);
  and (_34214_, _11453_, _03649_);
  or (_34215_, _34214_, _03778_);
  nor (_34216_, _34215_, _34213_);
  and (_34217_, _11607_, _03778_);
  or (_34218_, _34217_, _34216_);
  nand (_34219_, _34218_, _32301_);
  and (_34220_, _06313_, _03231_);
  nor (_34221_, _34220_, _11856_);
  nand (_34223_, _34221_, _34219_);
  and (_34224_, _34030_, _08820_);
  nor (_34225_, _11606_, _08820_);
  nor (_34226_, _34225_, _11857_);
  not (_34227_, _34226_);
  nor (_34228_, _34227_, _34224_);
  nor (_34229_, _34228_, _11865_);
  and (_34230_, _34229_, _34223_);
  or (_34231_, _34230_, _34005_);
  nand (_34232_, _34231_, _11367_);
  nor (_34234_, _11367_, _11606_);
  nor (_34235_, _34234_, _03655_);
  and (_34236_, _34235_, _34232_);
  and (_34237_, _11453_, _03655_);
  or (_34238_, _34237_, _03773_);
  nor (_34239_, _34238_, _34236_);
  and (_34240_, _11607_, _03773_);
  or (_34241_, _34240_, _34239_);
  nand (_34242_, _34241_, _32298_);
  and (_34243_, _06313_, _03238_);
  nor (_34245_, _34243_, _11363_);
  nand (_34246_, _34245_, _34242_);
  and (_34247_, _34030_, _07911_);
  nor (_34248_, _11606_, _07911_);
  nor (_34249_, _34248_, _11364_);
  not (_34250_, _34249_);
  nor (_34251_, _34250_, _34247_);
  nor (_34252_, _34251_, _11877_);
  and (_34253_, _34252_, _34246_);
  or (_34254_, _34253_, _34004_);
  nand (_34256_, _34254_, _11357_);
  nor (_34257_, _11606_, _11357_);
  nor (_34258_, _34257_, _03653_);
  and (_34259_, _34258_, _34256_);
  and (_34260_, _11453_, _03653_);
  or (_34261_, _34260_, _03786_);
  nor (_34262_, _34261_, _34259_);
  and (_34263_, _11607_, _03786_);
  or (_34264_, _34263_, _34262_);
  nand (_34265_, _34264_, _32295_);
  and (_34267_, _06313_, _03236_);
  nor (_34268_, _34267_, _11893_);
  nand (_34269_, _34268_, _34265_);
  and (_34270_, _34030_, \oc8051_golden_model_1.PSW [7]);
  nor (_34271_, _11606_, \oc8051_golden_model_1.PSW [7]);
  nor (_34272_, _34271_, _11894_);
  not (_34273_, _34272_);
  nor (_34274_, _34273_, _34270_);
  nor (_34275_, _34274_, _11898_);
  and (_34276_, _34275_, _34269_);
  or (_34278_, _34276_, _34003_);
  nand (_34279_, _34278_, _08570_);
  nor (_34280_, _11606_, _08570_);
  nor (_34281_, _34280_, _08600_);
  nand (_34282_, _34281_, _34279_);
  and (_34283_, _33999_, _08600_);
  nor (_34284_, _34283_, _03792_);
  and (_34285_, _34284_, _34282_);
  or (_34286_, _34285_, _34001_);
  nand (_34287_, _34286_, _06475_);
  and (_34289_, _06313_, _03248_);
  nor (_34290_, _34289_, _03652_);
  nand (_34291_, _34290_, _34287_);
  and (_34292_, _34045_, _09914_);
  nor (_34293_, _11453_, _09914_);
  or (_34294_, _34293_, _03796_);
  or (_34295_, _34294_, _34292_);
  and (_34296_, _34295_, _11353_);
  and (_34297_, _34296_, _34291_);
  or (_34298_, _34297_, _34000_);
  nand (_34300_, _34298_, _08721_);
  nor (_34301_, _11606_, _08721_);
  nor (_34302_, _34301_, _08769_);
  nand (_34303_, _34302_, _34300_);
  and (_34304_, _33999_, _08769_);
  nor (_34305_, _34304_, _03521_);
  and (_34306_, _34305_, _34303_);
  and (_34307_, _06761_, _03521_);
  or (_34308_, _34307_, _34306_);
  nand (_34309_, _34308_, _32287_);
  and (_34311_, _06313_, _03246_);
  nor (_34312_, _34311_, _03519_);
  nand (_34313_, _34312_, _34309_);
  and (_34314_, _11454_, _09914_);
  nor (_34315_, _34047_, _09914_);
  nor (_34316_, _34315_, _34314_);
  and (_34317_, _34316_, _03519_);
  nor (_34318_, _34317_, _11946_);
  nand (_34319_, _34318_, _34313_);
  nor (_34320_, _33999_, _11945_);
  nor (_34322_, _34320_, _03809_);
  and (_34323_, _34322_, _34319_);
  or (_34324_, _34323_, _33996_);
  nand (_34325_, _34324_, _11952_);
  nor (_34326_, _34008_, _11952_);
  nor (_34327_, _34326_, _05047_);
  nand (_34328_, _34327_, _34325_);
  and (_34329_, _06313_, _05047_);
  nor (_34330_, _34329_, _03205_);
  nand (_34331_, _34330_, _34328_);
  and (_34333_, _34316_, _03205_);
  nor (_34334_, _34333_, _11968_);
  nand (_34335_, _34334_, _34331_);
  nor (_34336_, _33999_, _11967_);
  nor (_34337_, _34336_, _03816_);
  and (_34338_, _34337_, _34335_);
  or (_34339_, _34338_, _33995_);
  nand (_34340_, _34339_, _11974_);
  nor (_34341_, _34008_, _11974_);
  nor (_34342_, _34341_, _11984_);
  nand (_34344_, _34342_, _34340_);
  and (_34345_, _11984_, _06313_);
  nor (_34346_, _34345_, _11982_);
  and (_34347_, _34346_, _34344_);
  and (_34348_, _33999_, _11982_);
  or (_34349_, _34348_, _34347_);
  or (_34350_, _34349_, _43231_);
  or (_34351_, _43227_, \oc8051_golden_model_1.PC [5]);
  and (_34352_, _34351_, _41991_);
  and (_43615_, _34352_, _34350_);
  and (_34354_, _11984_, _06281_);
  and (_34355_, _05915_, _11340_);
  nor (_34356_, _34355_, \oc8051_golden_model_1.PC [6]);
  nor (_34357_, _34356_, _11341_);
  not (_34358_, _34357_);
  nor (_34359_, _34358_, _11974_);
  and (_34360_, _06281_, _05047_);
  and (_34361_, _34358_, _08769_);
  and (_34362_, _11446_, _03653_);
  and (_34363_, _11446_, _03655_);
  and (_34365_, _11446_, _03649_);
  nor (_34366_, _32667_, _11598_);
  and (_34367_, _34358_, _10096_);
  nand (_34368_, _11445_, _10037_);
  and (_34369_, _11490_, _11450_);
  or (_34370_, _34369_, _11491_);
  or (_34371_, _34370_, _10037_);
  and (_34372_, _34371_, _34368_);
  and (_34373_, _34372_, _11706_);
  and (_34374_, _11599_, _03511_);
  nor (_34376_, _34357_, _11680_);
  and (_34377_, _06281_, _03947_);
  nor (_34378_, _34357_, _32309_);
  and (_34379_, _11599_, _03946_);
  nor (_34380_, _04499_, \oc8051_golden_model_1.PC [6]);
  and (_34381_, _34380_, _11531_);
  or (_34382_, _34381_, _34379_);
  and (_34383_, _34382_, _11537_);
  or (_34384_, _34383_, _34378_);
  and (_34385_, _34384_, _04868_);
  or (_34387_, _34385_, _32577_);
  or (_34388_, _34387_, _34377_);
  or (_34389_, _34358_, _11540_);
  and (_34390_, _34389_, _06054_);
  and (_34391_, _34390_, _34388_);
  and (_34392_, _11636_, _11603_);
  or (_34393_, _34392_, _11637_);
  or (_34394_, _34393_, _11554_);
  or (_34395_, _11599_, _11556_);
  and (_34396_, _34395_, _12226_);
  and (_34398_, _34396_, _34394_);
  nor (_34399_, _34398_, _34391_);
  nor (_34400_, _34399_, _11675_);
  or (_34401_, _11446_, _11526_);
  or (_34402_, _34370_, _11397_);
  and (_34403_, _34402_, _03599_);
  and (_34404_, _34403_, _34401_);
  or (_34405_, _34404_, _34400_);
  and (_34406_, _34405_, _11391_);
  or (_34407_, _34406_, _34376_);
  and (_34409_, _34407_, _03516_);
  and (_34410_, _11599_, _03515_);
  or (_34411_, _34410_, _04857_);
  or (_34412_, _34411_, _34409_);
  or (_34413_, _06281_, _03257_);
  and (_34414_, _34413_, _04524_);
  and (_34415_, _34414_, _34412_);
  and (_34416_, _11599_, _03597_);
  or (_34417_, _34416_, _34415_);
  and (_34418_, _34417_, _11684_);
  nor (_34420_, _34357_, _11684_);
  or (_34421_, _34420_, _34418_);
  and (_34422_, _34421_, _03611_);
  nand (_34423_, _11599_, _03603_);
  nand (_34424_, _34423_, _11692_);
  or (_34425_, _34424_, _34422_);
  or (_34426_, _34358_, _11692_);
  and (_34427_, _34426_, _03512_);
  and (_34428_, _34427_, _34425_);
  or (_34429_, _34428_, _34374_);
  and (_34431_, _34429_, _03260_);
  and (_34432_, _06281_, _11696_);
  or (_34433_, _34432_, _03510_);
  or (_34434_, _34433_, _34431_);
  nand (_34435_, _11598_, _03510_);
  and (_34436_, _34435_, _09988_);
  and (_34437_, _34436_, _34434_);
  or (_34438_, _34437_, _34373_);
  and (_34439_, _34438_, _32558_);
  nand (_34440_, _11445_, _10089_);
  or (_34442_, _34370_, _10089_);
  and (_34443_, _34442_, _32559_);
  and (_34444_, _34443_, _34440_);
  or (_34445_, _34444_, _03615_);
  or (_34446_, _34445_, _34439_);
  nand (_34447_, _11445_, _09946_);
  or (_34448_, _34370_, _09946_);
  and (_34449_, _34448_, _34447_);
  or (_34450_, _34449_, _04046_);
  and (_34451_, _34450_, _34446_);
  or (_34453_, _34451_, _03676_);
  nand (_34454_, _11445_, _10133_);
  or (_34455_, _34370_, _10133_);
  and (_34456_, _34455_, _34454_);
  or (_34457_, _34456_, _09916_);
  and (_34458_, _34457_, _11389_);
  and (_34459_, _34458_, _34453_);
  or (_34460_, _34459_, _34367_);
  and (_34461_, _34460_, _03505_);
  and (_34462_, _11599_, _03504_);
  or (_34464_, _34462_, _04998_);
  or (_34465_, _34464_, _34461_);
  or (_34466_, _06281_, _03253_);
  and (_34467_, _34466_, _32667_);
  and (_34468_, _34467_, _34465_);
  or (_34469_, _34468_, _34366_);
  and (_34470_, _34469_, _11386_);
  nor (_34471_, _34357_, _11386_);
  or (_34472_, _34471_, _03630_);
  or (_34473_, _34472_, _34470_);
  nand (_34475_, _11598_, _03630_);
  and (_34476_, _34475_, _03265_);
  and (_34477_, _34476_, _34473_);
  and (_34478_, _06281_, _32397_);
  or (_34479_, _34478_, _03629_);
  or (_34480_, _34479_, _34477_);
  nand (_34481_, _11598_, _03629_);
  and (_34482_, _34481_, _11381_);
  and (_34483_, _34482_, _34480_);
  nor (_34484_, _34357_, _11381_);
  or (_34486_, _34484_, _11380_);
  or (_34487_, _34486_, _34483_);
  or (_34488_, _11599_, _11379_);
  and (_34489_, _34488_, _03285_);
  and (_34490_, _34489_, _34487_);
  nor (_34491_, _34357_, _03285_);
  or (_34492_, _34491_, _34490_);
  and (_34493_, _34492_, _03501_);
  and (_34494_, _11599_, _03500_);
  or (_34495_, _34494_, _03497_);
  or (_34497_, _34495_, _34493_);
  or (_34498_, _06281_, _03278_);
  and (_34499_, _34498_, _08865_);
  and (_34500_, _34499_, _34497_);
  nand (_34501_, _11446_, _03656_);
  nand (_34502_, _34501_, _11759_);
  or (_34503_, _34502_, _34500_);
  or (_34504_, _11599_, _11759_);
  and (_34505_, _34504_, _03275_);
  and (_34506_, _34505_, _34503_);
  or (_34508_, _11445_, _03275_);
  nand (_34509_, _34508_, _11767_);
  or (_34510_, _34509_, _34506_);
  or (_34511_, _34358_, _11767_);
  and (_34512_, _34511_, _32716_);
  and (_34513_, _34512_, _34510_);
  and (_34514_, _11599_, _03562_);
  or (_34515_, _34514_, _03220_);
  or (_34516_, _34515_, _34513_);
  or (_34517_, _06281_, _03221_);
  and (_34519_, _34517_, _11373_);
  and (_34520_, _34519_, _34516_);
  and (_34521_, _34393_, _11372_);
  or (_34522_, _34521_, _34520_);
  or (_34523_, _34522_, _06246_);
  or (_34524_, _11599_, _05966_);
  and (_34525_, _34524_, _04582_);
  and (_34526_, _34525_, _34523_);
  and (_34527_, _11446_, _03650_);
  or (_34528_, _34527_, _08445_);
  or (_34530_, _34528_, _34526_);
  nand (_34531_, _11598_, _08445_);
  and (_34532_, _34531_, _11785_);
  and (_34533_, _34532_, _34530_);
  and (_34534_, _11807_, _11794_);
  or (_34535_, _34534_, _11808_);
  and (_34536_, _34535_, _11784_);
  or (_34537_, _34536_, _03561_);
  or (_34538_, _34537_, _34533_);
  nand (_34539_, _11598_, _03561_);
  and (_34541_, _34539_, _27673_);
  and (_34542_, _34541_, _34538_);
  and (_34543_, _06281_, _03227_);
  or (_34544_, _34543_, _11826_);
  or (_34545_, _34544_, _34542_);
  and (_34546_, _34393_, _11832_);
  or (_34547_, _11598_, _11832_);
  nand (_34548_, _34547_, _11826_);
  or (_34549_, _34548_, _34546_);
  and (_34550_, _34549_, _11841_);
  and (_34552_, _34550_, _34545_);
  nor (_34553_, _34357_, _11841_);
  or (_34554_, _34553_, _11844_);
  or (_34555_, _34554_, _34552_);
  or (_34556_, _11599_, _11843_);
  and (_34557_, _34556_, _04591_);
  and (_34558_, _34557_, _34555_);
  or (_34559_, _34558_, _34365_);
  and (_34560_, _34559_, _04589_);
  and (_34561_, _11599_, _03778_);
  or (_34563_, _34561_, _03231_);
  or (_34564_, _34563_, _34560_);
  or (_34565_, _06281_, _32301_);
  and (_34566_, _34565_, _34564_);
  or (_34567_, _34566_, _11856_);
  and (_34568_, _34393_, _08820_);
  or (_34569_, _11598_, _08820_);
  nand (_34570_, _34569_, _11856_);
  or (_34571_, _34570_, _34568_);
  and (_34572_, _34571_, _11370_);
  and (_34574_, _34572_, _34567_);
  nor (_34575_, _34357_, _11370_);
  or (_34576_, _34575_, _11368_);
  or (_34577_, _34576_, _34574_);
  or (_34578_, _11367_, _11599_);
  and (_34579_, _34578_, _04596_);
  and (_34580_, _34579_, _34577_);
  or (_34581_, _34580_, _34363_);
  and (_34582_, _34581_, _04594_);
  and (_34583_, _11599_, _03773_);
  or (_34585_, _34583_, _03238_);
  or (_34586_, _34585_, _34582_);
  or (_34587_, _06281_, _32298_);
  and (_34588_, _34587_, _34586_);
  or (_34589_, _34588_, _11363_);
  and (_34590_, _34393_, _07911_);
  or (_34591_, _11598_, _07911_);
  nand (_34592_, _34591_, _11363_);
  or (_34593_, _34592_, _34590_);
  and (_34594_, _34593_, _11361_);
  and (_34596_, _34594_, _34589_);
  nor (_34597_, _34357_, _11361_);
  or (_34598_, _34597_, _11358_);
  or (_34599_, _34598_, _34596_);
  or (_34600_, _11599_, _11357_);
  and (_34601_, _34600_, _04608_);
  and (_34602_, _34601_, _34599_);
  or (_34603_, _34602_, _34362_);
  and (_34604_, _34603_, _04606_);
  and (_34605_, _11599_, _03786_);
  or (_34607_, _34605_, _03236_);
  or (_34608_, _34607_, _34604_);
  or (_34609_, _06281_, _32295_);
  and (_34610_, _34609_, _34608_);
  or (_34611_, _34610_, _11893_);
  and (_34612_, _34393_, \oc8051_golden_model_1.PSW [7]);
  or (_34613_, _11598_, \oc8051_golden_model_1.PSW [7]);
  nand (_34614_, _34613_, _11893_);
  or (_34615_, _34614_, _34612_);
  and (_34616_, _34615_, _11355_);
  and (_34618_, _34616_, _34611_);
  nor (_34619_, _34357_, _11355_);
  or (_34620_, _34619_, _08571_);
  or (_34621_, _34620_, _34618_);
  or (_34622_, _11599_, _08570_);
  and (_34623_, _34622_, _08601_);
  and (_34624_, _34623_, _34621_);
  and (_34625_, _34358_, _08600_);
  or (_34626_, _34625_, _03792_);
  or (_34627_, _34626_, _34624_);
  nand (_34629_, _06531_, _03792_);
  and (_34630_, _34629_, _06475_);
  and (_34631_, _34630_, _34627_);
  and (_34632_, _06281_, _03248_);
  or (_34633_, _34632_, _03652_);
  or (_34634_, _34633_, _34631_);
  nor (_34635_, _11445_, _09914_);
  and (_34636_, _34370_, _09914_);
  or (_34637_, _34636_, _03796_);
  or (_34638_, _34637_, _34635_);
  and (_34640_, _34638_, _11353_);
  and (_34641_, _34640_, _34634_);
  nor (_34642_, _34357_, _11353_);
  or (_34643_, _34642_, _08722_);
  or (_34644_, _34643_, _34641_);
  or (_34645_, _11599_, _08721_);
  and (_34646_, _34645_, _08770_);
  and (_34647_, _34646_, _34644_);
  or (_34648_, _34647_, _34361_);
  and (_34649_, _34648_, _03522_);
  nor (_34651_, _06531_, _03522_);
  or (_34652_, _34651_, _03246_);
  or (_34653_, _34652_, _34649_);
  or (_34654_, _06281_, _32287_);
  and (_34655_, _34654_, _03520_);
  and (_34656_, _34655_, _34653_);
  nand (_34657_, _11445_, _09914_);
  or (_34658_, _34370_, _09914_);
  and (_34659_, _34658_, _34657_);
  and (_34660_, _34659_, _03519_);
  or (_34662_, _34660_, _34656_);
  and (_34663_, _34662_, _11945_);
  nor (_34664_, _34357_, _11945_);
  or (_34665_, _34664_, _34663_);
  and (_34666_, _34665_, _04260_);
  nand (_34667_, _11599_, _03809_);
  nand (_34668_, _34667_, _11952_);
  or (_34669_, _34668_, _34666_);
  or (_34670_, _34358_, _11952_);
  and (_34671_, _34670_, _04625_);
  and (_34673_, _34671_, _34669_);
  or (_34674_, _34673_, _34360_);
  and (_34675_, _34674_, _03206_);
  and (_34676_, _34659_, _03205_);
  or (_34677_, _34676_, _11968_);
  nor (_34678_, _34677_, _34675_);
  nor (_34679_, _34358_, _11967_);
  nor (_34680_, _34679_, _03816_);
  not (_34681_, _34680_);
  nor (_34682_, _34681_, _34678_);
  and (_34684_, _11599_, _03816_);
  nor (_34685_, _34684_, _33977_);
  not (_34686_, _34685_);
  nor (_34687_, _34686_, _34682_);
  or (_34688_, _34687_, _11984_);
  nor (_34689_, _34688_, _34359_);
  or (_34690_, _34689_, _11982_);
  nor (_34691_, _34690_, _34354_);
  and (_34692_, _34357_, _11982_);
  or (_34693_, _34692_, _34691_);
  or (_34695_, _34693_, _43231_);
  or (_34696_, _43227_, \oc8051_golden_model_1.PC [6]);
  and (_34697_, _34696_, _41991_);
  and (_43616_, _34697_, _34695_);
  and (_34698_, _11984_, _05958_);
  and (_34699_, _06059_, _03816_);
  and (_34700_, _06059_, _03809_);
  nor (_34701_, _11341_, \oc8051_golden_model_1.PC [7]);
  nor (_34702_, _34701_, _11342_);
  nor (_34703_, _34702_, _11353_);
  nor (_34705_, _34702_, _11355_);
  nor (_34706_, _34702_, _11361_);
  nor (_34707_, _34702_, _11370_);
  nor (_34708_, _34702_, _11841_);
  and (_34709_, _06221_, _03561_);
  and (_34710_, _05922_, _03656_);
  nor (_34711_, _34702_, _11381_);
  and (_34712_, _05958_, _32397_);
  or (_34713_, _34712_, _03629_);
  nor (_34714_, _32667_, _06059_);
  not (_34716_, _34702_);
  and (_34717_, _34716_, _10096_);
  or (_34718_, _11441_, _11442_);
  and (_34719_, _34718_, _11492_);
  nor (_34720_, _34718_, _11492_);
  nor (_34721_, _34720_, _34719_);
  or (_34722_, _34721_, _10089_);
  nand (_34723_, _10089_, _05923_);
  nand (_34724_, _34723_, _34722_);
  nand (_34725_, _34724_, _10041_);
  or (_34727_, _11526_, _05923_);
  not (_34728_, _34721_);
  or (_34729_, _34728_, _11397_);
  and (_34730_, _34729_, _03599_);
  and (_34731_, _34730_, _34727_);
  and (_34732_, _11554_, _06221_);
  or (_34733_, _11594_, _11595_);
  and (_34734_, _34733_, _11638_);
  nor (_34735_, _34733_, _11638_);
  nor (_34736_, _34735_, _34734_);
  not (_34738_, _34736_);
  and (_34739_, _34738_, _11556_);
  or (_34740_, _34739_, _06054_);
  or (_34741_, _34740_, _34732_);
  and (_34742_, _05958_, _03947_);
  nor (_34743_, _34702_, _32309_);
  and (_34744_, _06221_, _03946_);
  nor (_34745_, _04499_, \oc8051_golden_model_1.PC [7]);
  and (_34746_, _34745_, _11531_);
  nor (_34747_, _34746_, _34744_);
  nor (_34749_, _34747_, _11536_);
  nor (_34750_, _34749_, _34743_);
  nor (_34751_, _34750_, _34012_);
  nor (_34752_, _34702_, _11540_);
  or (_34753_, _34752_, _12226_);
  or (_34754_, _34753_, _34751_);
  or (_34755_, _34754_, _34742_);
  and (_34756_, _34755_, _34741_);
  or (_34757_, _34756_, _04509_);
  nand (_34758_, _34702_, _04509_);
  and (_34759_, _34758_, _04515_);
  and (_34760_, _34759_, _34757_);
  or (_34761_, _34760_, _34731_);
  nand (_34762_, _34761_, _11391_);
  nor (_34763_, _34702_, _11391_);
  nor (_34764_, _34763_, _03515_);
  nand (_34765_, _34764_, _34762_);
  and (_34766_, _06059_, _03515_);
  nor (_34767_, _34766_, _04857_);
  nand (_34768_, _34767_, _34765_);
  and (_34771_, _05958_, _04857_);
  nor (_34772_, _34771_, _03597_);
  nand (_34773_, _34772_, _34768_);
  and (_34774_, _06059_, _03597_);
  nor (_34775_, _34774_, _33003_);
  nand (_34776_, _34775_, _34773_);
  nor (_34777_, _34702_, _11684_);
  nor (_34778_, _34777_, _03603_);
  nand (_34779_, _34778_, _34776_);
  and (_34780_, _06059_, _03603_);
  nor (_34782_, _34780_, _11694_);
  nand (_34783_, _34782_, _34779_);
  nor (_34784_, _34702_, _11692_);
  nor (_34785_, _34784_, _03511_);
  nand (_34786_, _34785_, _34783_);
  and (_34787_, _06059_, _03511_);
  nor (_34788_, _34787_, _11696_);
  nand (_34789_, _34788_, _34786_);
  and (_34790_, _05958_, _11696_);
  nor (_34791_, _34790_, _03510_);
  nand (_34793_, _34791_, _34789_);
  and (_34794_, _06059_, _03510_);
  nor (_34795_, _34794_, _11706_);
  and (_34796_, _34795_, _34793_);
  and (_34797_, _10037_, _05922_);
  nor (_34798_, _34728_, _10037_);
  or (_34799_, _34798_, _09988_);
  nor (_34800_, _34799_, _34797_);
  or (_34801_, _34800_, _34796_);
  nand (_34802_, _34801_, _10042_);
  nand (_34804_, _34802_, _34725_);
  or (_34805_, _34804_, _03615_);
  and (_34806_, _09946_, _05922_);
  nor (_34807_, _34728_, _09946_);
  nor (_34808_, _34807_, _34806_);
  or (_34809_, _34808_, _04046_);
  and (_34810_, _34809_, _34805_);
  or (_34811_, _34810_, _03676_);
  nor (_34812_, _34721_, _10133_);
  and (_34813_, _10133_, _05923_);
  nor (_34815_, _34813_, _09916_);
  not (_34816_, _34815_);
  nor (_34817_, _34816_, _34812_);
  nor (_34818_, _34817_, _10096_);
  and (_34819_, _34818_, _34811_);
  or (_34820_, _34819_, _34717_);
  nand (_34821_, _34820_, _03505_);
  and (_34822_, _06221_, _03504_);
  nor (_34823_, _34822_, _04998_);
  nand (_34824_, _34823_, _34821_);
  nor (_34826_, _05958_, _03253_);
  nor (_34827_, _34826_, _32668_);
  and (_34828_, _34827_, _34824_);
  or (_34829_, _34828_, _34714_);
  nand (_34830_, _34829_, _11386_);
  nor (_34831_, _34702_, _11386_);
  nor (_34832_, _34831_, _03630_);
  nand (_34833_, _34832_, _34830_);
  and (_34834_, _06059_, _03630_);
  nor (_34835_, _34834_, _32397_);
  and (_34837_, _34835_, _34833_);
  or (_34838_, _34837_, _34713_);
  and (_34839_, _06059_, _03629_);
  nor (_34840_, _34839_, _33065_);
  and (_34841_, _34840_, _34838_);
  or (_34842_, _34841_, _34711_);
  nand (_34843_, _34842_, _11379_);
  nor (_34844_, _11379_, _06059_);
  nor (_34845_, _34844_, _03371_);
  and (_34846_, _34845_, _34843_);
  nor (_34848_, _34716_, _03285_);
  or (_34849_, _34848_, _03500_);
  nor (_34850_, _34849_, _34846_);
  and (_34851_, _06221_, _03500_);
  or (_34852_, _34851_, _34850_);
  nand (_34853_, _34852_, _03278_);
  and (_34854_, _05958_, _03497_);
  nor (_34855_, _34854_, _03656_);
  nand (_34856_, _34855_, _34853_);
  nand (_34857_, _34856_, _11759_);
  or (_34859_, _34857_, _34710_);
  nor (_34860_, _11759_, _06059_);
  nor (_34861_, _34860_, _03644_);
  nand (_34862_, _34861_, _34859_);
  nor (_34863_, _05923_, _03275_);
  nor (_34864_, _34863_, _11770_);
  nand (_34865_, _34864_, _34862_);
  nor (_34866_, _34702_, _11767_);
  nor (_34867_, _34866_, _03562_);
  and (_34868_, _34867_, _34865_);
  and (_34870_, _06059_, _03562_);
  or (_34871_, _34870_, _03220_);
  or (_34872_, _34871_, _34868_);
  and (_34873_, _05958_, _03220_);
  nor (_34874_, _34873_, _11372_);
  nand (_34875_, _34874_, _34872_);
  and (_34876_, _34736_, _11372_);
  nor (_34877_, _34876_, _06246_);
  nand (_34878_, _34877_, _34875_);
  nor (_34879_, _06059_, _05966_);
  nor (_34881_, _34879_, _03650_);
  nand (_34882_, _34881_, _34878_);
  and (_34883_, _05922_, _03650_);
  nor (_34884_, _34883_, _08445_);
  nand (_34885_, _34884_, _34882_);
  and (_34886_, _08445_, _06221_);
  nor (_34887_, _34886_, _11784_);
  nand (_34888_, _34887_, _34885_);
  or (_34889_, _11789_, _11790_);
  nor (_34890_, _34889_, _11809_);
  and (_34892_, _34889_, _11809_);
  nor (_34893_, _34892_, _34890_);
  and (_34894_, _34893_, _11784_);
  nor (_34895_, _34894_, _03561_);
  and (_34896_, _34895_, _34888_);
  or (_34897_, _34896_, _34709_);
  nand (_34898_, _34897_, _27673_);
  and (_34899_, _05958_, _03227_);
  nor (_34900_, _34899_, _11826_);
  nand (_34901_, _34900_, _34898_);
  and (_34903_, _08820_, _06059_);
  and (_34904_, _34736_, _11832_);
  or (_34905_, _34904_, _34903_);
  and (_34906_, _34905_, _11826_);
  nor (_34907_, _34906_, _11845_);
  and (_34908_, _34907_, _34901_);
  or (_34909_, _34908_, _34708_);
  nand (_34910_, _34909_, _11843_);
  nor (_34911_, _11843_, _06059_);
  nor (_34912_, _34911_, _03649_);
  and (_34914_, _34912_, _34910_);
  and (_34915_, _05922_, _03649_);
  or (_34916_, _34915_, _03778_);
  nor (_34917_, _34916_, _34914_);
  and (_34918_, _06221_, _03778_);
  or (_34919_, _34918_, _34917_);
  nand (_34920_, _34919_, _32301_);
  and (_34921_, _05958_, _03231_);
  nor (_34922_, _34921_, _11856_);
  nand (_34923_, _34922_, _34920_);
  nor (_34925_, _34736_, _11832_);
  nor (_34926_, _08820_, _06059_);
  nor (_34927_, _34926_, _11857_);
  not (_34928_, _34927_);
  nor (_34929_, _34928_, _34925_);
  nor (_34930_, _34929_, _11865_);
  and (_34931_, _34930_, _34923_);
  or (_34932_, _34931_, _34707_);
  nand (_34933_, _34932_, _11367_);
  nor (_34934_, _11367_, _06059_);
  nor (_34936_, _34934_, _03655_);
  and (_34937_, _34936_, _34933_);
  and (_34938_, _05922_, _03655_);
  or (_34939_, _34938_, _03773_);
  nor (_34940_, _34939_, _34937_);
  and (_34941_, _06221_, _03773_);
  or (_34942_, _34941_, _34940_);
  nand (_34943_, _34942_, _32298_);
  and (_34944_, _05958_, _03238_);
  nor (_34945_, _34944_, _11363_);
  nand (_34947_, _34945_, _34943_);
  and (_34948_, _06059_, \oc8051_golden_model_1.PSW [7]);
  and (_34949_, _34736_, _07911_);
  or (_34950_, _34949_, _34948_);
  and (_34951_, _34950_, _11363_);
  nor (_34952_, _34951_, _11877_);
  and (_34953_, _34952_, _34947_);
  or (_34954_, _34953_, _34706_);
  nand (_34955_, _34954_, _11357_);
  nor (_34956_, _11357_, _06059_);
  nor (_34958_, _34956_, _03653_);
  and (_34959_, _34958_, _34955_);
  and (_34960_, _05922_, _03653_);
  or (_34961_, _34960_, _03786_);
  nor (_34962_, _34961_, _34959_);
  and (_34963_, _06221_, _03786_);
  or (_34964_, _34963_, _34962_);
  nand (_34965_, _34964_, _32295_);
  and (_34966_, _05958_, _03236_);
  nor (_34967_, _34966_, _11893_);
  nand (_34969_, _34967_, _34965_);
  nor (_34970_, _34736_, _07911_);
  nor (_34971_, _06059_, \oc8051_golden_model_1.PSW [7]);
  nor (_34972_, _34971_, _11894_);
  not (_34973_, _34972_);
  nor (_34974_, _34973_, _34970_);
  nor (_34975_, _34974_, _11898_);
  and (_34976_, _34975_, _34969_);
  or (_34977_, _34976_, _34705_);
  nand (_34978_, _34977_, _08570_);
  nor (_34980_, _08570_, _06059_);
  nor (_34981_, _34980_, _08600_);
  nand (_34982_, _34981_, _34978_);
  and (_34983_, _34702_, _08600_);
  nor (_34984_, _34983_, _03792_);
  and (_34985_, _34984_, _34982_);
  nor (_34986_, _06171_, _10680_);
  or (_34987_, _34986_, _34985_);
  nand (_34988_, _34987_, _06475_);
  and (_34989_, _05958_, _03248_);
  nor (_34991_, _34989_, _03652_);
  nand (_34992_, _34991_, _34988_);
  and (_34993_, _34728_, _09914_);
  nor (_34994_, _09914_, _05922_);
  or (_34995_, _34994_, _03796_);
  or (_34996_, _34995_, _34993_);
  and (_34997_, _34996_, _11353_);
  and (_34998_, _34997_, _34992_);
  or (_34999_, _34998_, _34703_);
  nand (_35000_, _34999_, _08721_);
  nor (_35002_, _08721_, _06059_);
  nor (_35003_, _35002_, _08769_);
  nand (_35004_, _35003_, _35000_);
  and (_35005_, _34702_, _08769_);
  nor (_35006_, _35005_, _03521_);
  and (_35007_, _35006_, _35004_);
  nor (_35008_, _06171_, _03522_);
  or (_35009_, _35008_, _35007_);
  nand (_35010_, _35009_, _32287_);
  and (_35011_, _05958_, _03246_);
  nor (_35013_, _35011_, _03519_);
  nand (_35014_, _35013_, _35010_);
  nor (_35015_, _34721_, _09914_);
  and (_35016_, _09914_, _05923_);
  nor (_35017_, _35016_, _35015_);
  and (_35018_, _35017_, _03519_);
  nor (_35019_, _35018_, _11946_);
  nand (_35020_, _35019_, _35014_);
  nor (_35021_, _34702_, _11945_);
  nor (_35022_, _35021_, _03809_);
  and (_35024_, _35022_, _35020_);
  or (_35025_, _35024_, _34700_);
  nand (_35026_, _35025_, _11952_);
  nor (_35027_, _34716_, _11952_);
  nor (_35028_, _35027_, _05047_);
  nand (_35029_, _35028_, _35026_);
  and (_35030_, _05958_, _05047_);
  nor (_35031_, _35030_, _03205_);
  nand (_35032_, _35031_, _35029_);
  and (_35033_, _35017_, _03205_);
  nor (_35035_, _35033_, _11968_);
  nand (_35036_, _35035_, _35032_);
  nor (_35037_, _34702_, _11967_);
  nor (_35038_, _35037_, _03816_);
  and (_35039_, _35038_, _35036_);
  or (_35040_, _35039_, _34699_);
  nand (_35041_, _35040_, _11974_);
  nor (_35042_, _34716_, _11974_);
  nor (_35043_, _35042_, _11984_);
  and (_35044_, _35043_, _35041_);
  or (_35046_, _35044_, _34698_);
  and (_35047_, _35046_, _11990_);
  and (_35048_, _34716_, _11982_);
  nor (_35049_, _35048_, _35047_);
  or (_35050_, _35049_, _43231_);
  or (_35051_, _43227_, \oc8051_golden_model_1.PC [7]);
  and (_35052_, _35051_, _41991_);
  and (_43617_, _35052_, _35050_);
  nor (_35053_, _04042_, _11978_);
  nor (_35054_, _04042_, _11956_);
  and (_35056_, _11497_, _09914_);
  nor (_35057_, _11500_, _11494_);
  nor (_35058_, _35057_, _11501_);
  nor (_35059_, _35058_, _09914_);
  nor (_35060_, _35059_, _35056_);
  and (_35061_, _35060_, _03519_);
  and (_35062_, _04491_, _03521_);
  nand (_35063_, _11497_, _03655_);
  or (_35064_, _11642_, _05966_);
  nor (_35065_, _11372_, _03220_);
  and (_35067_, _11642_, _03562_);
  and (_35068_, _11642_, _03511_);
  nor (_35069_, _03597_, _04857_);
  and (_35070_, _11642_, _03515_);
  nor (_35071_, _11342_, \oc8051_golden_model_1.PC [8]);
  nor (_35072_, _35071_, _11343_);
  and (_35073_, _11540_, _11531_);
  or (_35074_, _35073_, _35072_);
  and (_35075_, _12206_, _03946_);
  nor (_35076_, _35075_, _11536_);
  nor (_35078_, _04499_, \oc8051_golden_model_1.PC [8]);
  nand (_35079_, _35078_, _11531_);
  nand (_35080_, _35079_, _35076_);
  nand (_35081_, _35080_, _32977_);
  and (_35082_, _35081_, _35074_);
  nand (_35083_, _35072_, _11536_);
  nand (_35084_, _35083_, _06054_);
  or (_35085_, _35084_, _35082_);
  nor (_35086_, _11645_, _11640_);
  nor (_35087_, _35086_, _11646_);
  and (_35089_, _35087_, _11556_);
  and (_35090_, _11642_, _11554_);
  or (_35091_, _35090_, _06054_);
  or (_35092_, _35091_, _35089_);
  and (_35093_, _35092_, _35085_);
  or (_35094_, _35093_, _04509_);
  not (_35095_, _35072_);
  nand (_35096_, _35095_, _04509_);
  and (_35097_, _35096_, _04515_);
  and (_35098_, _35097_, _35094_);
  or (_35100_, _35058_, _11397_);
  and (_35101_, _35100_, _03599_);
  or (_35102_, _11496_, _11526_);
  and (_35103_, _35102_, _35101_);
  or (_35104_, _35103_, _11392_);
  or (_35105_, _35104_, _35098_);
  or (_35106_, _35072_, _11391_);
  and (_35107_, _35106_, _03516_);
  and (_35108_, _35107_, _35105_);
  or (_35109_, _35108_, _35070_);
  and (_35111_, _35109_, _35069_);
  nand (_35112_, _11642_, _03597_);
  nand (_35113_, _35112_, _11684_);
  or (_35114_, _35113_, _35111_);
  or (_35115_, _35072_, _11684_);
  and (_35116_, _35115_, _03611_);
  and (_35117_, _35116_, _35114_);
  nand (_35118_, _11642_, _03603_);
  nand (_35119_, _35118_, _11692_);
  or (_35120_, _35119_, _35117_);
  or (_35122_, _35072_, _11692_);
  and (_35123_, _35122_, _03512_);
  and (_35124_, _35123_, _35120_);
  or (_35125_, _35124_, _35068_);
  and (_35126_, _35125_, _11697_);
  nand (_35127_, _11642_, _03510_);
  nand (_35128_, _35127_, _09988_);
  or (_35129_, _35128_, _35126_);
  and (_35130_, _11496_, _10037_);
  not (_35131_, _35058_);
  nor (_35133_, _35131_, _10037_);
  or (_35134_, _35133_, _35130_);
  or (_35135_, _35134_, _09988_);
  and (_35136_, _35135_, _10042_);
  and (_35137_, _35136_, _35129_);
  or (_35138_, _35058_, _10089_);
  nand (_35139_, _11497_, _10089_);
  and (_35140_, _35139_, _10041_);
  and (_35141_, _35140_, _35138_);
  or (_35142_, _35141_, _03615_);
  or (_35144_, _35142_, _35137_);
  and (_35145_, _11496_, _09946_);
  nor (_35146_, _35131_, _09946_);
  or (_35147_, _35146_, _04046_);
  or (_35148_, _35147_, _35145_);
  and (_35149_, _35148_, _09916_);
  and (_35150_, _35149_, _35144_);
  or (_35151_, _35058_, _10133_);
  nand (_35152_, _11497_, _10133_);
  and (_35153_, _35152_, _03676_);
  and (_35155_, _35153_, _35151_);
  or (_35156_, _35155_, _10096_);
  or (_35157_, _35156_, _35150_);
  nand (_35158_, _35095_, _10096_);
  and (_35159_, _35158_, _03505_);
  and (_35160_, _35159_, _35157_);
  and (_35161_, _11642_, _03504_);
  or (_35162_, _35161_, _04998_);
  or (_35163_, _35162_, _35160_);
  and (_35164_, _35163_, _32667_);
  nor (_35166_, _32667_, _12206_);
  or (_35167_, _35166_, _11387_);
  or (_35168_, _35167_, _35164_);
  or (_35169_, _35072_, _11386_);
  and (_35170_, _35169_, _09729_);
  and (_35171_, _35170_, _35168_);
  and (_35172_, _11642_, _03630_);
  or (_35173_, _35172_, _32397_);
  or (_35174_, _35173_, _35171_);
  and (_35175_, _35174_, _09728_);
  nand (_35177_, _11642_, _03629_);
  nand (_35178_, _35177_, _11381_);
  or (_35179_, _35178_, _35175_);
  or (_35180_, _35072_, _11381_);
  and (_35181_, _35180_, _11379_);
  and (_35182_, _35181_, _35179_);
  nor (_35183_, _12206_, _11379_);
  or (_35184_, _35183_, _35182_);
  and (_35185_, _35184_, _03285_);
  nor (_35186_, _35095_, _03285_);
  or (_35188_, _35186_, _03500_);
  or (_35189_, _35188_, _35185_);
  nand (_35190_, _12206_, _03500_);
  and (_35191_, _35190_, _23770_);
  and (_35192_, _35191_, _35189_);
  nand (_35193_, _11496_, _03656_);
  nand (_35194_, _35193_, _11759_);
  or (_35195_, _35194_, _35192_);
  or (_35196_, _11642_, _11759_);
  and (_35197_, _35196_, _03275_);
  and (_35199_, _35197_, _35195_);
  or (_35200_, _11497_, _03275_);
  nand (_35201_, _35200_, _11767_);
  or (_35202_, _35201_, _35199_);
  or (_35203_, _35072_, _11767_);
  and (_35204_, _35203_, _32716_);
  and (_35205_, _35204_, _35202_);
  or (_35206_, _35205_, _35067_);
  and (_35207_, _35206_, _35065_);
  and (_35208_, _35087_, _11372_);
  or (_35210_, _35208_, _06246_);
  or (_35211_, _35210_, _35207_);
  and (_35212_, _35211_, _35064_);
  or (_35213_, _35212_, _03650_);
  nand (_35214_, _11497_, _03650_);
  and (_35215_, _35214_, _08446_);
  and (_35216_, _35215_, _35213_);
  and (_35217_, _11642_, _08445_);
  or (_35218_, _35217_, _11784_);
  or (_35219_, _35218_, _35216_);
  and (_35221_, _11811_, \oc8051_golden_model_1.DPH [0]);
  nor (_35222_, _11811_, \oc8051_golden_model_1.DPH [0]);
  nor (_35223_, _35222_, _35221_);
  or (_35224_, _35223_, _11785_);
  and (_35225_, _35224_, _04181_);
  and (_35226_, _35225_, _35219_);
  and (_35227_, _11642_, _03561_);
  or (_35228_, _35227_, _03227_);
  or (_35229_, _35228_, _35226_);
  and (_35230_, _35229_, _11827_);
  or (_35232_, _35087_, _08820_);
  or (_35233_, _11642_, _11832_);
  and (_35234_, _35233_, _11826_);
  and (_35235_, _35234_, _35232_);
  or (_35236_, _35235_, _11845_);
  or (_35237_, _35236_, _35230_);
  or (_35238_, _35072_, _11841_);
  and (_35239_, _35238_, _11843_);
  and (_35240_, _35239_, _35237_);
  nor (_35241_, _12206_, _11843_);
  or (_35243_, _35241_, _03649_);
  or (_35244_, _35243_, _35240_);
  nand (_35245_, _11497_, _03649_);
  and (_35246_, _35245_, _04589_);
  and (_35247_, _35246_, _35244_);
  and (_35248_, _11642_, _03778_);
  or (_35249_, _35248_, _03231_);
  or (_35250_, _35249_, _35247_);
  and (_35251_, _35250_, _11857_);
  or (_35252_, _35087_, _11832_);
  or (_35254_, _11642_, _08820_);
  and (_35255_, _35254_, _11856_);
  and (_35256_, _35255_, _35252_);
  or (_35257_, _35256_, _11865_);
  or (_35258_, _35257_, _35251_);
  or (_35259_, _35072_, _11370_);
  and (_35260_, _35259_, _11367_);
  and (_35261_, _35260_, _35258_);
  nor (_35262_, _11367_, _12206_);
  or (_35263_, _35262_, _03655_);
  or (_35265_, _35263_, _35261_);
  and (_35266_, _35265_, _35063_);
  or (_35267_, _35266_, _03773_);
  nor (_35268_, _11363_, _03238_);
  nand (_35269_, _12206_, _03773_);
  and (_35270_, _35269_, _35268_);
  and (_35271_, _35270_, _35267_);
  or (_35272_, _35087_, \oc8051_golden_model_1.PSW [7]);
  or (_35273_, _11642_, _07911_);
  and (_35274_, _35273_, _11363_);
  and (_35276_, _35274_, _35272_);
  or (_35277_, _35276_, _11877_);
  or (_35278_, _35277_, _35271_);
  or (_35279_, _35072_, _11361_);
  and (_35280_, _35279_, _11357_);
  and (_35281_, _35280_, _35278_);
  nor (_35282_, _12206_, _11357_);
  or (_35283_, _35282_, _35281_);
  and (_35284_, _35283_, _04608_);
  and (_35285_, _11496_, _03653_);
  or (_35287_, _35285_, _03786_);
  or (_35288_, _35287_, _35284_);
  nor (_35289_, _11893_, _03236_);
  nand (_35290_, _12206_, _03786_);
  and (_35291_, _35290_, _35289_);
  and (_35292_, _35291_, _35288_);
  or (_35293_, _35087_, _07911_);
  or (_35294_, _11642_, \oc8051_golden_model_1.PSW [7]);
  and (_35295_, _35294_, _11893_);
  and (_35296_, _35295_, _35293_);
  or (_35298_, _35296_, _11898_);
  nor (_35299_, _35298_, _35292_);
  nor (_35300_, _35072_, _11355_);
  nor (_35301_, _35300_, _35299_);
  nor (_35302_, _35301_, _08571_);
  nor (_35303_, _11642_, _08570_);
  nor (_35304_, _35303_, _35302_);
  and (_35305_, _35304_, _08601_);
  and (_35306_, _35072_, _08600_);
  or (_35307_, _35306_, _35305_);
  and (_35309_, _35307_, _10680_);
  and (_35310_, _04491_, _03792_);
  or (_35311_, _35310_, _03248_);
  nor (_35312_, _35311_, _35309_);
  nor (_35313_, _35312_, _03652_);
  and (_35314_, _35131_, _09914_);
  nor (_35315_, _11496_, _09914_);
  or (_35316_, _35315_, _03796_);
  or (_35317_, _35316_, _35314_);
  and (_35318_, _35317_, _11353_);
  not (_35320_, _35318_);
  nor (_35321_, _35320_, _35313_);
  nor (_35322_, _35072_, _11353_);
  nor (_35323_, _35322_, _35321_);
  nor (_35324_, _35323_, _08722_);
  nor (_35325_, _11642_, _08721_);
  nor (_35326_, _35325_, _35324_);
  and (_35327_, _35326_, _08770_);
  and (_35328_, _35072_, _08769_);
  or (_35329_, _35328_, _35327_);
  and (_35331_, _35329_, _03522_);
  or (_35332_, _35331_, _03246_);
  nor (_35333_, _35332_, _35062_);
  nor (_35334_, _35333_, _03519_);
  or (_35335_, _35334_, _11946_);
  nor (_35336_, _35335_, _35061_);
  nor (_35337_, _35072_, _11945_);
  nor (_35338_, _35337_, _03809_);
  not (_35339_, _35338_);
  or (_35340_, _35339_, _35336_);
  not (_35342_, _11952_);
  and (_35343_, _11642_, _03809_);
  nor (_35344_, _35343_, _35342_);
  nand (_35345_, _35344_, _35340_);
  nor (_35346_, _35072_, _11952_);
  nor (_35347_, _35346_, _03686_);
  and (_35348_, _35347_, _35345_);
  or (_35349_, _35348_, _35054_);
  nor (_35350_, _03243_, _03205_);
  nand (_35351_, _35350_, _35349_);
  and (_35353_, _35060_, _03205_);
  nor (_35354_, _35353_, _11968_);
  nand (_35355_, _35354_, _35351_);
  nor (_35356_, _35072_, _11967_);
  nor (_35357_, _35356_, _03816_);
  nand (_35358_, _35357_, _35355_);
  and (_35359_, _11642_, _03816_);
  nor (_35360_, _35359_, _33977_);
  nand (_35361_, _35360_, _35358_);
  nor (_35362_, _35072_, _11974_);
  nor (_35364_, _35362_, _03684_);
  and (_35365_, _35364_, _35361_);
  or (_35366_, _35365_, _35053_);
  and (_35367_, _35366_, _24650_);
  and (_35368_, _35072_, _11982_);
  or (_35369_, _35368_, _35367_);
  or (_35370_, _35369_, _43231_);
  or (_35371_, _43227_, \oc8051_golden_model_1.PC [8]);
  and (_35372_, _35371_, _41991_);
  and (_43618_, _35372_, _35370_);
  nor (_35374_, _04434_, _11978_);
  nor (_35375_, _04434_, _11956_);
  nor (_35376_, _11343_, \oc8051_golden_model_1.PC [9]);
  nor (_35377_, _35376_, _11344_);
  nor (_35378_, _35377_, _11353_);
  nor (_35379_, _35377_, _11355_);
  and (_35380_, _11436_, _03653_);
  nor (_35381_, _35377_, _11361_);
  and (_35382_, _11436_, _03655_);
  nor (_35383_, _35377_, _11370_);
  and (_35385_, _11436_, _03649_);
  nor (_35386_, _35377_, _11841_);
  and (_35387_, _11590_, _03562_);
  and (_35388_, _11590_, _03629_);
  nor (_35389_, _35377_, _11386_);
  not (_35390_, _35377_);
  and (_35391_, _35390_, _10096_);
  and (_35392_, _11590_, _03510_);
  nor (_35393_, _11501_, _11498_);
  and (_35394_, _35393_, _11440_);
  nor (_35396_, _35393_, _11440_);
  nor (_35397_, _35396_, _35394_);
  and (_35398_, _35397_, _11526_);
  and (_35399_, _11437_, _11397_);
  nor (_35400_, _35399_, _35398_);
  or (_35401_, _35400_, _04515_);
  and (_35402_, _11590_, _11554_);
  nor (_35403_, _11646_, _11643_);
  and (_35404_, _35403_, _11593_);
  nor (_35405_, _35403_, _11593_);
  nor (_35407_, _35405_, _35404_);
  nor (_35408_, _35407_, _11554_);
  or (_35409_, _35408_, _06054_);
  nor (_35410_, _35409_, _35402_);
  and (_35411_, _32309_, _11540_);
  nor (_35412_, _35411_, _35377_);
  and (_35413_, _12402_, _03946_);
  nor (_35414_, _04499_, \oc8051_golden_model_1.PC [9]);
  and (_35415_, _35414_, _11531_);
  nor (_35416_, _35415_, _35413_);
  nor (_35418_, _35416_, _11536_);
  and (_35419_, _35418_, _32977_);
  nor (_35420_, _35419_, _35412_);
  nor (_35421_, _35420_, _12226_);
  or (_35422_, _35421_, _04509_);
  nor (_35423_, _35422_, _35410_);
  and (_35424_, _35377_, _04509_);
  or (_35425_, _35424_, _03599_);
  or (_35426_, _35425_, _35423_);
  and (_35427_, _35426_, _35401_);
  nor (_35429_, _35427_, _11392_);
  nor (_35430_, _35377_, _11391_);
  nor (_35431_, _35430_, _03515_);
  not (_35432_, _35431_);
  nor (_35433_, _35432_, _35429_);
  and (_35434_, _11590_, _03515_);
  or (_35435_, _35434_, _04857_);
  nor (_35436_, _35435_, _35433_);
  nor (_35437_, _35436_, _03597_);
  and (_35438_, _11590_, _03597_);
  nor (_35440_, _35438_, _33003_);
  not (_35441_, _35440_);
  nor (_35442_, _35441_, _35437_);
  nor (_35443_, _35377_, _11684_);
  nor (_35444_, _35443_, _03603_);
  not (_35445_, _35444_);
  nor (_35446_, _35445_, _35442_);
  and (_35447_, _11590_, _03603_);
  nor (_35448_, _35447_, _11694_);
  not (_35449_, _35448_);
  or (_35451_, _35449_, _35446_);
  nor (_35452_, _35377_, _11692_);
  nor (_35453_, _35452_, _03511_);
  and (_35454_, _35453_, _35451_);
  and (_35455_, _11590_, _03511_);
  or (_35456_, _35455_, _11696_);
  or (_35457_, _35456_, _35454_);
  and (_35458_, _35457_, _04650_);
  or (_35459_, _35458_, _11706_);
  or (_35460_, _35459_, _35392_);
  and (_35462_, _11436_, _10037_);
  nor (_35463_, _35397_, _10037_);
  or (_35464_, _35463_, _35462_);
  nor (_35465_, _35464_, _09988_);
  nor (_35466_, _35465_, _10041_);
  nand (_35467_, _35466_, _35460_);
  nor (_35468_, _35397_, _10089_);
  and (_35469_, _11436_, _10089_);
  nor (_35470_, _35469_, _35468_);
  nor (_35471_, _35470_, _10042_);
  nor (_35473_, _35471_, _03615_);
  nand (_35474_, _35473_, _35467_);
  and (_35475_, _11436_, _09946_);
  not (_35476_, _35475_);
  nor (_35477_, _35397_, _09946_);
  nor (_35478_, _35477_, _04046_);
  and (_35479_, _35478_, _35476_);
  nor (_35480_, _35479_, _03676_);
  nand (_35481_, _35480_, _35474_);
  and (_35482_, _11436_, _10133_);
  nor (_35485_, _35397_, _10133_);
  or (_35486_, _35485_, _35482_);
  and (_35487_, _35486_, _03676_);
  nor (_35488_, _35487_, _10096_);
  and (_35489_, _35488_, _35481_);
  or (_35490_, _35489_, _35391_);
  nand (_35491_, _35490_, _03505_);
  and (_35492_, _12402_, _03504_);
  nor (_35493_, _35492_, _04998_);
  and (_35494_, _35493_, _32667_);
  nand (_35496_, _35494_, _35491_);
  nor (_35497_, _32667_, _12402_);
  nor (_35498_, _35497_, _11387_);
  and (_35499_, _35498_, _35496_);
  or (_35500_, _35499_, _35389_);
  or (_35501_, _35500_, _03630_);
  nand (_35502_, _11590_, _03630_);
  and (_35503_, _35502_, _35501_);
  or (_35504_, _35503_, _32397_);
  nor (_35505_, _35504_, _03629_);
  or (_35508_, _35505_, _35388_);
  nand (_35509_, _35508_, _11381_);
  nor (_35510_, _35390_, _11381_);
  nor (_35511_, _35510_, _11380_);
  nand (_35512_, _35511_, _35509_);
  nor (_35513_, _11590_, _11379_);
  nor (_35514_, _35513_, _03371_);
  nand (_35515_, _35514_, _35512_);
  nor (_35516_, _35390_, _03285_);
  nor (_35517_, _35516_, _03500_);
  nand (_35519_, _35517_, _35515_);
  and (_35520_, _12402_, _03500_);
  nor (_35521_, _35520_, _23771_);
  nand (_35522_, _35521_, _35519_);
  and (_35523_, _11436_, _03656_);
  not (_35524_, _35523_);
  and (_35525_, _35524_, _11759_);
  nand (_35526_, _35525_, _35522_);
  nor (_35527_, _11590_, _11759_);
  nor (_35528_, _35527_, _03644_);
  nand (_35531_, _35528_, _35526_);
  nor (_35532_, _11437_, _03275_);
  nor (_35533_, _35532_, _11770_);
  nand (_35534_, _35533_, _35531_);
  nor (_35535_, _35377_, _11767_);
  nor (_35536_, _35535_, _03562_);
  and (_35537_, _35536_, _35534_);
  or (_35538_, _35537_, _35387_);
  nand (_35539_, _35538_, _35065_);
  nor (_35540_, _35407_, _11373_);
  nor (_35542_, _35540_, _06246_);
  nand (_35543_, _35542_, _35539_);
  nor (_35544_, _11590_, _05966_);
  nor (_35545_, _35544_, _03650_);
  nand (_35546_, _35545_, _35543_);
  and (_35547_, _11436_, _03650_);
  nor (_35548_, _35547_, _08445_);
  nand (_35549_, _35548_, _35546_);
  and (_35550_, _12402_, _08445_);
  nor (_35551_, _35550_, _11784_);
  and (_35554_, _35551_, _35549_);
  nor (_35555_, _35221_, \oc8051_golden_model_1.DPH [1]);
  not (_35556_, _35555_);
  nor (_35557_, _11812_, _11785_);
  and (_35558_, _35557_, _35556_);
  or (_35559_, _35558_, _35554_);
  nand (_35560_, _35559_, _04181_);
  and (_35561_, _11590_, _03561_);
  nor (_35562_, _35561_, _03227_);
  nand (_35563_, _35562_, _35560_);
  nand (_35565_, _35563_, _11827_);
  and (_35566_, _11590_, _08820_);
  nor (_35567_, _35407_, _08820_);
  or (_35568_, _35567_, _35566_);
  and (_35569_, _35568_, _11826_);
  nor (_35570_, _35569_, _11845_);
  and (_35571_, _35570_, _35565_);
  or (_35572_, _35571_, _35386_);
  nand (_35573_, _35572_, _11843_);
  nor (_35574_, _11590_, _11843_);
  nor (_35576_, _35574_, _03649_);
  and (_35577_, _35576_, _35573_);
  or (_35578_, _35577_, _35385_);
  nand (_35579_, _35578_, _04589_);
  and (_35580_, _11590_, _03778_);
  nor (_35581_, _35580_, _03231_);
  nand (_35582_, _35581_, _35579_);
  nand (_35583_, _35582_, _11857_);
  and (_35584_, _35407_, _08820_);
  nor (_35585_, _11590_, _08820_);
  nor (_35587_, _35585_, _11857_);
  not (_35588_, _35587_);
  nor (_35589_, _35588_, _35584_);
  nor (_35590_, _35589_, _11865_);
  and (_35591_, _35590_, _35583_);
  or (_35592_, _35591_, _35383_);
  nand (_35593_, _35592_, _11367_);
  nor (_35594_, _11367_, _11590_);
  nor (_35595_, _35594_, _03655_);
  and (_35596_, _35595_, _35593_);
  or (_35598_, _35596_, _35382_);
  nand (_35599_, _35598_, _04594_);
  and (_35600_, _11590_, _03773_);
  nor (_35601_, _35600_, _03238_);
  nand (_35602_, _35601_, _35599_);
  nand (_35603_, _35602_, _11364_);
  and (_35604_, _11590_, \oc8051_golden_model_1.PSW [7]);
  nor (_35605_, _35407_, \oc8051_golden_model_1.PSW [7]);
  or (_35606_, _35605_, _35604_);
  and (_35607_, _35606_, _11363_);
  nor (_35609_, _35607_, _11877_);
  and (_35610_, _35609_, _35603_);
  or (_35611_, _35610_, _35381_);
  nand (_35612_, _35611_, _11357_);
  nor (_35613_, _11590_, _11357_);
  nor (_35614_, _35613_, _03653_);
  and (_35615_, _35614_, _35612_);
  or (_35616_, _35615_, _35380_);
  nand (_35617_, _35616_, _04606_);
  and (_35618_, _11590_, _03786_);
  nor (_35620_, _35618_, _03236_);
  nand (_35621_, _35620_, _35617_);
  nand (_35622_, _35621_, _11894_);
  and (_35623_, _35407_, \oc8051_golden_model_1.PSW [7]);
  nor (_35624_, _11590_, \oc8051_golden_model_1.PSW [7]);
  nor (_35625_, _35624_, _11894_);
  not (_35626_, _35625_);
  nor (_35627_, _35626_, _35623_);
  nor (_35628_, _35627_, _11898_);
  and (_35629_, _35628_, _35622_);
  or (_35631_, _35629_, _35379_);
  nand (_35632_, _35631_, _08570_);
  nor (_35633_, _11590_, _08570_);
  nor (_35634_, _35633_, _08600_);
  nand (_35635_, _35634_, _35632_);
  and (_35636_, _35377_, _08600_);
  nor (_35637_, _35636_, _03792_);
  nand (_35638_, _35637_, _35635_);
  nor (_35639_, _03652_, _03248_);
  not (_35640_, _35639_);
  and (_35642_, _04699_, _03792_);
  nor (_35643_, _35642_, _35640_);
  nand (_35644_, _35643_, _35638_);
  and (_35645_, _35397_, _09914_);
  nor (_35646_, _11436_, _09914_);
  or (_35647_, _35646_, _03796_);
  nor (_35648_, _35647_, _35645_);
  nor (_35649_, _35648_, _11919_);
  and (_35650_, _35649_, _35644_);
  or (_35651_, _35650_, _35378_);
  nand (_35653_, _35651_, _08721_);
  nor (_35654_, _11590_, _08721_);
  nor (_35655_, _35654_, _08769_);
  nand (_35656_, _35655_, _35653_);
  and (_35657_, _35377_, _08769_);
  nor (_35658_, _35657_, _03521_);
  nand (_35659_, _35658_, _35656_);
  and (_35660_, _04699_, _03521_);
  nor (_35661_, _35660_, _24531_);
  nand (_35662_, _35661_, _35659_);
  and (_35664_, _11436_, _09914_);
  nor (_35665_, _35397_, _09914_);
  or (_35666_, _35665_, _35664_);
  and (_35667_, _35666_, _03519_);
  nor (_35668_, _35667_, _11946_);
  nand (_35669_, _35668_, _35662_);
  nor (_35670_, _35377_, _11945_);
  nor (_35671_, _35670_, _03809_);
  nand (_35672_, _35671_, _35669_);
  and (_35673_, _11590_, _03809_);
  nor (_35675_, _35673_, _35342_);
  nand (_35676_, _35675_, _35672_);
  nor (_35677_, _35377_, _11952_);
  nor (_35678_, _35677_, _03686_);
  and (_35679_, _35678_, _35676_);
  or (_35680_, _35679_, _35375_);
  nand (_35681_, _35680_, _35350_);
  and (_35682_, _35666_, _03205_);
  nor (_35683_, _35682_, _11968_);
  nand (_35684_, _35683_, _35681_);
  nor (_35686_, _35377_, _11967_);
  nor (_35687_, _35686_, _03816_);
  nand (_35688_, _35687_, _35684_);
  and (_35689_, _11590_, _03816_);
  nor (_35690_, _35689_, _33977_);
  nand (_35691_, _35690_, _35688_);
  nor (_35692_, _35377_, _11974_);
  nor (_35693_, _35692_, _03684_);
  and (_35694_, _35693_, _35691_);
  or (_35695_, _35694_, _35374_);
  and (_35697_, _35695_, _24650_);
  and (_35698_, _35377_, _11982_);
  or (_35699_, _35698_, _35697_);
  or (_35700_, _35699_, _43231_);
  or (_35701_, _43227_, \oc8051_golden_model_1.PC [9]);
  and (_35702_, _35701_, _41991_);
  and (_43619_, _35702_, _35700_);
  nor (_35703_, _11344_, \oc8051_golden_model_1.PC [10]);
  nor (_35704_, _35703_, _11345_);
  and (_35705_, _35704_, _11982_);
  or (_35707_, _35704_, _08770_);
  or (_35708_, _35704_, _08601_);
  nand (_35709_, _11423_, _03653_);
  nand (_35710_, _11423_, _03655_);
  nand (_35711_, _11423_, _03649_);
  and (_35712_, _35704_, _11770_);
  and (_35713_, _35704_, _11694_);
  or (_35714_, _35704_, _11684_);
  not (_35715_, _11680_);
  and (_35716_, _35704_, _35715_);
  nor (_35718_, _11505_, _11502_);
  not (_35719_, _35718_);
  and (_35720_, _35719_, _11433_);
  nor (_35721_, _35719_, _11433_);
  nor (_35722_, _35721_, _35720_);
  or (_35723_, _35722_, _11397_);
  or (_35724_, _11422_, _11526_);
  and (_35725_, _35724_, _03599_);
  and (_35726_, _35725_, _35723_);
  and (_35727_, _11578_, _11554_);
  nor (_35729_, _11650_, _11647_);
  not (_35730_, _35729_);
  and (_35731_, _35730_, _11587_);
  nor (_35732_, _35730_, _11587_);
  nor (_35733_, _35732_, _35731_);
  and (_35734_, _35733_, _11556_);
  or (_35735_, _35734_, _35727_);
  or (_35736_, _35735_, _06054_);
  or (_35737_, _35704_, _35411_);
  nand (_35738_, _12607_, _03946_);
  nor (_35740_, _04499_, \oc8051_golden_model_1.PC [10]);
  nand (_35741_, _35740_, _11531_);
  and (_35742_, _35741_, _35738_);
  or (_35743_, _35742_, _11536_);
  and (_35744_, _35743_, _35737_);
  and (_35745_, _35704_, _32577_);
  nand (_35746_, _06054_, _04868_);
  or (_35747_, _35746_, _35745_);
  or (_35748_, _35747_, _35744_);
  and (_35749_, _35748_, _11674_);
  and (_35751_, _35749_, _35736_);
  or (_35752_, _35751_, _35726_);
  and (_35753_, _35752_, _11391_);
  or (_35754_, _35753_, _35716_);
  and (_35755_, _35754_, _03604_);
  nor (_35756_, _12607_, _03604_);
  nor (_35757_, _35756_, _04857_);
  nand (_35758_, _35757_, _11684_);
  or (_35759_, _35758_, _35755_);
  and (_35760_, _35759_, _35714_);
  or (_35762_, _35760_, _03603_);
  nand (_35763_, _12607_, _03603_);
  and (_35764_, _35763_, _11692_);
  and (_35765_, _35764_, _35762_);
  or (_35766_, _35765_, _35713_);
  and (_35767_, _35766_, _03512_);
  and (_35768_, _11578_, _03511_);
  or (_35769_, _35768_, _11696_);
  or (_35770_, _35769_, _35767_);
  and (_35771_, _35770_, _04650_);
  nand (_35773_, _11578_, _03510_);
  nand (_35774_, _35773_, _09988_);
  or (_35775_, _35774_, _35771_);
  or (_35776_, _35722_, _10037_);
  nand (_35777_, _11423_, _10037_);
  and (_35778_, _35777_, _35776_);
  or (_35779_, _35778_, _09988_);
  and (_35780_, _35779_, _10042_);
  and (_35781_, _35780_, _35775_);
  and (_35782_, _35722_, _11713_);
  and (_35784_, _11422_, _10089_);
  or (_35785_, _35784_, _35782_);
  and (_35786_, _35785_, _10041_);
  or (_35787_, _35786_, _03615_);
  or (_35788_, _35787_, _35781_);
  and (_35789_, _11422_, _09946_);
  and (_35790_, _35722_, _11719_);
  or (_35791_, _35790_, _04046_);
  or (_35792_, _35791_, _35789_);
  and (_35793_, _35792_, _09916_);
  and (_35795_, _35793_, _35788_);
  or (_35796_, _35722_, _10133_);
  nand (_35797_, _11423_, _10133_);
  and (_35798_, _35797_, _03676_);
  and (_35799_, _35798_, _35796_);
  or (_35800_, _35799_, _10096_);
  or (_35801_, _35800_, _35795_);
  or (_35802_, _35704_, _11389_);
  and (_35803_, _32667_, _03505_);
  and (_35804_, _35803_, _35802_);
  and (_35806_, _35804_, _35801_);
  nor (_35807_, _35803_, _12607_);
  nand (_35808_, _11386_, _03253_);
  or (_35809_, _35808_, _35807_);
  or (_35810_, _35809_, _35806_);
  or (_35811_, _35704_, _11386_);
  and (_35812_, _35811_, _09729_);
  and (_35813_, _35812_, _35810_);
  or (_35814_, _35813_, _32397_);
  and (_35815_, _35814_, _09728_);
  or (_35817_, _12607_, _03631_);
  nand (_35818_, _35817_, _11381_);
  or (_35819_, _35818_, _35815_);
  or (_35820_, _35704_, _11381_);
  and (_35821_, _35820_, _11379_);
  and (_35822_, _35821_, _35819_);
  nor (_35823_, _12607_, _11379_);
  or (_35824_, _35823_, _03371_);
  or (_35825_, _35824_, _35822_);
  or (_35826_, _35704_, _03285_);
  and (_35828_, _35826_, _03501_);
  and (_35829_, _35828_, _35825_);
  nand (_35830_, _11578_, _03500_);
  nand (_35831_, _35830_, _23770_);
  or (_35832_, _35831_, _35829_);
  nand (_35833_, _11423_, _03656_);
  and (_35834_, _35833_, _11759_);
  and (_35835_, _35834_, _35832_);
  nor (_35836_, _12607_, _11759_);
  or (_35837_, _35836_, _03644_);
  or (_35839_, _35837_, _35835_);
  or (_35840_, _11422_, _03275_);
  and (_35841_, _35840_, _11767_);
  and (_35842_, _35841_, _35839_);
  or (_35843_, _35842_, _35712_);
  and (_35844_, _35843_, _32716_);
  nand (_35845_, _11578_, _03562_);
  nand (_35846_, _35845_, _35065_);
  or (_35847_, _35846_, _35844_);
  or (_35848_, _35733_, _11373_);
  and (_35850_, _35848_, _05966_);
  and (_35851_, _35850_, _35847_);
  nor (_35852_, _12607_, _05966_);
  or (_35853_, _35852_, _03650_);
  or (_35854_, _35853_, _35851_);
  nand (_35855_, _11423_, _03650_);
  and (_35856_, _35855_, _08446_);
  and (_35857_, _35856_, _35854_);
  and (_35858_, _11578_, _08445_);
  or (_35859_, _35858_, _11784_);
  or (_35861_, _35859_, _35857_);
  nor (_35862_, _11812_, \oc8051_golden_model_1.DPH [2]);
  nor (_35863_, _35862_, _11813_);
  or (_35864_, _35863_, _11785_);
  and (_35865_, _35864_, _04181_);
  and (_35866_, _35865_, _35861_);
  and (_35867_, _11578_, _03561_);
  or (_35868_, _35867_, _35866_);
  nand (_35869_, _04756_, _03136_);
  and (_35870_, _35869_, _35868_);
  or (_35872_, _35733_, _08820_);
  or (_35873_, _11578_, _11832_);
  and (_35874_, _35873_, _11826_);
  and (_35875_, _35874_, _35872_);
  or (_35876_, _35875_, _11845_);
  or (_35877_, _35876_, _35870_);
  or (_35878_, _35704_, _11841_);
  and (_35879_, _35878_, _11843_);
  and (_35880_, _35879_, _35877_);
  nor (_35881_, _12607_, _11843_);
  or (_35883_, _35881_, _03649_);
  or (_35884_, _35883_, _35880_);
  and (_35885_, _35884_, _35711_);
  or (_35886_, _35885_, _03778_);
  nand (_35887_, _12607_, _03778_);
  and (_35888_, _35887_, _24039_);
  and (_35889_, _35888_, _35886_);
  or (_35890_, _35733_, _11832_);
  or (_35891_, _11578_, _08820_);
  and (_35892_, _35891_, _11856_);
  and (_35894_, _35892_, _35890_);
  or (_35895_, _35894_, _11865_);
  or (_35896_, _35895_, _35889_);
  or (_35897_, _35704_, _11370_);
  and (_35898_, _35897_, _11367_);
  and (_35899_, _35898_, _35896_);
  nor (_35900_, _11367_, _12607_);
  or (_35901_, _35900_, _03655_);
  or (_35902_, _35901_, _35899_);
  and (_35903_, _35902_, _35710_);
  or (_35905_, _35903_, _03773_);
  nand (_35906_, _12607_, _03773_);
  and (_35907_, _35906_, _35268_);
  and (_35908_, _35907_, _35905_);
  or (_35909_, _35733_, \oc8051_golden_model_1.PSW [7]);
  or (_35910_, _11578_, _07911_);
  and (_35911_, _35910_, _11363_);
  and (_35912_, _35911_, _35909_);
  or (_35913_, _35912_, _11877_);
  or (_35914_, _35913_, _35908_);
  or (_35916_, _35704_, _11361_);
  and (_35917_, _35916_, _11357_);
  and (_35918_, _35917_, _35914_);
  nor (_35919_, _12607_, _11357_);
  or (_35920_, _35919_, _03653_);
  or (_35921_, _35920_, _35918_);
  and (_35922_, _35921_, _35709_);
  or (_35923_, _35922_, _03786_);
  nand (_35924_, _12607_, _03786_);
  and (_35925_, _35924_, _35289_);
  and (_35927_, _35925_, _35923_);
  or (_35928_, _35733_, _07911_);
  or (_35929_, _11578_, \oc8051_golden_model_1.PSW [7]);
  and (_35930_, _35929_, _11893_);
  and (_35931_, _35930_, _35928_);
  or (_35932_, _35931_, _11898_);
  or (_35933_, _35932_, _35927_);
  or (_35934_, _35704_, _11355_);
  and (_35935_, _35934_, _08570_);
  and (_35936_, _35935_, _35933_);
  nor (_35938_, _12607_, _08570_);
  or (_35939_, _35938_, _08600_);
  or (_35940_, _35939_, _35936_);
  and (_35941_, _35940_, _35708_);
  or (_35942_, _35941_, _03792_);
  nand (_35943_, _05130_, _03792_);
  and (_35944_, _35943_, _35639_);
  and (_35945_, _35944_, _35942_);
  or (_35946_, _35722_, _11920_);
  or (_35947_, _11422_, _09914_);
  and (_35949_, _35947_, _03652_);
  and (_35950_, _35949_, _35946_);
  or (_35951_, _35950_, _11919_);
  or (_35952_, _35951_, _35945_);
  or (_35953_, _35704_, _11353_);
  and (_35954_, _35953_, _08721_);
  and (_35955_, _35954_, _35952_);
  nor (_35956_, _12607_, _08721_);
  or (_35957_, _35956_, _08769_);
  or (_35958_, _35957_, _35955_);
  and (_35960_, _35958_, _35707_);
  or (_35961_, _35960_, _03521_);
  nand (_35962_, _05130_, _03521_);
  and (_35963_, _35962_, _24530_);
  and (_35964_, _35963_, _35961_);
  or (_35965_, _35722_, _09914_);
  nand (_35966_, _11423_, _09914_);
  and (_35967_, _35966_, _35965_);
  and (_35968_, _35967_, _03519_);
  or (_35969_, _35968_, _11946_);
  or (_35971_, _35969_, _35964_);
  or (_35972_, _35704_, _11945_);
  and (_35973_, _35972_, _35971_);
  or (_35974_, _35973_, _03809_);
  nand (_35975_, _12607_, _03809_);
  and (_35976_, _35975_, _11952_);
  and (_35977_, _35976_, _35974_);
  and (_35978_, _35704_, _35342_);
  or (_35979_, _35978_, _03686_);
  or (_35980_, _35979_, _35977_);
  nand (_35982_, _03898_, _03686_);
  and (_35983_, _35982_, _35350_);
  and (_35984_, _35983_, _35980_);
  and (_35985_, _35967_, _03205_);
  or (_35986_, _35985_, _11968_);
  or (_35987_, _35986_, _35984_);
  or (_35988_, _35704_, _11967_);
  and (_35989_, _35988_, _35987_);
  or (_35990_, _35989_, _03816_);
  nand (_35991_, _12607_, _03816_);
  and (_35993_, _35991_, _11974_);
  and (_35994_, _35993_, _35990_);
  and (_35995_, _35704_, _33977_);
  or (_35996_, _35995_, _03684_);
  or (_35997_, _35996_, _35994_);
  nand (_35998_, _03898_, _03684_);
  and (_35999_, _35998_, _24650_);
  and (_36000_, _35999_, _35997_);
  or (_36001_, _36000_, _35705_);
  or (_36002_, _36001_, _43231_);
  or (_36004_, _43227_, \oc8051_golden_model_1.PC [10]);
  and (_36005_, _36004_, _41991_);
  and (_43620_, _36005_, _36002_);
  nor (_36006_, _11345_, \oc8051_golden_model_1.PC [11]);
  nor (_36007_, _36006_, _11346_);
  or (_36008_, _36007_, _11353_);
  or (_36009_, _36007_, _11355_);
  or (_36010_, _36007_, _11361_);
  or (_36011_, _36007_, _11370_);
  or (_36012_, _36007_, _11841_);
  or (_36014_, _11582_, _05966_);
  nor (_36015_, _11428_, _03275_);
  nor (_36016_, _35720_, _11424_);
  and (_36017_, _36016_, _11431_);
  nor (_36018_, _36016_, _11431_);
  or (_36019_, _36018_, _36017_);
  or (_36020_, _36019_, _10133_);
  nand (_36021_, _11428_, _10133_);
  and (_36022_, _36021_, _03676_);
  and (_36023_, _36022_, _36020_);
  and (_36025_, _36019_, _11713_);
  and (_36026_, _11427_, _10089_);
  or (_36027_, _36026_, _10042_);
  or (_36028_, _36027_, _36025_);
  and (_36029_, _11582_, _03603_);
  or (_36030_, _36019_, _11397_);
  or (_36031_, _11427_, _11526_);
  and (_36032_, _36031_, _36030_);
  or (_36033_, _36032_, _04515_);
  or (_36034_, _36007_, _35411_);
  or (_36036_, _11582_, _03948_);
  nor (_36037_, _04499_, \oc8051_golden_model_1.PC [11]);
  nand (_36038_, _36037_, _11531_);
  and (_36039_, _36038_, _36036_);
  or (_36040_, _36039_, _11536_);
  and (_36041_, _36040_, _36034_);
  and (_36042_, _11582_, _03947_);
  and (_36043_, _36007_, _32577_);
  or (_36044_, _36043_, _12226_);
  or (_36045_, _36044_, _36042_);
  or (_36047_, _36045_, _36041_);
  and (_36048_, _11582_, _11554_);
  nor (_36049_, _35731_, _11579_);
  and (_36050_, _36049_, _11585_);
  nor (_36051_, _36049_, _11585_);
  or (_36052_, _36051_, _36050_);
  and (_36053_, _36052_, _11556_);
  or (_36054_, _36053_, _36048_);
  or (_36055_, _36054_, _06054_);
  and (_36056_, _36055_, _36047_);
  or (_36058_, _36056_, _11675_);
  and (_36059_, _36058_, _36033_);
  or (_36060_, _36059_, _11392_);
  or (_36061_, _36007_, _11680_);
  and (_36062_, _36061_, _11679_);
  and (_36063_, _36062_, _36060_);
  not (_36064_, _11679_);
  nand (_36065_, _36064_, _11582_);
  nand (_36066_, _36065_, _11684_);
  or (_36067_, _36066_, _36063_);
  or (_36069_, _36007_, _11684_);
  and (_36070_, _36069_, _03611_);
  and (_36071_, _36070_, _36067_);
  or (_36072_, _36071_, _36029_);
  and (_36073_, _36072_, _11692_);
  and (_36074_, _36007_, _11694_);
  or (_36075_, _36074_, _11699_);
  or (_36076_, _36075_, _36073_);
  or (_36077_, _11698_, _11582_);
  and (_36078_, _36077_, _09988_);
  and (_36080_, _36078_, _36076_);
  nand (_36081_, _11428_, _10037_);
  or (_36082_, _36019_, _10037_);
  and (_36083_, _36082_, _11706_);
  and (_36084_, _36083_, _36081_);
  or (_36085_, _36084_, _10041_);
  or (_36086_, _36085_, _36080_);
  and (_36087_, _36086_, _04046_);
  and (_36088_, _36087_, _36028_);
  and (_36089_, _36019_, _11719_);
  and (_36091_, _11427_, _09946_);
  or (_36092_, _36091_, _36089_);
  and (_36093_, _36092_, _03615_);
  or (_36094_, _36093_, _36088_);
  and (_36095_, _36094_, _09916_);
  or (_36096_, _36095_, _36023_);
  and (_36097_, _36096_, _11389_);
  nand (_36098_, _36007_, _10096_);
  nand (_36099_, _36098_, _11734_);
  or (_36100_, _36099_, _36097_);
  or (_36102_, _11734_, _11582_);
  and (_36103_, _36102_, _11386_);
  and (_36104_, _36103_, _36100_);
  not (_36105_, _11741_);
  and (_36106_, _36007_, _11387_);
  or (_36107_, _36106_, _36105_);
  or (_36108_, _36107_, _36104_);
  or (_36109_, _11741_, _11582_);
  and (_36110_, _36109_, _11381_);
  and (_36111_, _36110_, _36108_);
  and (_36113_, _36007_, _33065_);
  or (_36114_, _36113_, _11380_);
  or (_36115_, _36114_, _36111_);
  or (_36116_, _11582_, _11379_);
  and (_36117_, _36116_, _03285_);
  and (_36118_, _36117_, _36115_);
  nand (_36119_, _36007_, _03371_);
  nand (_36120_, _36119_, _11752_);
  or (_36121_, _36120_, _36118_);
  or (_36122_, _11752_, _11582_);
  and (_36124_, _36122_, _08865_);
  and (_36125_, _36124_, _36121_);
  nand (_36126_, _11427_, _03656_);
  nand (_36127_, _36126_, _11759_);
  or (_36128_, _36127_, _36125_);
  or (_36129_, _11582_, _11759_);
  and (_36130_, _36129_, _03275_);
  and (_36131_, _36130_, _36128_);
  or (_36132_, _36131_, _36015_);
  and (_36133_, _36132_, _11767_);
  and (_36135_, _36007_, _11770_);
  or (_36136_, _36135_, _11769_);
  or (_36137_, _36136_, _36133_);
  and (_36138_, _11582_, _11373_);
  or (_36139_, _36138_, _23286_);
  and (_36140_, _36139_, _36137_);
  and (_36141_, _36052_, _11372_);
  or (_36142_, _36141_, _06246_);
  or (_36143_, _36142_, _36140_);
  and (_36144_, _36143_, _36014_);
  or (_36146_, _36144_, _03650_);
  nand (_36147_, _11428_, _03650_);
  and (_36148_, _36147_, _08446_);
  and (_36149_, _36148_, _36146_);
  and (_36150_, _11582_, _08445_);
  or (_36151_, _36150_, _36149_);
  and (_36152_, _36151_, _11785_);
  or (_36153_, _11813_, \oc8051_golden_model_1.DPH [3]);
  nor (_36154_, _11814_, _11785_);
  and (_36155_, _36154_, _36153_);
  or (_36157_, _36155_, _11823_);
  or (_36158_, _36157_, _36152_);
  or (_36159_, _11822_, _11582_);
  and (_36160_, _36159_, _11827_);
  and (_36161_, _36160_, _36158_);
  or (_36162_, _36052_, _08820_);
  or (_36163_, _11582_, _11832_);
  and (_36164_, _36163_, _11826_);
  and (_36165_, _36164_, _36162_);
  or (_36166_, _36165_, _11845_);
  or (_36168_, _36166_, _36161_);
  and (_36169_, _36168_, _36012_);
  or (_36170_, _36169_, _11844_);
  or (_36171_, _11582_, _11843_);
  and (_36172_, _36171_, _04591_);
  and (_36173_, _36172_, _36170_);
  nand (_36174_, _11427_, _03649_);
  nand (_36175_, _36174_, _11853_);
  or (_36176_, _36175_, _36173_);
  or (_36177_, _11853_, _11582_);
  and (_36179_, _36177_, _11857_);
  and (_36180_, _36179_, _36176_);
  or (_36181_, _36052_, _11832_);
  or (_36182_, _11582_, _08820_);
  and (_36183_, _36182_, _11856_);
  and (_36184_, _36183_, _36181_);
  or (_36185_, _36184_, _11865_);
  or (_36186_, _36185_, _36180_);
  and (_36187_, _36186_, _36011_);
  or (_36188_, _36187_, _11368_);
  or (_36190_, _11367_, _11582_);
  and (_36191_, _36190_, _04596_);
  and (_36192_, _36191_, _36188_);
  nand (_36193_, _11427_, _03655_);
  nand (_36194_, _36193_, _10776_);
  or (_36195_, _36194_, _36192_);
  and (_36196_, _11582_, _11364_);
  or (_36197_, _36196_, _24139_);
  and (_36198_, _36197_, _36195_);
  or (_36199_, _36052_, \oc8051_golden_model_1.PSW [7]);
  or (_36201_, _11582_, _07911_);
  and (_36202_, _36201_, _11363_);
  and (_36203_, _36202_, _36199_);
  or (_36204_, _36203_, _11877_);
  or (_36205_, _36204_, _36198_);
  and (_36206_, _36205_, _36010_);
  or (_36207_, _36206_, _11358_);
  or (_36208_, _11582_, _11357_);
  and (_36209_, _36208_, _04608_);
  and (_36210_, _36209_, _36207_);
  nand (_36212_, _11427_, _03653_);
  nand (_36213_, _36212_, _11890_);
  or (_36214_, _36213_, _36210_);
  and (_36215_, _11894_, _11582_);
  or (_36216_, _36215_, _24294_);
  and (_36217_, _36216_, _36214_);
  or (_36218_, _36052_, _07911_);
  or (_36219_, _11582_, \oc8051_golden_model_1.PSW [7]);
  and (_36220_, _36219_, _11893_);
  and (_36221_, _36220_, _36218_);
  or (_36223_, _36221_, _11898_);
  or (_36224_, _36223_, _36217_);
  and (_36225_, _36224_, _36009_);
  or (_36226_, _36225_, _08571_);
  or (_36227_, _11582_, _08570_);
  and (_36228_, _36227_, _08601_);
  and (_36229_, _36228_, _36226_);
  and (_36230_, _36007_, _08600_);
  or (_36231_, _36230_, _03792_);
  or (_36232_, _36231_, _36229_);
  nand (_36234_, _04944_, _03792_);
  and (_36235_, _36234_, _36232_);
  or (_36236_, _36235_, _03248_);
  or (_36237_, _11582_, _06475_);
  and (_36238_, _36237_, _03796_);
  and (_36239_, _36238_, _36236_);
  or (_36240_, _36019_, _11920_);
  or (_36241_, _11427_, _09914_);
  and (_36242_, _36241_, _03652_);
  and (_36243_, _36242_, _36240_);
  or (_36245_, _36243_, _11919_);
  or (_36246_, _36245_, _36239_);
  and (_36247_, _36246_, _36008_);
  or (_36248_, _36247_, _08722_);
  or (_36249_, _11582_, _08721_);
  and (_36250_, _36249_, _08770_);
  and (_36251_, _36250_, _36248_);
  and (_36252_, _36007_, _08769_);
  or (_36253_, _36252_, _03521_);
  or (_36254_, _36253_, _36251_);
  nand (_36256_, _04944_, _03521_);
  and (_36257_, _36256_, _36254_);
  or (_36258_, _36257_, _03246_);
  or (_36259_, _11582_, _32287_);
  and (_36260_, _36259_, _03520_);
  and (_36261_, _36260_, _36258_);
  or (_36262_, _36019_, _09914_);
  nand (_36263_, _11428_, _09914_);
  and (_36264_, _36263_, _36262_);
  and (_36265_, _36264_, _03519_);
  or (_36267_, _36265_, _11946_);
  or (_36268_, _36267_, _36261_);
  or (_36269_, _36007_, _11945_);
  and (_36270_, _36269_, _04260_);
  and (_36271_, _36270_, _36268_);
  nand (_36272_, _11582_, _03809_);
  nand (_36273_, _36272_, _11952_);
  or (_36274_, _36273_, _36271_);
  or (_36275_, _36007_, _11952_);
  and (_36276_, _36275_, _11956_);
  and (_36278_, _36276_, _36274_);
  nor (_36279_, _11956_, _03494_);
  or (_36280_, _36279_, _03243_);
  or (_36281_, _36280_, _36278_);
  or (_36282_, _11582_, _12381_);
  and (_36283_, _36282_, _03206_);
  and (_36284_, _36283_, _36281_);
  and (_36285_, _36264_, _03205_);
  or (_36286_, _36285_, _11968_);
  or (_36287_, _36286_, _36284_);
  or (_36289_, _36007_, _11967_);
  and (_36290_, _36289_, _03820_);
  and (_36291_, _36290_, _36287_);
  nand (_36292_, _11582_, _03816_);
  nand (_36293_, _36292_, _11974_);
  or (_36294_, _36293_, _36291_);
  or (_36295_, _36007_, _11974_);
  and (_36296_, _36295_, _11978_);
  and (_36297_, _36296_, _36294_);
  not (_36298_, _03242_);
  nand (_36300_, _03494_, _36298_);
  and (_36301_, _36300_, _11984_);
  or (_36302_, _36301_, _11982_);
  or (_36303_, _36302_, _36297_);
  or (_36304_, _11582_, _36298_);
  or (_36305_, _36007_, _11990_);
  and (_36306_, _36305_, _36304_);
  and (_36307_, _36306_, _36303_);
  or (_36308_, _36307_, _43231_);
  or (_36309_, _43227_, \oc8051_golden_model_1.PC [11]);
  and (_36311_, _36309_, _41991_);
  and (_43623_, _36311_, _36308_);
  nand (_36312_, _13020_, _03246_);
  nor (_36313_, _11657_, _11655_);
  nor (_36314_, _36313_, _11658_);
  or (_36315_, _36314_, _08820_);
  or (_36316_, _11575_, _11832_);
  and (_36317_, _36316_, _11826_);
  and (_36318_, _36317_, _36315_);
  nor (_36319_, _11419_, _03275_);
  nor (_36321_, _11512_, _11510_);
  nor (_36322_, _36321_, _11513_);
  or (_36323_, _36322_, _10133_);
  nand (_36324_, _11419_, _10133_);
  and (_36325_, _36324_, _03676_);
  and (_36326_, _36325_, _36323_);
  and (_36327_, _11418_, _10089_);
  and (_36328_, _36322_, _11713_);
  or (_36329_, _36328_, _32558_);
  or (_36330_, _36329_, _36327_);
  or (_36332_, _11698_, _11575_);
  or (_36333_, _36322_, _11397_);
  or (_36334_, _11418_, _11526_);
  and (_36335_, _36334_, _03599_);
  and (_36336_, _36335_, _36333_);
  and (_36337_, _11575_, _11554_);
  and (_36338_, _36314_, _11556_);
  or (_36339_, _36338_, _06054_);
  or (_36340_, _36339_, _36337_);
  nand (_36341_, _13020_, _03947_);
  and (_36343_, _36341_, _11540_);
  nand (_36344_, _13020_, _03946_);
  nor (_36345_, _04499_, \oc8051_golden_model_1.PC [12]);
  nand (_36346_, _36345_, _11531_);
  and (_36347_, _36346_, _36344_);
  or (_36348_, _36347_, _11536_);
  nor (_36349_, _11346_, \oc8051_golden_model_1.PC [12]);
  nor (_36350_, _36349_, _11347_);
  or (_36351_, _36350_, _32309_);
  and (_36352_, _36351_, _36348_);
  or (_36354_, _36352_, _03947_);
  and (_36355_, _36354_, _36343_);
  and (_36356_, _36350_, _32577_);
  or (_36357_, _36356_, _12226_);
  or (_36358_, _36357_, _36355_);
  and (_36359_, _36358_, _11674_);
  and (_36360_, _36359_, _36340_);
  or (_36361_, _36360_, _36336_);
  and (_36362_, _36361_, _11391_);
  and (_36363_, _36350_, _35715_);
  or (_36365_, _36363_, _36064_);
  or (_36366_, _36365_, _36362_);
  or (_36367_, _11679_, _11575_);
  and (_36368_, _36367_, _11684_);
  and (_36369_, _36368_, _36366_);
  and (_36370_, _36350_, _33003_);
  or (_36371_, _36370_, _03603_);
  or (_36372_, _36371_, _36369_);
  nand (_36373_, _13020_, _03603_);
  and (_36374_, _36373_, _11692_);
  and (_36376_, _36374_, _36372_);
  and (_36377_, _36350_, _11694_);
  or (_36378_, _36377_, _11699_);
  or (_36379_, _36378_, _36376_);
  and (_36380_, _36379_, _36332_);
  or (_36381_, _36380_, _11706_);
  not (_36382_, _10037_);
  and (_36383_, _36322_, _36382_);
  and (_36384_, _11418_, _10037_);
  or (_36385_, _36384_, _09988_);
  or (_36387_, _36385_, _36383_);
  and (_36388_, _36387_, _36381_);
  or (_36389_, _36388_, _32559_);
  and (_36390_, _36389_, _04046_);
  and (_36391_, _36390_, _36330_);
  and (_36392_, _36322_, _11719_);
  and (_36393_, _11418_, _09946_);
  or (_36394_, _36393_, _36392_);
  and (_36395_, _36394_, _03615_);
  or (_36396_, _36395_, _36391_);
  and (_36398_, _36396_, _09916_);
  or (_36399_, _36398_, _36326_);
  and (_36400_, _36399_, _11389_);
  nand (_36401_, _36350_, _10096_);
  nand (_36402_, _36401_, _11734_);
  or (_36403_, _36402_, _36400_);
  or (_36404_, _11734_, _11575_);
  and (_36405_, _36404_, _11386_);
  and (_36406_, _36405_, _36403_);
  and (_36407_, _36350_, _11387_);
  or (_36409_, _36407_, _36105_);
  or (_36410_, _36409_, _36406_);
  or (_36411_, _11741_, _11575_);
  and (_36412_, _36411_, _11381_);
  and (_36413_, _36412_, _36410_);
  and (_36414_, _36350_, _33065_);
  or (_36415_, _36414_, _11380_);
  or (_36416_, _36415_, _36413_);
  or (_36417_, _11575_, _11379_);
  and (_36418_, _36417_, _03285_);
  and (_36420_, _36418_, _36416_);
  nand (_36421_, _36350_, _03371_);
  nand (_36422_, _36421_, _11752_);
  or (_36423_, _36422_, _36420_);
  or (_36424_, _11752_, _11575_);
  and (_36425_, _36424_, _08865_);
  and (_36426_, _36425_, _36423_);
  nand (_36427_, _11418_, _03656_);
  nand (_36428_, _36427_, _11759_);
  or (_36429_, _36428_, _36426_);
  or (_36431_, _11575_, _11759_);
  and (_36432_, _36431_, _03275_);
  and (_36433_, _36432_, _36429_);
  or (_36434_, _36433_, _36319_);
  and (_36435_, _36434_, _11767_);
  and (_36436_, _36350_, _11770_);
  or (_36437_, _36436_, _11769_);
  or (_36438_, _36437_, _36435_);
  or (_36439_, _11575_, _11374_);
  and (_36440_, _36439_, _11373_);
  and (_36442_, _36440_, _36438_);
  and (_36443_, _36314_, _11372_);
  or (_36444_, _36443_, _06246_);
  or (_36445_, _36444_, _36442_);
  or (_36446_, _11575_, _05966_);
  and (_36447_, _36446_, _04582_);
  and (_36448_, _36447_, _36445_);
  and (_36449_, _11418_, _03650_);
  or (_36450_, _36449_, _08445_);
  or (_36451_, _36450_, _36448_);
  nand (_36453_, _13020_, _08445_);
  and (_36454_, _36453_, _11785_);
  and (_36455_, _36454_, _36451_);
  nor (_36456_, _11814_, \oc8051_golden_model_1.DPH [4]);
  nor (_36457_, _36456_, _11815_);
  and (_36458_, _36457_, _11784_);
  or (_36459_, _36458_, _11823_);
  or (_36460_, _36459_, _36455_);
  or (_36461_, _11822_, _11575_);
  and (_36462_, _36461_, _11827_);
  and (_36464_, _36462_, _36460_);
  or (_36465_, _36464_, _36318_);
  and (_36466_, _36465_, _11841_);
  and (_36467_, _36350_, _11845_);
  or (_36468_, _36467_, _11844_);
  or (_36469_, _36468_, _36466_);
  or (_36470_, _11575_, _11843_);
  and (_36471_, _36470_, _04591_);
  and (_36472_, _36471_, _36469_);
  nand (_36473_, _11418_, _03649_);
  nand (_36475_, _36473_, _11853_);
  or (_36476_, _36475_, _36472_);
  or (_36477_, _11853_, _11575_);
  and (_36478_, _36477_, _11857_);
  and (_36479_, _36478_, _36476_);
  or (_36480_, _36314_, _11832_);
  or (_36481_, _11575_, _08820_);
  and (_36482_, _36481_, _11856_);
  and (_36483_, _36482_, _36480_);
  or (_36484_, _36483_, _36479_);
  and (_36486_, _36484_, _11370_);
  and (_36487_, _36350_, _11865_);
  or (_36488_, _36487_, _11368_);
  or (_36489_, _36488_, _36486_);
  or (_36490_, _11367_, _11575_);
  and (_36491_, _36490_, _04596_);
  and (_36492_, _36491_, _36489_);
  nand (_36493_, _11418_, _03655_);
  nand (_36494_, _36493_, _10776_);
  or (_36495_, _36494_, _36492_);
  nor (_36497_, _13020_, _11363_);
  or (_36498_, _36497_, _24139_);
  and (_36499_, _36498_, _36495_);
  or (_36500_, _36314_, \oc8051_golden_model_1.PSW [7]);
  or (_36501_, _11575_, _07911_);
  and (_36502_, _36501_, _11363_);
  and (_36503_, _36502_, _36500_);
  or (_36504_, _36503_, _36499_);
  and (_36505_, _36504_, _11361_);
  and (_36506_, _36350_, _11877_);
  or (_36508_, _36506_, _11358_);
  or (_36509_, _36508_, _36505_);
  or (_36510_, _11575_, _11357_);
  and (_36511_, _36510_, _04608_);
  and (_36512_, _36511_, _36509_);
  nand (_36513_, _11418_, _03653_);
  nand (_36514_, _36513_, _11890_);
  or (_36515_, _36514_, _36512_);
  nor (_36516_, _11893_, _13020_);
  or (_36517_, _36516_, _24294_);
  and (_36519_, _36517_, _36515_);
  or (_36520_, _36314_, _07911_);
  or (_36521_, _11575_, \oc8051_golden_model_1.PSW [7]);
  and (_36522_, _36521_, _11893_);
  and (_36523_, _36522_, _36520_);
  or (_36524_, _36523_, _36519_);
  and (_36525_, _36524_, _11355_);
  and (_36526_, _36350_, _11898_);
  or (_36527_, _36526_, _08571_);
  or (_36528_, _36527_, _36525_);
  or (_36530_, _11575_, _08570_);
  and (_36531_, _36530_, _08601_);
  and (_36532_, _36531_, _36528_);
  and (_36533_, _36350_, _08600_);
  or (_36534_, _36533_, _36532_);
  and (_36535_, _36534_, _10680_);
  nor (_36536_, _05840_, _10680_);
  or (_36537_, _36536_, _03248_);
  or (_36538_, _36537_, _36535_);
  nand (_36539_, _13020_, _03248_);
  and (_36541_, _36539_, _03796_);
  and (_36542_, _36541_, _36538_);
  and (_36543_, _36322_, _09914_);
  nor (_36544_, _11419_, _09914_);
  or (_36545_, _36544_, _36543_);
  and (_36546_, _36545_, _03652_);
  or (_36547_, _36546_, _36542_);
  and (_36548_, _36547_, _11353_);
  and (_36549_, _36350_, _11919_);
  or (_36550_, _36549_, _08722_);
  or (_36552_, _36550_, _36548_);
  or (_36553_, _11575_, _08721_);
  and (_36554_, _36553_, _08770_);
  and (_36555_, _36554_, _36552_);
  and (_36556_, _36350_, _08769_);
  or (_36557_, _36556_, _03521_);
  or (_36558_, _36557_, _36555_);
  nand (_36559_, _05840_, _03521_);
  and (_36560_, _36559_, _36558_);
  or (_36561_, _36560_, _03246_);
  and (_36563_, _36561_, _36312_);
  or (_36564_, _36563_, _03519_);
  nand (_36565_, _11419_, _09914_);
  or (_36566_, _36322_, _09914_);
  and (_36567_, _36566_, _36565_);
  or (_36568_, _36567_, _03520_);
  and (_36569_, _36568_, _11945_);
  and (_36570_, _36569_, _36564_);
  and (_36571_, _36350_, _11946_);
  or (_36572_, _36571_, _03809_);
  or (_36574_, _36572_, _36570_);
  nand (_36575_, _13020_, _03809_);
  and (_36576_, _36575_, _11952_);
  and (_36577_, _36576_, _36574_);
  and (_36578_, _36350_, _35342_);
  or (_36579_, _36578_, _03686_);
  or (_36580_, _36579_, _36577_);
  nand (_36581_, _04308_, _03686_);
  and (_36582_, _36581_, _12381_);
  and (_36583_, _36582_, _36580_);
  and (_36585_, _11575_, _03243_);
  or (_36586_, _36585_, _03205_);
  or (_36587_, _36586_, _36583_);
  or (_36588_, _36567_, _03206_);
  and (_36589_, _36588_, _11967_);
  and (_36590_, _36589_, _36587_);
  and (_36591_, _36350_, _11968_);
  or (_36592_, _36591_, _03816_);
  or (_36593_, _36592_, _36590_);
  nand (_36594_, _13020_, _03816_);
  and (_36596_, _36594_, _11974_);
  and (_36597_, _36596_, _36593_);
  and (_36598_, _36350_, _33977_);
  or (_36599_, _36598_, _03684_);
  or (_36600_, _36599_, _36597_);
  nand (_36601_, _04308_, _03684_);
  and (_36602_, _36601_, _24650_);
  and (_36603_, _36602_, _36600_);
  and (_36604_, _36350_, _11982_);
  and (_36605_, _11575_, _03242_);
  or (_36607_, _36605_, _36604_);
  or (_36608_, _36607_, _36603_);
  or (_36609_, _36608_, _43231_);
  or (_36610_, _43227_, \oc8051_golden_model_1.PC [12]);
  and (_36611_, _36610_, _41991_);
  and (_43624_, _36611_, _36609_);
  nor (_36612_, _11347_, \oc8051_golden_model_1.PC [13]);
  nor (_36613_, _36612_, _11348_);
  or (_36614_, _36613_, _11353_);
  or (_36615_, _36613_, _11355_);
  or (_36617_, _36613_, _11361_);
  or (_36618_, _36613_, _11370_);
  or (_36619_, _36613_, _11841_);
  and (_36620_, _11413_, _03644_);
  or (_36621_, _36613_, _11381_);
  and (_36622_, _36613_, _11387_);
  or (_36623_, _11416_, _11415_);
  not (_36624_, _36623_);
  nor (_36625_, _36624_, _11514_);
  and (_36626_, _36624_, _11514_);
  or (_36628_, _36626_, _36625_);
  or (_36629_, _36628_, _10133_);
  nand (_36630_, _11414_, _10133_);
  and (_36631_, _36630_, _03676_);
  and (_36632_, _36631_, _36629_);
  nand (_36633_, _11414_, _09946_);
  or (_36634_, _36628_, _09946_);
  and (_36635_, _36634_, _03615_);
  and (_36636_, _36635_, _36633_);
  nand (_36637_, _11414_, _10037_);
  or (_36639_, _36628_, _10037_);
  and (_36640_, _36639_, _11706_);
  and (_36641_, _36640_, _36637_);
  and (_36642_, _11571_, _03603_);
  or (_36643_, _11679_, _11571_);
  or (_36644_, _36628_, _11397_);
  or (_36645_, _11413_, _11526_);
  and (_36646_, _36645_, _03599_);
  and (_36647_, _36646_, _36644_);
  and (_36648_, _11571_, _11554_);
  or (_36650_, _11573_, _11572_);
  not (_36651_, _36650_);
  nor (_36652_, _36651_, _11659_);
  and (_36653_, _36651_, _11659_);
  or (_36654_, _36653_, _36652_);
  and (_36655_, _36654_, _11556_);
  or (_36656_, _36655_, _06054_);
  or (_36657_, _36656_, _36648_);
  or (_36658_, _36613_, _35411_);
  or (_36659_, _11571_, _03948_);
  nor (_36661_, _04499_, \oc8051_golden_model_1.PC [13]);
  nand (_36662_, _36661_, _11531_);
  and (_36663_, _36662_, _36659_);
  or (_36664_, _36663_, _11536_);
  and (_36665_, _36664_, _36658_);
  and (_36666_, _11571_, _03947_);
  and (_36667_, _36613_, _32577_);
  or (_36668_, _36667_, _12226_);
  or (_36669_, _36668_, _36666_);
  or (_36670_, _36669_, _36665_);
  and (_36672_, _36670_, _11674_);
  and (_36673_, _36672_, _36657_);
  or (_36674_, _36673_, _36647_);
  and (_36675_, _36674_, _11391_);
  and (_36676_, _36613_, _35715_);
  or (_36677_, _36676_, _36064_);
  or (_36678_, _36677_, _36675_);
  and (_36679_, _36678_, _36643_);
  or (_36680_, _36679_, _33003_);
  or (_36681_, _36613_, _11684_);
  and (_36683_, _36681_, _03611_);
  and (_36684_, _36683_, _36680_);
  or (_36685_, _36684_, _36642_);
  and (_36686_, _36685_, _11692_);
  and (_36687_, _36613_, _11694_);
  or (_36688_, _36687_, _11699_);
  or (_36689_, _36688_, _36686_);
  or (_36690_, _11698_, _11571_);
  and (_36691_, _36690_, _09988_);
  and (_36692_, _36691_, _36689_);
  or (_36694_, _36692_, _36641_);
  or (_36695_, _36694_, _32559_);
  and (_36696_, _11413_, _10089_);
  and (_36697_, _36628_, _11713_);
  or (_36698_, _36697_, _32558_);
  or (_36699_, _36698_, _36696_);
  and (_36700_, _36699_, _04046_);
  and (_36701_, _36700_, _36695_);
  or (_36702_, _36701_, _36636_);
  and (_36703_, _36702_, _09916_);
  or (_36705_, _36703_, _36632_);
  and (_36706_, _36705_, _11389_);
  nand (_36707_, _36613_, _10096_);
  nand (_36708_, _36707_, _11734_);
  or (_36709_, _36708_, _36706_);
  or (_36710_, _11734_, _11571_);
  and (_36711_, _36710_, _11386_);
  and (_36712_, _36711_, _36709_);
  or (_36713_, _36712_, _36622_);
  and (_36714_, _36713_, _11741_);
  nand (_36716_, _36105_, _11571_);
  nand (_36717_, _36716_, _11381_);
  or (_36718_, _36717_, _36714_);
  and (_36719_, _36718_, _36621_);
  or (_36720_, _36719_, _11380_);
  or (_36721_, _11571_, _11379_);
  and (_36722_, _36721_, _03285_);
  and (_36723_, _36722_, _36720_);
  nand (_36724_, _36613_, _03371_);
  nand (_36725_, _36724_, _11752_);
  or (_36727_, _36725_, _36723_);
  or (_36728_, _11752_, _11571_);
  and (_36729_, _36728_, _08865_);
  and (_36730_, _36729_, _36727_);
  nand (_36731_, _11413_, _03656_);
  nand (_36732_, _36731_, _11759_);
  or (_36733_, _36732_, _36730_);
  or (_36734_, _11571_, _11759_);
  and (_36735_, _36734_, _03275_);
  and (_36736_, _36735_, _36733_);
  or (_36738_, _36736_, _36620_);
  and (_36739_, _36738_, _11767_);
  and (_36740_, _36613_, _11770_);
  or (_36741_, _36740_, _11769_);
  or (_36742_, _36741_, _36739_);
  and (_36743_, _11571_, _11373_);
  or (_36744_, _36743_, _23286_);
  and (_36745_, _36744_, _36742_);
  and (_36746_, _36654_, _11372_);
  or (_36747_, _36746_, _06246_);
  or (_36749_, _36747_, _36745_);
  or (_36750_, _11571_, _05966_);
  and (_36751_, _36750_, _04582_);
  and (_36752_, _36751_, _36749_);
  and (_36753_, _11413_, _03650_);
  or (_36754_, _36753_, _08445_);
  or (_36755_, _36754_, _36752_);
  or (_36756_, _11571_, _08446_);
  and (_36757_, _36756_, _11785_);
  and (_36758_, _36757_, _36755_);
  or (_36760_, _11815_, \oc8051_golden_model_1.DPH [5]);
  nor (_36761_, _11816_, _11785_);
  and (_36762_, _36761_, _36760_);
  or (_36763_, _36762_, _11823_);
  or (_36764_, _36763_, _36758_);
  or (_36765_, _11822_, _11571_);
  and (_36766_, _36765_, _11827_);
  and (_36767_, _36766_, _36764_);
  or (_36768_, _36654_, _08820_);
  or (_36769_, _11571_, _11832_);
  and (_36771_, _36769_, _11826_);
  and (_36772_, _36771_, _36768_);
  or (_36773_, _36772_, _11845_);
  or (_36774_, _36773_, _36767_);
  and (_36775_, _36774_, _36619_);
  or (_36776_, _36775_, _11844_);
  or (_36777_, _11571_, _11843_);
  and (_36778_, _36777_, _04591_);
  and (_36779_, _36778_, _36776_);
  nand (_36780_, _11413_, _03649_);
  nand (_36782_, _36780_, _11853_);
  or (_36783_, _36782_, _36779_);
  or (_36784_, _11853_, _11571_);
  and (_36785_, _36784_, _11857_);
  and (_36786_, _36785_, _36783_);
  or (_36787_, _36654_, _11832_);
  or (_36788_, _11571_, _08820_);
  and (_36789_, _36788_, _11856_);
  and (_36790_, _36789_, _36787_);
  or (_36791_, _36790_, _11865_);
  or (_36793_, _36791_, _36786_);
  and (_36794_, _36793_, _36618_);
  or (_36795_, _36794_, _11368_);
  or (_36796_, _11367_, _11571_);
  and (_36797_, _36796_, _04596_);
  and (_36798_, _36797_, _36795_);
  nand (_36799_, _11413_, _03655_);
  nand (_36800_, _36799_, _10776_);
  or (_36801_, _36800_, _36798_);
  and (_36802_, _11571_, _11364_);
  or (_36804_, _36802_, _24139_);
  and (_36805_, _36804_, _36801_);
  or (_36806_, _36654_, \oc8051_golden_model_1.PSW [7]);
  or (_36807_, _11571_, _07911_);
  and (_36808_, _36807_, _11363_);
  and (_36809_, _36808_, _36806_);
  or (_36810_, _36809_, _11877_);
  or (_36811_, _36810_, _36805_);
  and (_36812_, _36811_, _36617_);
  or (_36813_, _36812_, _11358_);
  or (_36815_, _11571_, _11357_);
  and (_36816_, _36815_, _04608_);
  and (_36817_, _36816_, _36813_);
  nand (_36818_, _11413_, _03653_);
  nand (_36819_, _36818_, _11890_);
  or (_36820_, _36819_, _36817_);
  and (_36821_, _11894_, _11571_);
  or (_36822_, _36821_, _24294_);
  and (_36823_, _36822_, _36820_);
  or (_36824_, _36654_, _07911_);
  or (_36826_, _11571_, \oc8051_golden_model_1.PSW [7]);
  and (_36827_, _36826_, _11893_);
  and (_36828_, _36827_, _36824_);
  or (_36829_, _36828_, _11898_);
  or (_36830_, _36829_, _36823_);
  and (_36831_, _36830_, _36615_);
  or (_36832_, _36831_, _08571_);
  or (_36833_, _11571_, _08570_);
  and (_36834_, _36833_, _08601_);
  and (_36835_, _36834_, _36832_);
  and (_36837_, _36613_, _08600_);
  or (_36838_, _36837_, _03792_);
  or (_36839_, _36838_, _36835_);
  nand (_36840_, _05552_, _03792_);
  and (_36841_, _36840_, _36839_);
  or (_36842_, _36841_, _03248_);
  or (_36843_, _11571_, _06475_);
  and (_36844_, _36843_, _03796_);
  and (_36845_, _36844_, _36842_);
  or (_36846_, _36628_, _11920_);
  or (_36848_, _11413_, _09914_);
  and (_36849_, _36848_, _03652_);
  and (_36850_, _36849_, _36846_);
  or (_36851_, _36850_, _11919_);
  or (_36852_, _36851_, _36845_);
  and (_36853_, _36852_, _36614_);
  or (_36854_, _36853_, _08722_);
  or (_36855_, _11571_, _08721_);
  and (_36856_, _36855_, _08770_);
  and (_36857_, _36856_, _36854_);
  and (_36859_, _36613_, _08769_);
  or (_36860_, _36859_, _03521_);
  or (_36861_, _36860_, _36857_);
  nand (_36862_, _05552_, _03521_);
  and (_36863_, _36862_, _36861_);
  or (_36864_, _36863_, _03246_);
  or (_36865_, _11571_, _32287_);
  and (_36866_, _36865_, _03520_);
  and (_36867_, _36866_, _36864_);
  nand (_36868_, _11414_, _09914_);
  or (_36870_, _36628_, _09914_);
  and (_36871_, _36870_, _36868_);
  and (_36872_, _36871_, _03519_);
  or (_36873_, _36872_, _11946_);
  or (_36874_, _36873_, _36867_);
  or (_36875_, _36613_, _11945_);
  and (_36876_, _36875_, _04260_);
  and (_36877_, _36876_, _36874_);
  nand (_36878_, _11571_, _03809_);
  nand (_36879_, _36878_, _11952_);
  or (_36881_, _36879_, _36877_);
  or (_36882_, _36613_, _11952_);
  and (_36883_, _36882_, _11956_);
  and (_36884_, _36883_, _36881_);
  nor (_36885_, _03853_, _11956_);
  or (_36886_, _36885_, _03243_);
  or (_36887_, _36886_, _36884_);
  or (_36888_, _11571_, _12381_);
  and (_36889_, _36888_, _03206_);
  and (_36890_, _36889_, _36887_);
  and (_36892_, _36871_, _03205_);
  or (_36893_, _36892_, _11968_);
  or (_36894_, _36893_, _36890_);
  or (_36895_, _36613_, _11967_);
  and (_36896_, _36895_, _03820_);
  and (_36897_, _36896_, _36894_);
  nand (_36898_, _11571_, _03816_);
  nand (_36899_, _36898_, _11974_);
  or (_36900_, _36899_, _36897_);
  or (_36901_, _36613_, _11974_);
  and (_36903_, _36901_, _11978_);
  and (_36904_, _36903_, _36900_);
  nor (_36905_, _03853_, _11978_);
  or (_36906_, _36905_, _03242_);
  or (_36907_, _36906_, _36904_);
  or (_36908_, _11571_, _36298_);
  and (_36909_, _36908_, _11990_);
  and (_36910_, _36909_, _36907_);
  and (_36911_, _36613_, _11982_);
  or (_36912_, _36911_, _36910_);
  or (_36914_, _36912_, _43231_);
  or (_36915_, _43227_, \oc8051_golden_model_1.PC [13]);
  and (_36916_, _36915_, _41991_);
  and (_43625_, _36916_, _36914_);
  nor (_36917_, _11348_, \oc8051_golden_model_1.PC [14]);
  nor (_36918_, _36917_, _11349_);
  nor (_36919_, _36918_, _08770_);
  not (_36920_, _11565_);
  nor (_36921_, _11890_, _36920_);
  nor (_36922_, _11406_, _04608_);
  nor (_36924_, _36920_, _10776_);
  nor (_36925_, _11853_, _36920_);
  nor (_36926_, _11406_, _04591_);
  nor (_36927_, _11822_, _36920_);
  nor (_36928_, _11406_, _08865_);
  nor (_36929_, _11565_, _11379_);
  nor (_36930_, _36918_, _11386_);
  nor (_36931_, _36918_, _11389_);
  nor (_36932_, _11698_, _36920_);
  not (_36933_, _36918_);
  nor (_36935_, _36933_, _11692_);
  nor (_36936_, _36918_, _11684_);
  and (_36937_, _11516_, _11411_);
  nor (_36938_, _36937_, _11517_);
  or (_36939_, _36938_, _11397_);
  or (_36940_, _11406_, _11526_);
  and (_36941_, _36940_, _36939_);
  nor (_36942_, _36941_, _04515_);
  and (_36943_, _11661_, _11569_);
  nor (_36944_, _36943_, _11662_);
  nand (_36946_, _36944_, _11556_);
  or (_36947_, _36920_, _11556_);
  and (_36948_, _36947_, _12226_);
  nand (_36949_, _36948_, _36946_);
  nor (_36950_, _11565_, _04868_);
  or (_36951_, _36950_, _32577_);
  nand (_36952_, _36920_, _03946_);
  nor (_36953_, _04499_, \oc8051_golden_model_1.PC [14]);
  nand (_36954_, _36953_, _11531_);
  and (_36955_, _36954_, _36952_);
  or (_36957_, _36955_, _11536_);
  or (_36958_, _36918_, _32309_);
  and (_36959_, _36958_, _36957_);
  nor (_36960_, _36959_, _03947_);
  nor (_36961_, _36960_, _36951_);
  nor (_36962_, _36933_, _11540_);
  nor (_36963_, _36962_, _12226_);
  not (_36964_, _36963_);
  nor (_36965_, _36964_, _36961_);
  nor (_36966_, _36965_, _04509_);
  nand (_36968_, _36966_, _36949_);
  and (_36969_, _36918_, _04509_);
  nor (_36970_, _36969_, _03599_);
  and (_36971_, _36970_, _36968_);
  or (_36972_, _36971_, _36942_);
  nand (_36973_, _36972_, _11391_);
  nor (_36974_, _36918_, _11391_);
  nor (_36975_, _36974_, _36064_);
  and (_36976_, _36975_, _36973_);
  nor (_36977_, _11679_, _36920_);
  nor (_36979_, _36977_, _36976_);
  and (_36980_, _36979_, _11684_);
  or (_36981_, _36980_, _36936_);
  nand (_36982_, _36981_, _03611_);
  nor (_36983_, _11565_, _03611_);
  nor (_36984_, _36983_, _11694_);
  and (_36985_, _36984_, _36982_);
  or (_36986_, _36985_, _36935_);
  and (_36987_, _36986_, _11698_);
  or (_36988_, _36987_, _11706_);
  nor (_36990_, _36988_, _36932_);
  nand (_36991_, _11406_, _10037_);
  not (_36992_, _36938_);
  or (_36993_, _36992_, _10037_);
  and (_36994_, _36993_, _11706_);
  and (_36995_, _36994_, _36991_);
  or (_36996_, _36995_, _36990_);
  or (_36997_, _36996_, _10041_);
  nor (_36998_, _36938_, _10089_);
  and (_36999_, _11407_, _10089_);
  or (_37001_, _36999_, _10042_);
  or (_37002_, _37001_, _36998_);
  and (_37003_, _37002_, _04046_);
  and (_37004_, _37003_, _36997_);
  and (_37005_, _11406_, _09946_);
  nor (_37006_, _36992_, _09946_);
  or (_37007_, _37006_, _04046_);
  nor (_37008_, _37007_, _37005_);
  or (_37009_, _37008_, _03676_);
  or (_37010_, _37009_, _37004_);
  nor (_37012_, _36938_, _10133_);
  and (_37013_, _11407_, _10133_);
  nor (_37014_, _37013_, _09916_);
  not (_37015_, _37014_);
  nor (_37016_, _37015_, _37012_);
  nor (_37017_, _37016_, _10096_);
  nand (_37018_, _37017_, _37010_);
  nand (_37019_, _37018_, _11734_);
  or (_37020_, _37019_, _36931_);
  nor (_37021_, _11734_, _36920_);
  nor (_37023_, _37021_, _11387_);
  and (_37024_, _37023_, _37020_);
  or (_37025_, _37024_, _36930_);
  nand (_37026_, _37025_, _11741_);
  nor (_37027_, _11741_, _11565_);
  nor (_37028_, _37027_, _33065_);
  nand (_37029_, _37028_, _37026_);
  nor (_37030_, _36933_, _11381_);
  nor (_37031_, _37030_, _11380_);
  and (_37032_, _37031_, _37029_);
  or (_37034_, _37032_, _36929_);
  nand (_37035_, _37034_, _03285_);
  nor (_37036_, _36918_, _03285_);
  nor (_37037_, _37036_, _11753_);
  nand (_37038_, _37037_, _37035_);
  nor (_37039_, _11752_, _36920_);
  nor (_37040_, _37039_, _03656_);
  nand (_37041_, _37040_, _37038_);
  nand (_37042_, _37041_, _11759_);
  or (_37043_, _37042_, _36928_);
  nor (_37045_, _36920_, _11759_);
  nor (_37046_, _37045_, _03644_);
  nand (_37047_, _37046_, _37043_);
  nor (_37048_, _11406_, _03275_);
  nor (_37049_, _37048_, _11770_);
  nand (_37050_, _37049_, _37047_);
  nor (_37051_, _36933_, _11767_);
  nor (_37052_, _37051_, _11769_);
  nand (_37053_, _37052_, _37050_);
  nor (_37054_, _11565_, _11374_);
  nor (_37056_, _37054_, _11372_);
  and (_37057_, _37056_, _37053_);
  and (_37058_, _36944_, _11372_);
  nor (_37059_, _37058_, _37057_);
  or (_37060_, _37059_, _06246_);
  or (_37061_, _36920_, _05966_);
  and (_37062_, _37061_, _04582_);
  nand (_37063_, _37062_, _37060_);
  nor (_37064_, _11406_, _04582_);
  nor (_37065_, _37064_, _08445_);
  nand (_37067_, _37065_, _37063_);
  and (_37068_, _11565_, _08445_);
  nor (_37069_, _37068_, _11784_);
  nand (_37070_, _37069_, _37067_);
  nor (_37071_, _11816_, \oc8051_golden_model_1.DPH [6]);
  nor (_37072_, _37071_, _11817_);
  nor (_37073_, _37072_, _11785_);
  nor (_37074_, _37073_, _11823_);
  and (_37075_, _37074_, _37070_);
  or (_37076_, _37075_, _36927_);
  nand (_37078_, _37076_, _11827_);
  and (_37079_, _11565_, _08820_);
  and (_37080_, _36944_, _11832_);
  or (_37081_, _37080_, _37079_);
  and (_37082_, _37081_, _11826_);
  nor (_37083_, _37082_, _11845_);
  nand (_37084_, _37083_, _37078_);
  nor (_37085_, _36918_, _11841_);
  nor (_37086_, _37085_, _11844_);
  nand (_37087_, _37086_, _37084_);
  nor (_37089_, _36920_, _11843_);
  nor (_37090_, _37089_, _03649_);
  nand (_37091_, _37090_, _37087_);
  nand (_37092_, _37091_, _11853_);
  nor (_37093_, _37092_, _36926_);
  or (_37094_, _37093_, _36925_);
  nand (_37095_, _37094_, _11857_);
  nor (_37096_, _36944_, _11832_);
  nor (_37097_, _11565_, _08820_);
  nor (_37098_, _37097_, _11857_);
  not (_37100_, _37098_);
  nor (_37101_, _37100_, _37096_);
  nor (_37102_, _37101_, _11865_);
  nand (_37103_, _37102_, _37095_);
  nor (_37104_, _36918_, _11370_);
  nor (_37105_, _37104_, _11368_);
  nand (_37106_, _37105_, _37103_);
  nor (_37107_, _11367_, _36920_);
  nor (_37108_, _37107_, _03655_);
  nand (_37109_, _37108_, _37106_);
  nor (_37111_, _11406_, _04596_);
  nor (_37112_, _37111_, _10777_);
  and (_37113_, _37112_, _37109_);
  or (_37114_, _37113_, _36924_);
  nand (_37115_, _37114_, _11364_);
  and (_37116_, _11565_, \oc8051_golden_model_1.PSW [7]);
  and (_37117_, _36944_, _07911_);
  or (_37118_, _37117_, _37116_);
  and (_37119_, _37118_, _11363_);
  nor (_37120_, _37119_, _11877_);
  nand (_37122_, _37120_, _37115_);
  nor (_37123_, _36918_, _11361_);
  nor (_37124_, _37123_, _11358_);
  nand (_37125_, _37124_, _37122_);
  nor (_37126_, _36920_, _11357_);
  nor (_37127_, _37126_, _03653_);
  nand (_37128_, _37127_, _37125_);
  nand (_37129_, _37128_, _11890_);
  nor (_37130_, _37129_, _36922_);
  or (_37131_, _37130_, _36921_);
  nand (_37133_, _37131_, _11894_);
  nand (_37134_, _11565_, _07911_);
  nand (_37135_, _36944_, \oc8051_golden_model_1.PSW [7]);
  and (_37136_, _37135_, _37134_);
  or (_37137_, _37136_, _11894_);
  and (_37138_, _37137_, _37133_);
  nand (_37139_, _37138_, _11355_);
  nor (_37140_, _36918_, _11355_);
  nor (_37141_, _37140_, _08571_);
  nand (_37142_, _37141_, _37139_);
  nor (_37144_, _36920_, _08570_);
  nor (_37145_, _37144_, _08600_);
  nand (_37146_, _37145_, _37142_);
  nor (_37147_, _36918_, _08601_);
  nor (_37148_, _37147_, _03792_);
  and (_37149_, _37148_, _37146_);
  nor (_37150_, _05442_, _10680_);
  or (_37151_, _37150_, _03248_);
  or (_37152_, _37151_, _37149_);
  nor (_37153_, _11565_, _06475_);
  nor (_37155_, _37153_, _03652_);
  nand (_37156_, _37155_, _37152_);
  nor (_37157_, _11406_, _09914_);
  and (_37158_, _36992_, _09914_);
  or (_37159_, _37158_, _03796_);
  or (_37160_, _37159_, _37157_);
  and (_37161_, _37160_, _11353_);
  nand (_37162_, _37161_, _37156_);
  nor (_37163_, _36918_, _11353_);
  nor (_37164_, _37163_, _08722_);
  nand (_37166_, _37164_, _37162_);
  nor (_37167_, _36920_, _08721_);
  nor (_37168_, _37167_, _08769_);
  and (_37169_, _37168_, _37166_);
  or (_37170_, _37169_, _36919_);
  nand (_37171_, _37170_, _03522_);
  and (_37172_, _05442_, _03521_);
  nor (_37173_, _37172_, _03246_);
  and (_37174_, _37173_, _37171_);
  and (_37175_, _11565_, _03246_);
  or (_37177_, _37175_, _03519_);
  nor (_37178_, _37177_, _37174_);
  and (_37179_, _11407_, _09914_);
  nor (_37180_, _36938_, _09914_);
  nor (_37181_, _37180_, _37179_);
  nor (_37182_, _37181_, _03520_);
  or (_37183_, _37182_, _37178_);
  and (_37184_, _37183_, _11945_);
  nor (_37185_, _36918_, _11945_);
  or (_37186_, _37185_, _37184_);
  nand (_37188_, _37186_, _04260_);
  and (_37189_, _36920_, _03809_);
  nor (_37190_, _37189_, _35342_);
  nand (_37191_, _37190_, _37188_);
  nor (_37192_, _36933_, _11952_);
  nor (_37193_, _37192_, _03686_);
  nand (_37194_, _37193_, _37191_);
  and (_37195_, _03686_, _03556_);
  nor (_37196_, _37195_, _03243_);
  nand (_37197_, _37196_, _37194_);
  and (_37199_, _11565_, _03243_);
  nor (_37200_, _37199_, _03205_);
  nand (_37201_, _37200_, _37197_);
  nor (_37202_, _37181_, _03206_);
  nor (_37203_, _37202_, _11968_);
  nand (_37204_, _37203_, _37201_);
  nor (_37205_, _36933_, _11967_);
  nor (_37206_, _37205_, _03816_);
  nand (_37207_, _37206_, _37204_);
  and (_37208_, _36920_, _03816_);
  nor (_37210_, _37208_, _33977_);
  nand (_37211_, _37210_, _37207_);
  nor (_37212_, _36933_, _11974_);
  nor (_37213_, _37212_, _03684_);
  nand (_37214_, _37213_, _37211_);
  and (_37215_, _03684_, _03556_);
  nor (_37216_, _37215_, _03242_);
  and (_37217_, _37216_, _37214_);
  and (_37218_, _11565_, _03242_);
  or (_37219_, _37218_, _37217_);
  and (_37221_, _37219_, _11990_);
  and (_37222_, _36918_, _11982_);
  or (_37223_, _37222_, _37221_);
  or (_37224_, _37223_, _43231_);
  or (_37225_, _43227_, \oc8051_golden_model_1.PC [14]);
  and (_37226_, _37225_, _41991_);
  and (_43626_, _37226_, _37224_);
  and (_37227_, _43231_, \oc8051_golden_model_1.P0INREG [0]);
  or (_37228_, _37227_, _01128_);
  and (_43627_, _37228_, _41991_);
  and (_37230_, _43231_, \oc8051_golden_model_1.P0INREG [1]);
  or (_37231_, _37230_, _01135_);
  and (_43628_, _37231_, _41991_);
  and (_37232_, _43231_, \oc8051_golden_model_1.P0INREG [2]);
  or (_37233_, _37232_, _01103_);
  and (_43629_, _37233_, _41991_);
  and (_37234_, _43231_, \oc8051_golden_model_1.P0INREG [3]);
  or (_37235_, _37234_, _01096_);
  and (_43630_, _37235_, _41991_);
  and (_37236_, _43231_, \oc8051_golden_model_1.P0INREG [4]);
  or (_37238_, _37236_, _01144_);
  and (_43631_, _37238_, _41991_);
  and (_37239_, _43231_, \oc8051_golden_model_1.P0INREG [5]);
  or (_37240_, _37239_, _01151_);
  and (_43632_, _37240_, _41991_);
  and (_37241_, _43231_, \oc8051_golden_model_1.P0INREG [6]);
  or (_37242_, _37241_, _01110_);
  and (_43633_, _37242_, _41991_);
  and (_37243_, _43231_, \oc8051_golden_model_1.P1INREG [0]);
  or (_37244_, _37243_, _00919_);
  and (_43636_, _37244_, _41991_);
  and (_37246_, _43231_, \oc8051_golden_model_1.P1INREG [1]);
  or (_37247_, _37246_, _00936_);
  and (_43637_, _37247_, _41991_);
  and (_37248_, _43231_, \oc8051_golden_model_1.P1INREG [2]);
  or (_37249_, _37248_, _00952_);
  and (_43638_, _37249_, _41991_);
  and (_37250_, _43231_, \oc8051_golden_model_1.P1INREG [3]);
  or (_37251_, _37250_, _00928_);
  and (_43639_, _37251_, _41991_);
  and (_37253_, _43231_, \oc8051_golden_model_1.P1INREG [4]);
  or (_37254_, _37253_, _00911_);
  and (_43640_, _37254_, _41991_);
  and (_37255_, _43231_, \oc8051_golden_model_1.P1INREG [5]);
  or (_37256_, _37255_, _00943_);
  and (_43643_, _37256_, _41991_);
  and (_37257_, _43231_, \oc8051_golden_model_1.P1INREG [6]);
  or (_37258_, _37257_, _00959_);
  and (_43644_, _37258_, _41991_);
  and (_37259_, _43231_, \oc8051_golden_model_1.P2INREG [0]);
  or (_37261_, _37259_, _01193_);
  and (_43645_, _37261_, _41991_);
  and (_37262_, _43231_, \oc8051_golden_model_1.P2INREG [1]);
  or (_37263_, _37262_, _01227_);
  and (_43646_, _37263_, _41991_);
  and (_37264_, _43231_, \oc8051_golden_model_1.P2INREG [2]);
  or (_37265_, _37264_, _01211_);
  and (_43647_, _37265_, _41991_);
  and (_37266_, _43231_, \oc8051_golden_model_1.P2INREG [3]);
  or (_37267_, _37266_, _01202_);
  and (_43648_, _37267_, _41991_);
  and (_37269_, _43231_, \oc8051_golden_model_1.P2INREG [4]);
  or (_37270_, _37269_, _01186_);
  and (_43649_, _37270_, _41991_);
  and (_37271_, _43231_, \oc8051_golden_model_1.P2INREG [5]);
  or (_37272_, _37271_, _01234_);
  and (_43650_, _37272_, _41991_);
  and (_37273_, _43231_, \oc8051_golden_model_1.P2INREG [6]);
  or (_37274_, _37273_, _01218_);
  and (_43651_, _37274_, _41991_);
  and (_37276_, _43231_, \oc8051_golden_model_1.P3INREG [0]);
  or (_37277_, _37276_, _01042_);
  and (_43654_, _37277_, _41991_);
  and (_37278_, _43231_, \oc8051_golden_model_1.P3INREG [1]);
  or (_37279_, _37278_, _01076_);
  and (_43655_, _37279_, _41991_);
  and (_37280_, _43231_, \oc8051_golden_model_1.P3INREG [2]);
  or (_37281_, _37280_, _01060_);
  and (_43656_, _37281_, _41991_);
  and (_37282_, _43231_, \oc8051_golden_model_1.P3INREG [3]);
  or (_37284_, _37282_, _01051_);
  and (_43657_, _37284_, _41991_);
  and (_37285_, _43231_, \oc8051_golden_model_1.P3INREG [4]);
  or (_37286_, _37285_, _01035_);
  and (_43658_, _37286_, _41991_);
  and (_37287_, _43231_, \oc8051_golden_model_1.P3INREG [5]);
  or (_37288_, _37287_, _01083_);
  and (_43659_, _37288_, _41991_);
  and (_37289_, _43231_, \oc8051_golden_model_1.P3INREG [6]);
  or (_37290_, _37289_, _01067_);
  and (_43660_, _37290_, _41991_);
  and (_00005_[6], _01068_, _41991_);
  and (_00005_[5], _01084_, _41991_);
  and (_00005_[4], _01036_, _41991_);
  and (_00005_[3], _01052_, _41991_);
  and (_00005_[2], _01061_, _41991_);
  and (_00005_[1], _01077_, _41991_);
  and (_00005_[0], _01043_, _41991_);
  and (_00004_[6], _01219_, _41991_);
  and (_00004_[5], _01235_, _41991_);
  and (_00004_[4], _01187_, _41991_);
  and (_00004_[3], _01203_, _41991_);
  and (_00004_[2], _01212_, _41991_);
  and (_00004_[1], _01228_, _41991_);
  and (_00004_[0], _01194_, _41991_);
  and (_00003_[6], _00960_, _41991_);
  and (_00003_[5], _00944_, _41991_);
  and (_00003_[4], _00912_, _41991_);
  and (_00003_[3], _00929_, _41991_);
  and (_00003_[2], _00953_, _41991_);
  and (_00003_[1], _00937_, _41991_);
  and (_00003_[0], _00920_, _41991_);
  and (_00002_[6], _01111_, _41991_);
  and (_00002_[5], _01152_, _41991_);
  and (_00002_[4], _01145_, _41991_);
  and (_00002_[3], _01097_, _41991_);
  and (_00002_[2], _01104_, _41991_);
  and (_00002_[1], _01136_, _41991_);
  and (_00002_[0], _01129_, _41991_);
  and (_37294_, _27785_, _40731_);
  or (_37296_, _27661_, _40573_);
  nand (_37297_, _27661_, _40573_);
  and (_37298_, _37297_, _37296_);
  nor (_37299_, _27785_, _40731_);
  or (_37300_, _37299_, _37298_);
  or (_37301_, _37300_, _37294_);
  and (_37302_, _28038_, _38651_);
  nor (_37303_, _28038_, _38651_);
  or (_37304_, _37303_, _37302_);
  and (_37305_, _27909_, _38645_);
  nor (_37307_, _27909_, _38645_);
  or (_37308_, _37307_, _37305_);
  or (_37309_, _37308_, _37304_);
  or (_37310_, _37309_, _37301_);
  nor (_37311_, _28304_, _38663_);
  and (_37312_, _28304_, _38663_);
  or (_37313_, _37312_, _37311_);
  and (_37314_, _28171_, _38657_);
  nor (_37315_, _28171_, _38657_);
  or (_37316_, _37315_, _37314_);
  or (_37318_, _37316_, _37313_);
  nor (_37319_, _28439_, _38669_);
  and (_37320_, _28439_, _38669_);
  or (_37321_, _37320_, _37319_);
  and (_37322_, _10818_, _38625_);
  nor (_37323_, _10818_, _38625_);
  or (_37324_, _37323_, _37322_);
  or (_37325_, _37324_, _37321_);
  or (_37326_, _37325_, _37318_);
  or (_37327_, _37326_, _37310_);
  or (_37329_, _10668_, _09262_);
  nor (_37330_, _37329_, _10925_);
  or (_37331_, _29118_, _28888_);
  nor (_37332_, _37331_, _29233_);
  nor (_37333_, _27577_, _27462_);
  not (_37334_, _28773_);
  and (_37335_, _37334_, _28657_);
  and (_37336_, _37335_, _37333_);
  nor (_37337_, _20031_, _19918_);
  nor (_37338_, _27231_, _26999_);
  and (_37340_, _37338_, _37337_);
  and (_37341_, _37340_, _37336_);
  and (_37342_, _37341_, _37332_);
  nor (_37343_, _10560_, _10479_);
  nor (_37344_, _11089_, _11007_);
  and (_37345_, _37344_, _37343_);
  nor (_37346_, _30542_, _29921_);
  nor (_37347_, _31752_, _31147_);
  and (_37348_, _37347_, _37346_);
  or (_37349_, _11372_, _02995_);
  nor (_37351_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_37352_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_37353_, _37352_, _37351_);
  nor (_37354_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor (_37355_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and (_37356_, _37355_, _37354_);
  and (_37357_, _37356_, _37353_);
  nor (_37358_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_37359_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_37360_, _37359_, _37358_);
  nor (_37362_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_37363_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_37364_, _37363_, _37362_);
  and (_37365_, _37364_, _37360_);
  and (_37366_, _37365_, _37357_);
  nor (_37367_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_37368_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_37369_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_37370_, _37369_, _37368_);
  and (_37371_, _37370_, _37367_);
  nor (_37373_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_37374_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_37375_, _37374_, _37373_);
  nor (_37376_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_37377_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_37378_, _37377_, _37376_);
  and (_37379_, _37378_, _37375_);
  and (_37380_, _37379_, _37371_);
  and (_37381_, _37380_, _37366_);
  nor (_37382_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  nor (_37384_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  and (_37385_, _37384_, _37382_);
  nor (_37386_, \oc8051_golden_model_1.TH0 [3], \oc8051_golden_model_1.TH0 [2]);
  nor (_37387_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [1]);
  and (_37388_, _37387_, _37386_);
  and (_37389_, _37388_, _37385_);
  nor (_37390_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_37391_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_37392_, _37391_, _37390_);
  nor (_37393_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_37395_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_37396_, _37395_, _37393_);
  and (_37397_, _37396_, _37392_);
  and (_37398_, _37397_, _37389_);
  nor (_37399_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_37400_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_37401_, _37400_, _37399_);
  nor (_37402_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  nor (_37403_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  and (_37404_, _37403_, _37402_);
  and (_37406_, _37404_, _37401_);
  nor (_37407_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_37408_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_37409_, _37408_, _37407_);
  nor (_37410_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_37411_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_37412_, _37411_, _37410_);
  and (_37413_, _37412_, _37409_);
  and (_37414_, _37413_, _37406_);
  and (_37415_, _37414_, _37398_);
  nor (_37417_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_37418_, _37417_, op0_cnst);
  nor (_37419_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_37420_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_37421_, _37420_, _37419_);
  nor (_37422_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_37423_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_37424_, _37423_, _37422_);
  and (_37425_, _37424_, _37421_);
  and (_37426_, _37425_, _37418_);
  nor (_37428_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_37429_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_37430_, _37429_, _37428_);
  nor (_37431_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_37432_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_37433_, _37432_, _37431_);
  and (_37434_, _37433_, _37430_);
  and (_37435_, \oc8051_golden_model_1.TCON [1], _28443_);
  nor (_37436_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_37437_, _37436_, _37435_);
  nor (_37439_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_37440_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_37441_, _37440_, _37439_);
  and (_37442_, _37441_, _37437_);
  and (_37443_, _37442_, _37434_);
  and (_37444_, _37443_, _37426_);
  and (_37445_, _37444_, _37415_);
  and (_37446_, _37445_, _37381_);
  nand (_37447_, _37446_, _37349_);
  nor (_37448_, _37447_, _25642_);
  nor (_37450_, _29315_, _26250_);
  and (_37451_, _37450_, _37448_);
  nand (_37452_, _37451_, _37348_);
  nor (_37453_, _37452_, _25729_);
  nor (_37454_, _26338_, _25906_);
  and (_37455_, _37454_, _37453_);
  nor (_37456_, _30094_, _30006_);
  nor (_37457_, _30803_, _30717_);
  and (_37458_, _37457_, _37456_);
  nor (_37459_, _26428_, _25818_);
  nor (_37461_, _29488_, _26515_);
  and (_37462_, _37461_, _37459_);
  and (_37463_, _37462_, _37458_);
  and (_37464_, _37463_, _37455_);
  or (_37465_, _31840_, _31234_);
  nor (_37466_, _37465_, _32016_);
  nor (_37467_, _29577_, _29401_);
  nor (_37468_, _30629_, _30182_);
  and (_37469_, _37468_, _37467_);
  and (_37470_, _37469_, _37466_);
  and (_37472_, _37470_, _37464_);
  nor (_37473_, _29753_, _26780_);
  nor (_37474_, _30360_, _29841_);
  and (_37475_, _37474_, _37473_);
  or (_37476_, _31410_, _31323_);
  or (_37477_, _37476_, _31929_);
  nor (_37478_, _37477_, _26080_);
  nor (_37479_, _26693_, _26168_);
  and (_37480_, _37479_, _37478_);
  and (_37481_, _37480_, _37475_);
  and (_37483_, _37481_, _37472_);
  or (_37484_, _31499_, _30890_);
  nor (_37485_, _37484_, _32105_);
  nor (_37486_, _26604_, _25994_);
  nor (_37487_, _30272_, _29667_);
  and (_37488_, _37487_, _37486_);
  and (_37489_, _37488_, _37485_);
  and (_37490_, _37489_, _37483_);
  and (_37491_, _37490_, _37345_);
  not (_37492_, _19344_);
  nor (_37494_, _19572_, _37492_);
  not (_37495_, _26887_);
  nor (_37496_, _27114_, _37495_);
  and (_37497_, _37496_, _37494_);
  nor (_37498_, _11255_, _11172_);
  not (_37499_, _11336_);
  and (_37500_, _18548_, _37499_);
  and (_37501_, _37500_, _37498_);
  and (_37502_, _37501_, _37497_);
  and (_37503_, _37502_, _37491_);
  nor (_37505_, _19236_, _19122_);
  nor (_37506_, _19689_, _19455_);
  and (_37507_, _37506_, _37505_);
  or (_37508_, _32191_, _31671_);
  nor (_37509_, _37508_, _32277_);
  nor (_37510_, _30977_, _30447_);
  nor (_37511_, _31585_, _31064_);
  and (_37512_, _37511_, _37510_);
  nand (_37513_, _37512_, _37509_);
  or (_37514_, _37513_, _28547_);
  nor (_37516_, _37514_, _18660_);
  nor (_37517_, _18893_, _18776_);
  and (_37518_, _37517_, _37516_);
  and (_37519_, _37518_, _37507_);
  and (_37520_, _37519_, _37503_);
  nor (_37521_, _19804_, _19008_);
  nor (_37522_, _29004_, _27348_);
  nand (_37523_, _37522_, _37521_);
  nor (_37524_, _37523_, _09155_);
  and (_37525_, _37524_, _37520_);
  and (_37527_, _37525_, _37342_);
  and (_37528_, _37527_, _37330_);
  and (_37529_, _37528_, _43227_);
  and (_37530_, _37529_, _41991_);
  and (_00007_, _37530_, _37327_);
  or (_37531_, _25029_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_37532_, _25029_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_37533_, _37532_, _37531_);
  or (_37534_, _25559_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_37535_, _25559_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_37537_, _37535_, _37534_);
  nor (_37538_, _24789_, _39047_);
  and (_37539_, _24789_, _39047_);
  or (_37540_, _37539_, _37538_);
  nor (_37541_, _25143_, _40431_);
  and (_37542_, _25143_, _40431_);
  or (_37543_, _37542_, _37541_);
  or (_37544_, _37543_, _37540_);
  and (_37545_, _25261_, _39132_);
  nor (_37546_, _25261_, _39132_);
  not (_37548_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_37549_, _25376_, _37548_);
  and (_37550_, _25376_, _37548_);
  or (_37551_, _37550_, _37549_);
  or (_37552_, _37551_, _37546_);
  or (_37553_, _37552_, _37545_);
  or (_37554_, _37553_, _37544_);
  or (_37555_, _37554_, _37537_);
  or (_37556_, _37555_, _37533_);
  and (_37557_, _10397_, _39018_);
  nor (_37559_, _10397_, _39018_);
  or (_37560_, _37559_, _37557_);
  or (_37561_, _37560_, _37556_);
  and (_00006_, _37561_, _37530_);
  or (_00001_, _37528_, rst);
  and (_00005_[7], _01029_, _41991_);
  and (_00004_[7], _01180_, _41991_);
  and (_00003_[7], _00969_, _41991_);
  and (_00002_[7], _01120_, _41991_);
  and (_37562_, _37528_, inst_finished_r);
  and (_37564_, _37562_, property_invalid_sp_1_r);
  and (property_invalid_sp, _37564_, _37327_);
  and (_37565_, _25149_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_37566_, \oc8051_golden_model_1.PSW [4], _39132_);
  or (_37567_, _37566_, _37565_);
  and (_37568_, _04957_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_37569_, \oc8051_golden_model_1.PSW [3], _40431_);
  or (_37570_, _37569_, _37568_);
  or (_37571_, _37570_, _37567_);
  and (_37572_, _24681_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_37574_, \oc8051_golden_model_1.PSW [1], _39047_);
  or (_37575_, _37574_, _37572_);
  nand (_37576_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_37577_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_37578_, _37577_, _37576_);
  or (_37579_, _37578_, _37575_);
  or (_37580_, _37579_, _37571_);
  and (_37581_, _07911_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_37582_, \oc8051_golden_model_1.PSW [7], _39018_);
  or (_37583_, _37582_, _37581_);
  and (_37585_, _25266_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_37586_, \oc8051_golden_model_1.PSW [5], _37548_);
  or (_37587_, _37586_, _37585_);
  nand (_37588_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_37589_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_37590_, _37589_, _37588_);
  or (_37591_, _37590_, _37587_);
  or (_37592_, _37591_, _37583_);
  or (_37593_, _37592_, _37580_);
  and (_37594_, _37593_, property_invalid_psw_1_r);
  and (property_invalid_psw, _37594_, _37562_);
  nand (_37596_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_37597_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_37598_, _37597_, _37596_);
  and (_37599_, _22664_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_37600_, \oc8051_golden_model_1.P3 [2], _39879_);
  or (_37601_, _37600_, _37599_);
  or (_37602_, _37601_, _37598_);
  and (_37603_, \oc8051_golden_model_1.P3 [0], _39853_);
  and (_37604_, _22448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_37606_, _37604_, _37603_);
  and (_37607_, _22552_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_37608_, \oc8051_golden_model_1.P3 [1], _39866_);
  or (_37609_, _37608_, _37607_);
  or (_37610_, _37609_, _37606_);
  or (_37611_, _37610_, _37602_);
  or (_37612_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_37613_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_37614_, _37613_, _37612_);
  or (_37615_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_37617_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_37618_, _37617_, _37615_);
  or (_37619_, _37618_, _37614_);
  and (_37620_, _09588_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_37621_, \oc8051_golden_model_1.P3 [7], _39372_);
  or (_37622_, _37621_, _37620_);
  nand (_37623_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_37624_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_37625_, _37624_, _37623_);
  or (_37626_, _37625_, _37622_);
  or (_37628_, _37626_, _37619_);
  or (_37629_, _37628_, _37611_);
  and (property_invalid_p3, _37629_, _37562_);
  nand (_37630_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_37631_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_37632_, _37631_, _37630_);
  and (_37633_, _21892_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_37634_, \oc8051_golden_model_1.P2 [2], _39786_);
  or (_37635_, _37634_, _37633_);
  or (_37636_, _37635_, _37632_);
  and (_37638_, \oc8051_golden_model_1.P2 [0], _39760_);
  and (_37639_, _21676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_37640_, _37639_, _37638_);
  and (_37641_, _21781_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_37642_, \oc8051_golden_model_1.P2 [1], _39773_);
  or (_37643_, _37642_, _37641_);
  or (_37644_, _37643_, _37640_);
  or (_37645_, _37644_, _37636_);
  or (_37646_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_37647_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_37649_, _37647_, _37646_);
  or (_37650_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_37651_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_37652_, _37651_, _37650_);
  or (_37653_, _37652_, _37649_);
  and (_37654_, _09484_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_37655_, \oc8051_golden_model_1.P2 [7], _39354_);
  or (_37656_, _37655_, _37654_);
  nand (_37657_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_37658_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_37660_, _37658_, _37657_);
  or (_37661_, _37660_, _37656_);
  or (_37662_, _37661_, _37653_);
  or (_37663_, _37662_, _37645_);
  and (property_invalid_p2, _37663_, _37562_);
  nand (_37664_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_37665_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_37666_, _37665_, _37664_);
  and (_37667_, _21116_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_37668_, \oc8051_golden_model_1.P1 [2], _39699_);
  or (_37670_, _37668_, _37667_);
  or (_37671_, _37670_, _37666_);
  and (_37672_, \oc8051_golden_model_1.P1 [0], _39673_);
  and (_37673_, _20906_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_37674_, _37673_, _37672_);
  and (_37675_, _21007_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_37676_, \oc8051_golden_model_1.P1 [1], _39686_);
  or (_37677_, _37676_, _37675_);
  or (_37678_, _37677_, _37674_);
  or (_37679_, _37678_, _37671_);
  or (_37681_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_37682_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_37683_, _37682_, _37681_);
  or (_37684_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_37685_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_37686_, _37685_, _37684_);
  or (_37687_, _37686_, _37683_);
  and (_37688_, _09382_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_37689_, \oc8051_golden_model_1.P1 [7], _39336_);
  or (_37690_, _37689_, _37688_);
  nand (_37692_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_37693_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_37694_, _37693_, _37692_);
  or (_37695_, _37694_, _37690_);
  or (_37696_, _37695_, _37687_);
  or (_37697_, _37696_, _37679_);
  and (property_invalid_p1, _37697_, _37562_);
  nand (_37698_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_37699_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_37700_, _37699_, _37698_);
  and (_37702_, _20290_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_37703_, \oc8051_golden_model_1.P0 [2], _39610_);
  or (_37704_, _37703_, _37702_);
  or (_37705_, _37704_, _37700_);
  and (_37706_, \oc8051_golden_model_1.P0 [0], _39419_);
  and (_37707_, _20036_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_37708_, _37707_, _37706_);
  and (_37709_, _20163_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_37710_, \oc8051_golden_model_1.P0 [1], _39594_);
  or (_37711_, _37710_, _37709_);
  or (_37713_, _37711_, _37708_);
  or (_37714_, _37713_, _37705_);
  or (_37715_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_37716_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_37717_, _37716_, _37715_);
  or (_37718_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_37719_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_37720_, _37719_, _37718_);
  or (_37721_, _37720_, _37717_);
  and (_37722_, _09266_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_37724_, \oc8051_golden_model_1.P0 [7], _39322_);
  or (_37725_, _37724_, _37722_);
  nand (_37726_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_37727_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_37728_, _37727_, _37726_);
  or (_37729_, _37728_, _37725_);
  or (_37730_, _37729_, _37721_);
  or (_37731_, _37730_, _37714_);
  and (property_invalid_p0, _37731_, _37562_);
  not (_37732_, word_in[1]);
  and (_37734_, _37732_, word_in[0]);
  and (_37735_, _37734_, \oc8051_golden_model_1.IRAM[1] [1]);
  nor (_37736_, _37732_, word_in[0]);
  and (_37737_, _37736_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor (_37738_, _37737_, _37735_);
  nor (_37739_, word_in[1], word_in[0]);
  and (_37740_, _37739_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_37741_, word_in[1], word_in[0]);
  and (_37742_, _37741_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor (_37743_, _37742_, _37740_);
  and (_37745_, _37743_, _37738_);
  nor (_37746_, word_in[3], word_in[2]);
  not (_37747_, _37746_);
  nor (_37748_, _37747_, _37745_);
  and (_37749_, _37734_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_37750_, _37736_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor (_37751_, _37750_, _37749_);
  and (_37752_, _37739_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_37753_, _37741_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_37754_, _37753_, _37752_);
  and (_37756_, _37754_, _37751_);
  and (_37757_, word_in[3], word_in[2]);
  not (_37758_, _37757_);
  nor (_37759_, _37758_, _37756_);
  nor (_37760_, _37759_, _37748_);
  and (_37761_, _37734_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_37762_, _37736_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor (_37763_, _37762_, _37761_);
  and (_37764_, _37739_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_37765_, _37741_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_37767_, _37765_, _37764_);
  and (_37768_, _37767_, _37763_);
  not (_37769_, word_in[3]);
  and (_37770_, _37769_, word_in[2]);
  not (_37771_, _37770_);
  nor (_37772_, _37771_, _37768_);
  and (_37773_, _37734_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_37774_, _37736_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor (_37775_, _37774_, _37773_);
  and (_37776_, _37739_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_37778_, _37741_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor (_37779_, _37778_, _37776_);
  and (_37780_, _37779_, _37775_);
  nor (_37781_, _37769_, word_in[2]);
  not (_37782_, _37781_);
  nor (_37783_, _37782_, _37780_);
  nor (_37784_, _37783_, _37772_);
  and (_37785_, _37784_, _37760_);
  and (_37786_, _37781_, _37741_);
  and (_37787_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_37789_, _37746_, _37739_);
  and (_37790_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_37791_, _37790_, _37787_);
  and (_37792_, _37757_, _37741_);
  and (_37793_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_37794_, _37770_, _37736_);
  and (_37795_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_37796_, _37795_, _37793_);
  and (_37797_, _37796_, _37791_);
  and (_37798_, _37781_, _37736_);
  and (_37800_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_37801_, _37781_, _37734_);
  and (_37802_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_37803_, _37802_, _37800_);
  and (_37804_, _37757_, _37736_);
  and (_37805_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_37806_, _37746_, _37736_);
  and (_37807_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_37808_, _37807_, _37805_);
  and (_37809_, _37808_, _37803_);
  and (_37811_, _37809_, _37797_);
  and (_37812_, _37770_, _37734_);
  and (_37813_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_37814_, _37746_, _37734_);
  and (_37815_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37816_, _37815_, _37813_);
  and (_37817_, _37770_, _37741_);
  and (_37818_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37819_, _37770_, _37739_);
  and (_37820_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_37822_, _37820_, _37818_);
  and (_37823_, _37822_, _37816_);
  and (_37824_, _37781_, _37739_);
  and (_37825_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_37826_, _37746_, _37741_);
  and (_37827_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_37828_, _37827_, _37825_);
  and (_37829_, _37757_, _37734_);
  and (_37830_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_37831_, _37757_, _37739_);
  and (_37833_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_37834_, _37833_, _37830_);
  and (_37835_, _37834_, _37828_);
  and (_37836_, _37835_, _37823_);
  and (_37837_, _37836_, _37811_);
  nand (_37838_, _37837_, _37785_);
  or (_37839_, _37837_, _37785_);
  and (_37840_, _37839_, _37838_);
  and (_37841_, _37734_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_37842_, _37736_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_37844_, _37842_, _37841_);
  and (_37845_, _37739_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_37846_, _37741_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor (_37847_, _37846_, _37845_);
  and (_37848_, _37847_, _37844_);
  nor (_37849_, _37848_, _37747_);
  and (_37850_, _37734_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_37851_, _37736_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor (_37852_, _37851_, _37850_);
  and (_37853_, _37739_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_37855_, _37741_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor (_37856_, _37855_, _37853_);
  and (_37857_, _37856_, _37852_);
  nor (_37858_, _37857_, _37782_);
  nor (_37859_, _37858_, _37849_);
  and (_37860_, _37734_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_37861_, _37736_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_37862_, _37861_, _37860_);
  and (_37863_, _37739_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_37864_, _37741_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor (_37866_, _37864_, _37863_);
  and (_37867_, _37866_, _37862_);
  nor (_37868_, _37867_, _37771_);
  and (_37869_, _37734_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_37870_, _37736_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor (_37871_, _37870_, _37869_);
  and (_37872_, _37739_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_37873_, _37741_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_37874_, _37873_, _37872_);
  and (_37875_, _37874_, _37871_);
  nor (_37877_, _37875_, _37758_);
  nor (_37878_, _37877_, _37868_);
  and (_37879_, _37878_, _37859_);
  and (_37880_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_37881_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37882_, _37881_, _37880_);
  and (_37883_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_37884_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_37885_, _37884_, _37883_);
  and (_37886_, _37885_, _37882_);
  and (_37888_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_37889_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_37890_, _37889_, _37888_);
  and (_37891_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_37892_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_37893_, _37892_, _37891_);
  and (_37894_, _37893_, _37890_);
  and (_37895_, _37894_, _37886_);
  and (_37896_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_37897_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_37899_, _37897_, _37896_);
  and (_37900_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_37901_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_37902_, _37901_, _37900_);
  and (_37903_, _37902_, _37899_);
  and (_37904_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_37905_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_37906_, _37905_, _37904_);
  and (_37907_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_37908_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_37910_, _37908_, _37907_);
  and (_37911_, _37910_, _37906_);
  and (_37912_, _37911_, _37903_);
  and (_37913_, _37912_, _37895_);
  nand (_37914_, _37913_, _37879_);
  or (_37915_, _37913_, _37879_);
  and (_37916_, _37915_, _37914_);
  or (_37917_, _37916_, _37840_);
  and (_37918_, _37734_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_37919_, _37736_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor (_37921_, _37919_, _37918_);
  and (_37922_, _37739_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_37923_, _37741_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor (_37924_, _37923_, _37922_);
  and (_37925_, _37924_, _37921_);
  nor (_37926_, _37925_, _37747_);
  and (_37927_, _37734_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_37928_, _37736_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor (_37929_, _37928_, _37927_);
  and (_37930_, _37739_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_37932_, _37741_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_37933_, _37932_, _37930_);
  and (_37934_, _37933_, _37929_);
  nor (_37935_, _37934_, _37782_);
  nor (_37936_, _37935_, _37926_);
  and (_37937_, _37734_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_37938_, _37736_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_37939_, _37938_, _37937_);
  and (_37940_, _37739_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_37941_, _37741_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor (_37943_, _37941_, _37940_);
  and (_37944_, _37943_, _37939_);
  nor (_37945_, _37944_, _37771_);
  and (_37946_, _37734_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_37947_, _37736_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor (_37948_, _37947_, _37946_);
  and (_37949_, _37739_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_37950_, _37741_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_37951_, _37950_, _37949_);
  and (_37952_, _37951_, _37948_);
  nor (_37954_, _37952_, _37758_);
  nor (_37955_, _37954_, _37945_);
  and (_37956_, _37955_, _37936_);
  and (_37957_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_37958_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_37959_, _37958_, _37957_);
  and (_37960_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_37961_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_37962_, _37961_, _37960_);
  and (_37963_, _37962_, _37959_);
  and (_37965_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_37966_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_37967_, _37966_, _37965_);
  and (_37968_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_37969_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_37970_, _37969_, _37968_);
  and (_37971_, _37970_, _37967_);
  and (_37972_, _37971_, _37963_);
  and (_37973_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_37974_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37976_, _37974_, _37973_);
  and (_37977_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_37978_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_37979_, _37978_, _37977_);
  and (_37980_, _37979_, _37976_);
  and (_37981_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_37982_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_37983_, _37982_, _37981_);
  and (_37984_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_37985_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_37987_, _37985_, _37984_);
  and (_37988_, _37987_, _37983_);
  and (_37989_, _37988_, _37980_);
  and (_37990_, _37989_, _37972_);
  or (_37991_, _37990_, _37956_);
  nand (_37992_, _37990_, _37956_);
  and (_37993_, _37992_, _37991_);
  and (_37994_, _37734_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_37995_, _37736_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor (_37996_, _37995_, _37994_);
  and (_37997_, _37739_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_37998_, _37741_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_37999_, _37998_, _37997_);
  and (_38000_, _37999_, _37996_);
  nor (_38001_, _38000_, _37771_);
  and (_38002_, _37734_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_38003_, _37736_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor (_38004_, _38003_, _38002_);
  and (_38005_, _37739_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_38006_, _37741_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor (_38008_, _38006_, _38005_);
  and (_38009_, _38008_, _38004_);
  nor (_38010_, _38009_, _37782_);
  nor (_38011_, _38010_, _38001_);
  and (_38012_, _37734_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_38013_, _37736_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor (_38014_, _38013_, _38012_);
  and (_38015_, _37739_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_38016_, _37741_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor (_38017_, _38016_, _38015_);
  and (_38019_, _38017_, _38014_);
  nor (_38020_, _38019_, _37747_);
  and (_38021_, _37734_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_38022_, _37736_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_38023_, _38022_, _38021_);
  and (_38024_, _37739_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_38025_, _37741_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_38026_, _38025_, _38024_);
  and (_38027_, _38026_, _38023_);
  nor (_38028_, _38027_, _37758_);
  nor (_38030_, _38028_, _38020_);
  and (_38031_, _38030_, _38011_);
  not (_38032_, _38031_);
  and (_38033_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_38034_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_38035_, _38034_, _38033_);
  and (_38036_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_38037_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_38038_, _38037_, _38036_);
  and (_38039_, _38038_, _38035_);
  and (_38041_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_38042_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_38043_, _38042_, _38041_);
  and (_38044_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_38045_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_38046_, _38045_, _38044_);
  and (_38047_, _38046_, _38043_);
  and (_38048_, _38047_, _38039_);
  and (_38049_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_38050_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_38052_, _38050_, _38049_);
  and (_38053_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_38054_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_38055_, _38054_, _38053_);
  and (_38056_, _38055_, _38052_);
  and (_38057_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_38058_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_38059_, _38058_, _38057_);
  and (_38060_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_38061_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_38063_, _38061_, _38060_);
  and (_38064_, _38063_, _38059_);
  and (_38065_, _38064_, _38056_);
  and (_38066_, _38065_, _38048_);
  nor (_38067_, _38066_, _38032_);
  and (_38068_, _38066_, _38032_);
  or (_38069_, _38068_, _38067_);
  or (_38070_, _38069_, _37993_);
  or (_38071_, _38070_, _37917_);
  and (_38072_, _37734_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_38074_, _37736_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_38075_, _38074_, _38072_);
  and (_38076_, _37739_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_38077_, _37741_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor (_38078_, _38077_, _38076_);
  and (_38079_, _38078_, _38075_);
  nor (_38080_, _38079_, _37771_);
  and (_38081_, _37734_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_38082_, _37736_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_38083_, _38082_, _38081_);
  and (_38085_, _37739_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_38086_, _37741_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_38087_, _38086_, _38085_);
  and (_38088_, _38087_, _38083_);
  nor (_38089_, _38088_, _37758_);
  nor (_38090_, _38089_, _38080_);
  and (_38091_, _37734_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_38092_, _37736_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor (_38093_, _38092_, _38091_);
  and (_38094_, _37739_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_38096_, _37741_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor (_38097_, _38096_, _38094_);
  and (_38098_, _38097_, _38093_);
  nor (_38099_, _38098_, _37747_);
  and (_38100_, _37734_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_38101_, _37736_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor (_38102_, _38101_, _38100_);
  and (_38103_, _37739_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_38104_, _37741_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor (_38105_, _38104_, _38103_);
  and (_38107_, _38105_, _38102_);
  nor (_38108_, _38107_, _37782_);
  nor (_38109_, _38108_, _38099_);
  and (_38110_, _38109_, _38090_);
  and (_38111_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_38112_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_38113_, _38112_, _38111_);
  and (_38114_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_38115_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_38116_, _38115_, _38114_);
  and (_38118_, _38116_, _38113_);
  and (_38119_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_38120_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_38121_, _38120_, _38119_);
  and (_38122_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_38123_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_38124_, _38123_, _38122_);
  and (_38125_, _38124_, _38121_);
  and (_38126_, _38125_, _38118_);
  and (_38127_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_38129_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_38130_, _38129_, _38127_);
  and (_38131_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_38132_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_38133_, _38132_, _38131_);
  and (_38134_, _38133_, _38130_);
  and (_38135_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_38136_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_38137_, _38136_, _38135_);
  and (_38138_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_38140_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_38141_, _38140_, _38138_);
  and (_38142_, _38141_, _38137_);
  and (_38143_, _38142_, _38134_);
  and (_38144_, _38143_, _38126_);
  nand (_38145_, _38144_, _38110_);
  or (_38146_, _38144_, _38110_);
  and (_38147_, _38146_, _38145_);
  and (_38148_, _37734_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_38149_, _37736_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor (_38151_, _38149_, _38148_);
  and (_38152_, _37739_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_38153_, _37741_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor (_38154_, _38153_, _38152_);
  and (_38155_, _38154_, _38151_);
  nor (_38156_, _38155_, _37771_);
  and (_38157_, _37734_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_38158_, _37736_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor (_38159_, _38158_, _38157_);
  and (_38160_, _37739_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_38162_, _37741_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor (_38163_, _38162_, _38160_);
  and (_38164_, _38163_, _38159_);
  nor (_38165_, _38164_, _37782_);
  nor (_38166_, _38165_, _38156_);
  and (_38167_, _37734_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_38168_, _37736_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor (_38169_, _38168_, _38167_);
  and (_38170_, _37739_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_38171_, _37741_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor (_38173_, _38171_, _38170_);
  and (_38174_, _38173_, _38169_);
  nor (_38175_, _38174_, _37747_);
  and (_38176_, _37734_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_38177_, _37736_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_38178_, _38177_, _38176_);
  and (_38179_, _37739_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_38180_, _37741_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_38181_, _38180_, _38179_);
  and (_38182_, _38181_, _38178_);
  nor (_38184_, _38182_, _37758_);
  nor (_38185_, _38184_, _38175_);
  and (_38186_, _38185_, _38166_);
  and (_38187_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_38188_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_38189_, _38188_, _38187_);
  and (_38190_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_38191_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_38192_, _38191_, _38190_);
  and (_38193_, _38192_, _38189_);
  and (_38195_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_38196_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_38197_, _38196_, _38195_);
  and (_38198_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_38199_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_38200_, _38199_, _38198_);
  and (_38201_, _38200_, _38197_);
  and (_38202_, _38201_, _38193_);
  and (_38203_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_38204_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_38206_, _38204_, _38203_);
  and (_38207_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_38208_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_38209_, _38208_, _38207_);
  and (_38210_, _38209_, _38206_);
  and (_38211_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_38212_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_38213_, _38212_, _38211_);
  and (_38214_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_38215_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_38217_, _38215_, _38214_);
  and (_38218_, _38217_, _38213_);
  and (_38219_, _38218_, _38210_);
  and (_38220_, _38219_, _38202_);
  nand (_38221_, _38220_, _38186_);
  or (_38222_, _38220_, _38186_);
  and (_38223_, _38222_, _38221_);
  or (_38224_, _38223_, _38147_);
  and (_38225_, _37734_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_38226_, _37736_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor (_38228_, _38226_, _38225_);
  and (_38229_, _37739_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_38230_, _37741_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor (_38231_, _38230_, _38229_);
  and (_38232_, _38231_, _38228_);
  nor (_38233_, _38232_, _37771_);
  and (_38234_, _37734_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_38235_, _37736_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_38236_, _38235_, _38234_);
  and (_38237_, _37739_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_38239_, _37741_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor (_38240_, _38239_, _38237_);
  and (_38241_, _38240_, _38236_);
  nor (_38242_, _38241_, _37758_);
  nor (_38243_, _38242_, _38233_);
  and (_38244_, _37734_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_38245_, _37736_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor (_38246_, _38245_, _38244_);
  and (_38247_, _37739_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_38248_, _37741_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor (_38250_, _38248_, _38247_);
  and (_38251_, _38250_, _38246_);
  nor (_38252_, _38251_, _37747_);
  and (_38253_, _37734_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_38254_, _37736_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor (_38255_, _38254_, _38253_);
  and (_38256_, _37739_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_38257_, _37741_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_38258_, _38257_, _38256_);
  and (_38259_, _38258_, _38255_);
  nor (_38261_, _38259_, _37782_);
  nor (_38262_, _38261_, _38252_);
  and (_38263_, _38262_, _38243_);
  and (_38264_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_38265_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_38266_, _38265_, _38264_);
  and (_38267_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_38268_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_38269_, _38268_, _38267_);
  and (_38270_, _38269_, _38266_);
  and (_38272_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_38273_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_38274_, _38273_, _38272_);
  and (_38275_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_38276_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_38277_, _38276_, _38275_);
  and (_38278_, _38277_, _38274_);
  and (_38279_, _38278_, _38270_);
  and (_38280_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_38281_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_38283_, _38281_, _38280_);
  and (_38284_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_38285_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_38286_, _38285_, _38284_);
  and (_38287_, _38286_, _38283_);
  and (_38288_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_38289_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_38290_, _38289_, _38288_);
  and (_38291_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_38292_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_38294_, _38292_, _38291_);
  and (_38295_, _38294_, _38290_);
  and (_38296_, _38295_, _38287_);
  and (_38297_, _38296_, _38279_);
  or (_38298_, _38297_, _38263_);
  nand (_38299_, _38297_, _38263_);
  and (_38300_, _38299_, _38298_);
  and (_38301_, _37734_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_38302_, _37736_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor (_38303_, _38302_, _38301_);
  and (_38305_, _37739_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_38306_, _37741_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor (_38307_, _38306_, _38305_);
  and (_38308_, _38307_, _38303_);
  nor (_38309_, _38308_, _37771_);
  and (_38310_, _37734_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_38311_, _37736_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_38312_, _38311_, _38310_);
  and (_38313_, _37739_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_38314_, _37741_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_38316_, _38314_, _38313_);
  and (_38317_, _38316_, _38312_);
  nor (_38318_, _38317_, _37782_);
  nor (_38319_, _38318_, _38309_);
  and (_38320_, _37734_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_38321_, _37736_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor (_38322_, _38321_, _38320_);
  and (_38323_, _37739_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_38324_, _37741_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor (_38325_, _38324_, _38323_);
  and (_38327_, _38325_, _38322_);
  nor (_38328_, _38327_, _37747_);
  and (_38329_, _37734_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_38330_, _37736_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_38331_, _38330_, _38329_);
  and (_38332_, _37739_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_38333_, _37741_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_38334_, _38333_, _38332_);
  and (_38335_, _38334_, _38331_);
  nor (_38336_, _38335_, _37758_);
  nor (_38338_, _38336_, _38328_);
  and (_38339_, _38338_, _38319_);
  and (_38340_, _37794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_38341_, _37812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_38342_, _38341_, _38340_);
  and (_38343_, _37792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_38344_, _37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_38345_, _38344_, _38343_);
  and (_38346_, _38345_, _38342_);
  and (_38347_, _37804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_38349_, _37829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_38350_, _38349_, _38347_);
  and (_38351_, _37798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_38352_, _37801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_38353_, _38352_, _38351_);
  and (_38354_, _38353_, _38350_);
  and (_38355_, _38354_, _38346_);
  and (_38356_, _37789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_38357_, _37806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_38358_, _38357_, _38356_);
  and (_38360_, _37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_38361_, _37819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_38362_, _38361_, _38360_);
  and (_38363_, _38362_, _38358_);
  and (_38364_, _37831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_38365_, _37824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_38366_, _38365_, _38364_);
  and (_38367_, _37826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_38368_, _37814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_38369_, _38368_, _38367_);
  and (_38371_, _38369_, _38366_);
  and (_38372_, _38371_, _38363_);
  and (_38373_, _38372_, _38355_);
  not (_38374_, _38373_);
  nor (_38375_, _38374_, _38339_);
  and (_38376_, _38374_, _38339_);
  or (_38377_, _38376_, _38375_);
  or (_38378_, _38377_, _38300_);
  or (_38379_, _38378_, _38224_);
  or (_38380_, _38379_, _38071_);
  and (property_invalid_iram, _38380_, _37562_);
  nand (_38382_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_38383_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_38384_, _38383_, _38382_);
  and (_38385_, _17978_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_38386_, _17978_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_38387_, _38386_, _38385_);
  or (_38388_, _38387_, _38384_);
  nor (_38389_, _17794_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_38390_, _17794_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_38392_, _38390_, _38389_);
  and (_38393_, _17884_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_38394_, _17884_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_38395_, _38394_, _38393_);
  or (_38396_, _38395_, _38392_);
  or (_38397_, _38396_, _38388_);
  or (_38398_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_38399_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_38400_, _38399_, _38398_);
  or (_38401_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_38403_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_38404_, _38403_, _38401_);
  or (_38405_, _38404_, _38400_);
  and (_38406_, _08955_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_38407_, _08955_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_38408_, _38407_, _38406_);
  nand (_38409_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_38410_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_38411_, _38410_, _38409_);
  or (_38412_, _38411_, _38408_);
  or (_38414_, _38412_, _38405_);
  or (_38415_, _38414_, _38397_);
  and (property_invalid_dph, _38415_, _37562_);
  nand (_38416_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_38417_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38418_, _38417_, _38416_);
  and (_38419_, _17326_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38420_, \oc8051_golden_model_1.DPL [2], _38979_);
  or (_38421_, _38420_, _38419_);
  or (_38422_, _38421_, _38418_);
  and (_38424_, \oc8051_golden_model_1.DPL [0], _38971_);
  and (_38425_, _17143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_38426_, _38425_, _38424_);
  and (_38427_, _17231_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38428_, \oc8051_golden_model_1.DPL [1], _38975_);
  or (_38429_, _38428_, _38427_);
  or (_38430_, _38429_, _38426_);
  or (_38431_, _38430_, _38422_);
  or (_38432_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_38433_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38435_, _38433_, _38432_);
  or (_38436_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_38437_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38438_, _38437_, _38436_);
  or (_38439_, _38438_, _38435_);
  and (_38440_, _08854_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38441_, \oc8051_golden_model_1.DPL [7], _38768_);
  or (_38442_, _38441_, _38440_);
  nand (_38443_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_38444_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38446_, _38444_, _38443_);
  or (_38447_, _38446_, _38442_);
  or (_38448_, _38447_, _38439_);
  or (_38449_, _38448_, _38431_);
  and (property_invalid_dpl, _38449_, _37562_);
  nand (_38450_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_38451_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_38452_, _38451_, _38450_);
  and (_38453_, _07475_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_38454_, \oc8051_golden_model_1.B [2], _30611_);
  or (_38456_, _38454_, _38453_);
  or (_38457_, _38456_, _38452_);
  and (_38458_, \oc8051_golden_model_1.B [0], _29253_);
  and (_38459_, _07467_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_38460_, _38459_, _38458_);
  and (_38461_, _07461_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_38462_, \oc8051_golden_model_1.B [1], _29926_);
  or (_38463_, _38462_, _38461_);
  or (_38464_, _38463_, _38460_);
  or (_38465_, _38464_, _38457_);
  or (_38467_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_38468_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_38469_, _38468_, _38467_);
  or (_38470_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_38471_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_38472_, _38471_, _38470_);
  or (_38473_, _38472_, _38469_);
  and (_38474_, _06880_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_38475_, \oc8051_golden_model_1.B [7], _28098_);
  or (_38476_, _38475_, _38474_);
  nand (_38478_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_38479_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_38480_, _38479_, _38478_);
  or (_38481_, _38480_, _38476_);
  or (_38482_, _38481_, _38473_);
  or (_38483_, _38482_, _38465_);
  and (property_invalid_b_reg, _38483_, _37562_);
  nand (_38484_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_38485_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_38486_, _38485_, _38484_);
  and (_38488_, _07634_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_38489_, \oc8051_golden_model_1.ACC [2], _39256_);
  or (_38490_, _38489_, _38488_);
  or (_38491_, _38490_, _38486_);
  nor (_38492_, _03320_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_38493_, _03320_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_38494_, _38493_, _38492_);
  and (_38495_, _03397_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38496_, _03397_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_38497_, _38496_, _38495_);
  or (_38499_, _38497_, _38494_);
  or (_38500_, _38499_, _38491_);
  or (_38501_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38502_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_38503_, _38502_, _38501_);
  or (_38504_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_38505_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_38506_, _38505_, _38504_);
  or (_38507_, _38506_, _38503_);
  and (_38508_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_38510_, \oc8051_golden_model_1.ACC [6], _01245_);
  or (_38511_, _38510_, _38508_);
  nand (_38512_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_38513_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_38514_, _38513_, _38512_);
  or (_38515_, _38514_, _38511_);
  or (_38516_, _38515_, _38507_);
  or (_38517_, _38516_, _38500_);
  and (property_invalid_acc, _38517_, _37562_);
  nor (_38518_, _32926_, _44168_);
  and (_38520_, _32926_, _44168_);
  and (_38521_, _34693_, _43417_);
  nor (_38522_, _34693_, _43417_);
  and (_38523_, _33990_, _43483_);
  or (_38524_, _38523_, _38522_);
  or (_38525_, _38524_, _38521_);
  and (_38526_, _35049_, _43411_);
  and (_38527_, _34349_, _43445_);
  nor (_38528_, _35699_, _38727_);
  and (_38529_, _35699_, _38727_);
  and (_38531_, _36912_, _38713_);
  and (_38532_, _11993_, _38749_);
  nor (_38533_, _36307_, _38717_);
  or (_38534_, _38533_, _38532_);
  and (_38535_, _36608_, _38738_);
  and (_38536_, _36307_, _38717_);
  or (_38537_, _38536_, _38535_);
  or (_38538_, _38537_, _38534_);
  nor (_38539_, _36001_, _38732_);
  and (_38540_, _36001_, _38732_);
  nor (_38542_, _32541_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_38543_, _32541_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_38544_, _38543_, _38542_);
  or (_38545_, _38544_, _38540_);
  or (_38546_, _38545_, _38539_);
  nor (_38547_, _36608_, _38738_);
  nor (_38548_, _11993_, _38749_);
  or (_38549_, _38548_, _38547_);
  or (_38550_, _38549_, _38546_);
  or (_38551_, _38550_, _38538_);
  or (_38553_, _38551_, _38531_);
  nand (_38554_, _35369_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_38555_, _35369_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38556_, _38555_, _38554_);
  nand (_38557_, _37223_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_38558_, _37223_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38559_, _38558_, _38557_);
  nor (_38560_, _36912_, _38713_);
  or (_38561_, _38560_, _38559_);
  or (_38562_, _38561_, _38556_);
  or (_38564_, _38562_, _38553_);
  or (_38565_, _38564_, _38529_);
  or (_38566_, _38565_, _38528_);
  or (_38567_, _38566_, _38527_);
  nor (_38568_, _34349_, _43445_);
  nor (_38569_, _33638_, _43511_);
  and (_38570_, _33638_, _43511_);
  or (_38571_, _38570_, _38569_);
  or (_38572_, _38571_, _38568_);
  or (_38573_, _38572_, _38567_);
  or (_38575_, _38573_, _38526_);
  nor (_38576_, _33990_, _43483_);
  nor (_38577_, _35049_, _43411_);
  or (_38578_, _38577_, _38576_);
  or (_38579_, _38578_, _38575_);
  and (_38580_, _33288_, _43547_);
  nor (_38581_, _33288_, _43547_);
  or (_38582_, _38581_, _38580_);
  or (_38583_, _38582_, _38579_);
  or (_38584_, _38583_, _38525_);
  or (_38586_, _38584_, _38520_);
  or (_38587_, _38586_, _38518_);
  and (property_invalid_pc, _38587_, _37529_);
  buf (_01418_, _41991_);
  buf (_01470_, _41991_);
  buf (_01521_, _41991_);
  buf (_01573_, _41991_);
  buf (_01625_, _41991_);
  buf (_01670_, _41991_);
  buf (_01716_, _41991_);
  buf (_01769_, _41991_);
  buf (_01820_, _41991_);
  buf (_01872_, _41991_);
  buf (_01924_, _41991_);
  buf (_01976_, _41991_);
  buf (_02028_, _41991_);
  buf (_02080_, _41991_);
  buf (_02132_, _41991_);
  buf (_02184_, _41991_);
  buf (_39095_, _38992_);
  buf (_39096_, _38993_);
  buf (_39109_, _38992_);
  buf (_39110_, _38993_);
  buf (_39422_, _39011_);
  buf (_39423_, _39013_);
  buf (_39424_, _39014_);
  buf (_39425_, _39015_);
  buf (_39426_, _39016_);
  buf (_39427_, _39017_);
  buf (_39428_, _39019_);
  buf (_39430_, _39020_);
  buf (_39431_, _39021_);
  buf (_39432_, _39022_);
  buf (_39433_, _39023_);
  buf (_39434_, _39025_);
  buf (_39435_, _39026_);
  buf (_39436_, _39027_);
  buf (_39488_, _39011_);
  buf (_39489_, _39013_);
  buf (_39490_, _39014_);
  buf (_39491_, _39015_);
  buf (_39492_, _39016_);
  buf (_39493_, _39017_);
  buf (_39494_, _39019_);
  buf (_39496_, _39020_);
  buf (_39497_, _39021_);
  buf (_39498_, _39022_);
  buf (_39499_, _39023_);
  buf (_39500_, _39025_);
  buf (_39501_, _39026_);
  buf (_39502_, _39027_);
  buf (_39829_, _39795_);
  buf (_39944_, _39795_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (property_invalid_psw_1_r, _00006_);
  dff (property_invalid_sp_1_r, _00007_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _01422_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _01426_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _01430_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _01434_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _01438_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _01442_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _01446_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _01415_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _01418_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _01474_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _01478_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _01482_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _01485_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _01489_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _01493_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _01497_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _01467_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _01470_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _01928_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _01932_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _01936_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _01940_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _01944_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _01948_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _01951_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _01921_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _01924_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _01980_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _01984_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _01988_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _01992_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _01996_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _02000_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _02004_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _01973_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _01976_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _02032_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _02036_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _02040_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _02044_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _02048_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _02052_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _02056_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _02025_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _02028_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _02084_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _02088_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _02092_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _02096_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _02100_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _02104_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _02108_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _02077_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _02080_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _02136_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _02140_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _02144_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _02148_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _02152_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _02156_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _02160_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _02129_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _02132_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _02188_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _02192_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _02196_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _02200_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _02204_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _02208_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _02212_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _02181_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _02184_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _01525_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _01529_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _01533_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _01537_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _01541_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _01545_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _01549_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _01518_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _01521_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _01577_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _01581_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _01585_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _01589_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _01593_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _01596_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _01600_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _01570_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _01573_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _01629_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _01632_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _01636_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _01640_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _01644_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _01648_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _01652_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _01622_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _01625_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _01671_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _01672_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _01675_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _01679_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _01683_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _01687_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _01691_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _01669_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _01670_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _01720_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _01724_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _01728_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _01732_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _01736_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _01740_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _01744_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _01713_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _01716_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _01773_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _01777_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _01781_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _01785_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _01788_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _01792_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _01796_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _01766_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _01769_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _01824_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _01828_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _01832_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _01836_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _01840_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _01844_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _01848_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _01818_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _01820_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _01876_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _01880_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _01884_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _01888_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _01892_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _01895_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _01899_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _01869_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _01872_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40976_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40977_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40978_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40979_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40981_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40982_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40983_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40744_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40964_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40965_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40966_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40967_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40969_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40970_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40971_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40972_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40952_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40953_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40954_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40955_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40957_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40958_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40959_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40960_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40940_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40941_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40942_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40943_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40944_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40946_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40947_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40948_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40927_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40929_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40930_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40931_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40932_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40933_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40935_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40936_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40915_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40916_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40918_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40919_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40920_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40921_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40922_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40924_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40903_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40904_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40906_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40907_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40908_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40909_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40910_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40912_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40891_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40892_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40893_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40895_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40896_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40897_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40898_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40899_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40878_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40880_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40881_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40882_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40883_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40884_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40886_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40887_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40866_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40867_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40869_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40870_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40871_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40872_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40873_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40875_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40854_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40855_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40857_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40858_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40859_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40860_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40861_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40863_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40842_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40843_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40844_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40846_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40847_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40848_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40849_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40850_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40829_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40831_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40832_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40833_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40834_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40835_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40837_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40838_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40817_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40818_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40819_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40821_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40822_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40823_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40824_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40825_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40804_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40806_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40807_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40808_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40809_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40810_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40812_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40813_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40790_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40792_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40793_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40795_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40796_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40797_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40799_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40800_);
  dff (\oc8051_golden_model_1.B [0], _43424_);
  dff (\oc8051_golden_model_1.B [1], _43425_);
  dff (\oc8051_golden_model_1.B [2], _43426_);
  dff (\oc8051_golden_model_1.B [3], _43428_);
  dff (\oc8051_golden_model_1.B [4], _43429_);
  dff (\oc8051_golden_model_1.B [5], _43430_);
  dff (\oc8051_golden_model_1.B [6], _43431_);
  dff (\oc8051_golden_model_1.B [7], _40745_);
  dff (\oc8051_golden_model_1.ACC [0], _43433_);
  dff (\oc8051_golden_model_1.ACC [1], _43434_);
  dff (\oc8051_golden_model_1.ACC [2], _43435_);
  dff (\oc8051_golden_model_1.ACC [3], _43436_);
  dff (\oc8051_golden_model_1.ACC [4], _43437_);
  dff (\oc8051_golden_model_1.ACC [5], _43438_);
  dff (\oc8051_golden_model_1.ACC [6], _43439_);
  dff (\oc8051_golden_model_1.ACC [7], _40746_);
  dff (\oc8051_golden_model_1.DPL [0], _43440_);
  dff (\oc8051_golden_model_1.DPL [1], _43441_);
  dff (\oc8051_golden_model_1.DPL [2], _43442_);
  dff (\oc8051_golden_model_1.DPL [3], _43443_);
  dff (\oc8051_golden_model_1.DPL [4], _43444_);
  dff (\oc8051_golden_model_1.DPL [5], _43447_);
  dff (\oc8051_golden_model_1.DPL [6], _43448_);
  dff (\oc8051_golden_model_1.DPL [7], _40747_);
  dff (\oc8051_golden_model_1.DPH [0], _43449_);
  dff (\oc8051_golden_model_1.DPH [1], _43452_);
  dff (\oc8051_golden_model_1.DPH [2], _43453_);
  dff (\oc8051_golden_model_1.DPH [3], _43454_);
  dff (\oc8051_golden_model_1.DPH [4], _43455_);
  dff (\oc8051_golden_model_1.DPH [5], _43456_);
  dff (\oc8051_golden_model_1.DPH [6], _43457_);
  dff (\oc8051_golden_model_1.DPH [7], _40748_);
  dff (\oc8051_golden_model_1.IE [0], _43458_);
  dff (\oc8051_golden_model_1.IE [1], _43459_);
  dff (\oc8051_golden_model_1.IE [2], _43460_);
  dff (\oc8051_golden_model_1.IE [3], _43461_);
  dff (\oc8051_golden_model_1.IE [4], _43462_);
  dff (\oc8051_golden_model_1.IE [5], _43463_);
  dff (\oc8051_golden_model_1.IE [6], _43464_);
  dff (\oc8051_golden_model_1.IE [7], _40750_);
  dff (\oc8051_golden_model_1.IP [0], _43467_);
  dff (\oc8051_golden_model_1.IP [1], _43468_);
  dff (\oc8051_golden_model_1.IP [2], _43469_);
  dff (\oc8051_golden_model_1.IP [3], _43472_);
  dff (\oc8051_golden_model_1.IP [4], _43473_);
  dff (\oc8051_golden_model_1.IP [5], _43474_);
  dff (\oc8051_golden_model_1.IP [6], _43475_);
  dff (\oc8051_golden_model_1.IP [7], _40751_);
  dff (\oc8051_golden_model_1.P0 [0], _43476_);
  dff (\oc8051_golden_model_1.P0 [1], _43477_);
  dff (\oc8051_golden_model_1.P0 [2], _43478_);
  dff (\oc8051_golden_model_1.P0 [3], _43479_);
  dff (\oc8051_golden_model_1.P0 [4], _43480_);
  dff (\oc8051_golden_model_1.P0 [5], _43481_);
  dff (\oc8051_golden_model_1.P0 [6], _43482_);
  dff (\oc8051_golden_model_1.P0 [7], _40752_);
  dff (\oc8051_golden_model_1.P1 [0], _43485_);
  dff (\oc8051_golden_model_1.P1 [1], _43486_);
  dff (\oc8051_golden_model_1.P1 [2], _43487_);
  dff (\oc8051_golden_model_1.P1 [3], _43488_);
  dff (\oc8051_golden_model_1.P1 [4], _43489_);
  dff (\oc8051_golden_model_1.P1 [5], _43492_);
  dff (\oc8051_golden_model_1.P1 [6], _43493_);
  dff (\oc8051_golden_model_1.P1 [7], _40753_);
  dff (\oc8051_golden_model_1.P2 [0], _43494_);
  dff (\oc8051_golden_model_1.P2 [1], _43495_);
  dff (\oc8051_golden_model_1.P2 [2], _43496_);
  dff (\oc8051_golden_model_1.P2 [3], _43497_);
  dff (\oc8051_golden_model_1.P2 [4], _43498_);
  dff (\oc8051_golden_model_1.P2 [5], _43499_);
  dff (\oc8051_golden_model_1.P2 [6], _43500_);
  dff (\oc8051_golden_model_1.P2 [7], _40754_);
  dff (\oc8051_golden_model_1.P3 [0], _43503_);
  dff (\oc8051_golden_model_1.P3 [1], _43504_);
  dff (\oc8051_golden_model_1.P3 [2], _43505_);
  dff (\oc8051_golden_model_1.P3 [3], _43506_);
  dff (\oc8051_golden_model_1.P3 [4], _43507_);
  dff (\oc8051_golden_model_1.P3 [5], _43508_);
  dff (\oc8051_golden_model_1.P3 [6], _43509_);
  dff (\oc8051_golden_model_1.P3 [7], _40756_);
  dff (\oc8051_golden_model_1.PSW [0], _43512_);
  dff (\oc8051_golden_model_1.PSW [1], _43513_);
  dff (\oc8051_golden_model_1.PSW [2], _43514_);
  dff (\oc8051_golden_model_1.PSW [3], _43515_);
  dff (\oc8051_golden_model_1.PSW [4], _43516_);
  dff (\oc8051_golden_model_1.PSW [5], _43517_);
  dff (\oc8051_golden_model_1.PSW [6], _43518_);
  dff (\oc8051_golden_model_1.PSW [7], _40757_);
  dff (\oc8051_golden_model_1.PCON [0], _43521_);
  dff (\oc8051_golden_model_1.PCON [1], _43522_);
  dff (\oc8051_golden_model_1.PCON [2], _43523_);
  dff (\oc8051_golden_model_1.PCON [3], _43524_);
  dff (\oc8051_golden_model_1.PCON [4], _43525_);
  dff (\oc8051_golden_model_1.PCON [5], _43526_);
  dff (\oc8051_golden_model_1.PCON [6], _43527_);
  dff (\oc8051_golden_model_1.PCON [7], _40758_);
  dff (\oc8051_golden_model_1.SBUF [0], _43530_);
  dff (\oc8051_golden_model_1.SBUF [1], _43531_);
  dff (\oc8051_golden_model_1.SBUF [2], _43532_);
  dff (\oc8051_golden_model_1.SBUF [3], _43533_);
  dff (\oc8051_golden_model_1.SBUF [4], _43534_);
  dff (\oc8051_golden_model_1.SBUF [5], _43535_);
  dff (\oc8051_golden_model_1.SBUF [6], _43536_);
  dff (\oc8051_golden_model_1.SBUF [7], _40759_);
  dff (\oc8051_golden_model_1.SCON [0], _43537_);
  dff (\oc8051_golden_model_1.SCON [1], _43540_);
  dff (\oc8051_golden_model_1.SCON [2], _43541_);
  dff (\oc8051_golden_model_1.SCON [3], _43542_);
  dff (\oc8051_golden_model_1.SCON [4], _43543_);
  dff (\oc8051_golden_model_1.SCON [5], _43544_);
  dff (\oc8051_golden_model_1.SCON [6], _43545_);
  dff (\oc8051_golden_model_1.SCON [7], _40760_);
  dff (\oc8051_golden_model_1.SP [0], _43548_);
  dff (\oc8051_golden_model_1.SP [1], _43549_);
  dff (\oc8051_golden_model_1.SP [2], _43550_);
  dff (\oc8051_golden_model_1.SP [3], _43551_);
  dff (\oc8051_golden_model_1.SP [4], _43552_);
  dff (\oc8051_golden_model_1.SP [5], _43553_);
  dff (\oc8051_golden_model_1.SP [6], _43554_);
  dff (\oc8051_golden_model_1.SP [7], _40762_);
  dff (\oc8051_golden_model_1.TCON [0], _43555_);
  dff (\oc8051_golden_model_1.TCON [1], _43556_);
  dff (\oc8051_golden_model_1.TCON [2], _43557_);
  dff (\oc8051_golden_model_1.TCON [3], _43560_);
  dff (\oc8051_golden_model_1.TCON [4], _43561_);
  dff (\oc8051_golden_model_1.TCON [5], _43562_);
  dff (\oc8051_golden_model_1.TCON [6], _43563_);
  dff (\oc8051_golden_model_1.TCON [7], _40763_);
  dff (\oc8051_golden_model_1.TH0 [0], _43566_);
  dff (\oc8051_golden_model_1.TH0 [1], _43567_);
  dff (\oc8051_golden_model_1.TH0 [2], _43568_);
  dff (\oc8051_golden_model_1.TH0 [3], _43569_);
  dff (\oc8051_golden_model_1.TH0 [4], _43570_);
  dff (\oc8051_golden_model_1.TH0 [5], _43571_);
  dff (\oc8051_golden_model_1.TH0 [6], _43572_);
  dff (\oc8051_golden_model_1.TH0 [7], _40764_);
  dff (\oc8051_golden_model_1.TH1 [0], _43574_);
  dff (\oc8051_golden_model_1.TH1 [1], _43575_);
  dff (\oc8051_golden_model_1.TH1 [2], _43576_);
  dff (\oc8051_golden_model_1.TH1 [3], _43577_);
  dff (\oc8051_golden_model_1.TH1 [4], _43578_);
  dff (\oc8051_golden_model_1.TH1 [5], _43581_);
  dff (\oc8051_golden_model_1.TH1 [6], _43582_);
  dff (\oc8051_golden_model_1.TH1 [7], _40765_);
  dff (\oc8051_golden_model_1.TL0 [0], _43583_);
  dff (\oc8051_golden_model_1.TL0 [1], _43585_);
  dff (\oc8051_golden_model_1.TL0 [2], _43586_);
  dff (\oc8051_golden_model_1.TL0 [3], _43587_);
  dff (\oc8051_golden_model_1.TL0 [4], _43588_);
  dff (\oc8051_golden_model_1.TL0 [5], _43589_);
  dff (\oc8051_golden_model_1.TL0 [6], _43590_);
  dff (\oc8051_golden_model_1.TL0 [7], _40766_);
  dff (\oc8051_golden_model_1.TL1 [0], _43592_);
  dff (\oc8051_golden_model_1.TL1 [1], _43593_);
  dff (\oc8051_golden_model_1.TL1 [2], _43594_);
  dff (\oc8051_golden_model_1.TL1 [3], _43595_);
  dff (\oc8051_golden_model_1.TL1 [4], _43596_);
  dff (\oc8051_golden_model_1.TL1 [5], _43597_);
  dff (\oc8051_golden_model_1.TL1 [6], _43598_);
  dff (\oc8051_golden_model_1.TL1 [7], _40768_);
  dff (\oc8051_golden_model_1.TMOD [0], _43600_);
  dff (\oc8051_golden_model_1.TMOD [1], _43601_);
  dff (\oc8051_golden_model_1.TMOD [2], _43602_);
  dff (\oc8051_golden_model_1.TMOD [3], _43604_);
  dff (\oc8051_golden_model_1.TMOD [4], _43605_);
  dff (\oc8051_golden_model_1.TMOD [5], _43606_);
  dff (\oc8051_golden_model_1.TMOD [6], _43607_);
  dff (\oc8051_golden_model_1.TMOD [7], _40769_);
  dff (\oc8051_golden_model_1.PC [0], _43608_);
  dff (\oc8051_golden_model_1.PC [1], _43611_);
  dff (\oc8051_golden_model_1.PC [2], _43612_);
  dff (\oc8051_golden_model_1.PC [3], _43613_);
  dff (\oc8051_golden_model_1.PC [4], _43614_);
  dff (\oc8051_golden_model_1.PC [5], _43615_);
  dff (\oc8051_golden_model_1.PC [6], _43616_);
  dff (\oc8051_golden_model_1.PC [7], _43617_);
  dff (\oc8051_golden_model_1.PC [8], _43618_);
  dff (\oc8051_golden_model_1.PC [9], _43619_);
  dff (\oc8051_golden_model_1.PC [10], _43620_);
  dff (\oc8051_golden_model_1.PC [11], _43623_);
  dff (\oc8051_golden_model_1.PC [12], _43624_);
  dff (\oc8051_golden_model_1.PC [13], _43625_);
  dff (\oc8051_golden_model_1.PC [14], _43626_);
  dff (\oc8051_golden_model_1.PC [15], _40770_);
  dff (\oc8051_golden_model_1.P0INREG [0], _43627_);
  dff (\oc8051_golden_model_1.P0INREG [1], _43628_);
  dff (\oc8051_golden_model_1.P0INREG [2], _43629_);
  dff (\oc8051_golden_model_1.P0INREG [3], _43630_);
  dff (\oc8051_golden_model_1.P0INREG [4], _43631_);
  dff (\oc8051_golden_model_1.P0INREG [5], _43632_);
  dff (\oc8051_golden_model_1.P0INREG [6], _43633_);
  dff (\oc8051_golden_model_1.P0INREG [7], _40771_);
  dff (\oc8051_golden_model_1.P1INREG [0], _43636_);
  dff (\oc8051_golden_model_1.P1INREG [1], _43637_);
  dff (\oc8051_golden_model_1.P1INREG [2], _43638_);
  dff (\oc8051_golden_model_1.P1INREG [3], _43639_);
  dff (\oc8051_golden_model_1.P1INREG [4], _43640_);
  dff (\oc8051_golden_model_1.P1INREG [5], _43643_);
  dff (\oc8051_golden_model_1.P1INREG [6], _43644_);
  dff (\oc8051_golden_model_1.P1INREG [7], _40772_);
  dff (\oc8051_golden_model_1.P2INREG [0], _43645_);
  dff (\oc8051_golden_model_1.P2INREG [1], _43646_);
  dff (\oc8051_golden_model_1.P2INREG [2], _43647_);
  dff (\oc8051_golden_model_1.P2INREG [3], _43648_);
  dff (\oc8051_golden_model_1.P2INREG [4], _43649_);
  dff (\oc8051_golden_model_1.P2INREG [5], _43650_);
  dff (\oc8051_golden_model_1.P2INREG [6], _43651_);
  dff (\oc8051_golden_model_1.P2INREG [7], _40774_);
  dff (\oc8051_golden_model_1.P3INREG [0], _43654_);
  dff (\oc8051_golden_model_1.P3INREG [1], _43655_);
  dff (\oc8051_golden_model_1.P3INREG [2], _43656_);
  dff (\oc8051_golden_model_1.P3INREG [3], _43657_);
  dff (\oc8051_golden_model_1.P3INREG [4], _43658_);
  dff (\oc8051_golden_model_1.P3INREG [5], _43659_);
  dff (\oc8051_golden_model_1.P3INREG [6], _43660_);
  dff (\oc8051_golden_model_1.P3INREG [7], _40775_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03002_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03013_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03034_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03056_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03077_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00881_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03088_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00850_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03099_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03110_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03121_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03132_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03143_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03154_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03165_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00902_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02454_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22423_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02649_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02844_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03045_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03256_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03457_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03658_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03859_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04060_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04161_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04262_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04363_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04464_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04565_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04666_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04767_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24609_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _39004_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _39005_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _39006_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _39007_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _39008_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _39009_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _39010_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38991_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _39011_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _39013_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _39014_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _39015_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _39016_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _39017_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _39019_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38992_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _39020_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _39021_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _39022_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _39023_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _39025_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _39026_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _39027_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38993_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _30457_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05999_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _30460_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _06002_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _30462_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _30464_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _06005_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _30466_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _30468_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06008_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _30470_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _06011_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _30472_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _30474_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _30476_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _06014_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _30478_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _06017_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _06020_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _06079_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _06081_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _05984_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _06084_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _06087_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05987_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _06090_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _05990_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _06093_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _06096_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _06099_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _06102_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _06105_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _06108_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _06111_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _05993_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _05996_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39168_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39171_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39173_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39176_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39052_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39187_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39192_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39054_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39376_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39377_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39378_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39379_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39381_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39383_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39384_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39385_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39386_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39387_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39388_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39389_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39390_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39391_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39392_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39394_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39395_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39396_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39397_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39398_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39399_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39401_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39402_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39403_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39405_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39406_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39407_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39408_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39117_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39091_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39410_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39411_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39412_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39413_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39092_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39414_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39415_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39416_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39417_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39418_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39420_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39421_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39093_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39422_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39423_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39425_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39426_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39095_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39430_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39432_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39433_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39096_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39097_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39098_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39437_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39438_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39439_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39441_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39442_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39099_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39446_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39448_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39450_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39452_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39453_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39454_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39455_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39456_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39457_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39458_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39459_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39460_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39101_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39461_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39463_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39464_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39465_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39466_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39468_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39469_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39470_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39471_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39472_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39474_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39475_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39476_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39477_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39102_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39103_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39106_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39104_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39478_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39479_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39480_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39481_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39482_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39483_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39485_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39107_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39486_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39487_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39108_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39488_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39489_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39490_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39491_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39492_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39493_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39494_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39109_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39496_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39497_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39498_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39499_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39500_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39501_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39110_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _39111_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39503_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39504_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39505_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39507_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39508_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39509_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39510_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39113_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _39114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39115_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39511_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39512_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39513_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39116_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39514_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39515_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39516_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39518_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39519_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39520_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39521_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39524_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39525_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39526_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39527_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39529_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39530_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39531_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39532_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39533_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39534_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39535_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39536_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39537_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39538_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39540_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39541_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39542_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39543_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39544_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39545_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39546_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39547_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39118_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39548_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39549_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39550_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39551_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39552_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39553_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39554_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39120_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39122_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39555_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39556_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39557_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39558_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39559_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39561_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39562_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39563_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39564_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39565_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39567_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39568_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39570_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39125_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39126_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39572_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39573_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39574_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39575_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39576_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39577_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39578_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39580_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39581_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39583_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39584_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39585_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39586_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39127_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39128_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39942_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39960_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39961_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39962_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39963_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39964_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39965_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39966_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39943_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39944_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39967_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39968_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _44007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _44011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _44015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _44019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _44023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _44027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _44031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _43059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _43975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _43979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _43983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _43987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _43991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _43995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _43999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _44002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _43315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _43321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _43327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _43333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _43339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _43345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _43348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _43351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _43359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _43363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _43367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _43371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _43375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _43379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _43383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _43386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _43394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _43398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _43402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _43406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _43410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _43414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _43418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _43421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _43610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _43635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _43653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _43664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _43668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _43672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _43676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _43679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _43446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _43466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _43484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _43502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _43520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _43539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _43559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _43573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _43814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _43818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _43822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _43826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _43830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _43834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _43838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _43841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _43782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _43786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _43790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _43794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _43798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _43802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _43806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _43809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _43748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _43752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _43756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _43760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _43764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _43767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _43771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _43774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _43716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _43720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _43724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _43728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _43732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _43736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _43740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _43743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _43684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _43688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _43692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _43696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _43700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _43704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _43708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _43711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _43846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _43850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _43854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _43858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _43862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _43866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _43870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _43873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _43943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _43947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _43951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _43955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _43959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _43963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _43967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _43970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _43911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _43915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _43919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _43923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _43927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _43931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _43935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _43938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _43878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _43882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _43886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _43890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _43894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _43898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _43902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _43905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _01396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _01397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _01399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _01401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _01403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _01405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _01407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _43047_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39826_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39827_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39891_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39892_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39893_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39894_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39895_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39896_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39897_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39828_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24198_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24210_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24222_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08932_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08943_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08975_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08986_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13674_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13713_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _41991_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _42909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _42911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42913_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _42915_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _42917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41989_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _42923_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _41987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _41985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _42925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _42927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _41983_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _42929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _42931_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _41981_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _42933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _42935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _41946_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _41944_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _41942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _41940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _42937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _42939_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _42941_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _41938_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _42943_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _42945_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _42947_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _42949_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _42951_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _42953_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _42954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41936_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _42956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _42958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _42960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _42962_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _42964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _42966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _42968_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _41933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41393_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41394_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41396_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41398_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41400_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41401_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41403_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35472_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41405_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41407_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41408_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41410_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41414_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35495_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41417_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41422_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41426_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41428_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35518_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41429_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41431_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41436_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41438_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41440_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35541_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21467_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21491_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21515_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21527_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16533_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09532_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10678_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10689_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10733_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10744_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09553_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0988 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0988 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0988 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0988 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0988 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0988 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0988 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0989 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0990 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0991 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0992 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0993 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0995 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0996 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1011 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1011 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1011 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1011 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1011 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1011 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1011 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1018 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1019 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.n1027 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1027 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1027 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1027 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1027 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1043 , \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.n1044 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1044 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1044 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1044 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1044 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1044 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1044 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1137 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1137 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1137 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1137 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1139 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1141 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1141 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1142 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1142 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1143 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1144 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1144 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1145 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1145 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1146 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1194 , \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n1239 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1240 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1240 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1240 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1240 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1240 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1240 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1240 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1241 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1241 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1241 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1241 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1241 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1241 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1241 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1242 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1242 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1242 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1242 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1242 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1242 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1242 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1242 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1243 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1244 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1244 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1244 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1247 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1247 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1247 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1247 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1247 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1248 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1248 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1248 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1248 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1248 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1248 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1248 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1249 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1251 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1252 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1253 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1254 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1255 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1264 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1280 , \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.n1281 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1281 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1281 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1281 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1281 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1281 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1281 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1323 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1323 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1323 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1323 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1323 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1323 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1323 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1323 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1323 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1323 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1323 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1323 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1323 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1323 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1323 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1323 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1325 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1325 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1325 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1325 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1325 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1325 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1325 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1327 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1328 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1329 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1330 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1331 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1332 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1340 , \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.n1341 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1341 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1341 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1341 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1341 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1341 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1343 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1347 [8], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1349 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1349 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1349 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1349 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1350 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1354 [4], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1356 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1356 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1356 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1356 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1356 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1356 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1356 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1356 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1356 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1364 , \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1365 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1365 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1365 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1365 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1365 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1365 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1366 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1366 [6], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1381 , \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.n1382 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1382 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1382 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1382 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1404 [8], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1405 , \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1410 [4], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1411 , \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1419 , \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1420 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1420 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1420 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1420 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1420 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1420 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1421 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1421 [1], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1421 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1421 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1421 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1421 [5], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1421 [6], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1436 , \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.n1437 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1437 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1437 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1437 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1439 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1439 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1439 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1439 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1439 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1439 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1439 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1439 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1439 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1441 [8], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1442 , \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1443 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1443 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1443 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1443 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1444 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1444 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1444 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1446 [4], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1447 , \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1448 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1448 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1448 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1448 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1448 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1448 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1448 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1448 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1448 [8], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1455 , \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1456 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1456 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1456 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1456 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1456 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1456 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1457 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1457 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1457 [6], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1472 , \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1473 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1473 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1473 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1473 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1476 [8], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1477 , \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1484 , \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1485 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1485 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1485 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1485 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1485 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1485 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1486 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1486 [1], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1486 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1486 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1486 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1486 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1486 [6], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1489 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1489 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1489 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1489 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1489 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1489 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1489 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1489 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1489 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1491 [8], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1493 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1495 [4], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1496 , \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1497 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1497 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1497 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1497 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1497 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1497 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1497 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1497 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1497 [8], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1521 , \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1522 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1524 [4], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1525 , \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1527 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1527 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1527 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1527 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1527 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1527 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1527 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1528 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1528 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1530 [8], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1531 , \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1538 , \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1539 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1539 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1539 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1539 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1539 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1539 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1540 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1540 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1540 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1540 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1540 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1540 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1540 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1541 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1541 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1541 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1541 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1541 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1541 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1541 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1543 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1543 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1543 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1543 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1543 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1543 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1543 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1544 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1544 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1544 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1547 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1547 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1548 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1548 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1548 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1549 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1549 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1549 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1549 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1549 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1549 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1549 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1549 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1550 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1550 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1550 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1550 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1550 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1550 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1550 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1550 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1551 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1552 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1553 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1555 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1557 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1559 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1566 , \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1571 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [8], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1575 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1575 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [4], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1585 , \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1586 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1586 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1586 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1586 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1586 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1586 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1587 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1602 , \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.n1603 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1603 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1603 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1603 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [8], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1608 , \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1610 [4], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1611 , \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1618 , \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1619 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1619 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1619 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1619 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1619 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1619 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1620 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1620 [1], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1620 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1620 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1620 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1620 [5], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1620 [6], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1635 , \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.n1636 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1636 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1636 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1636 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [8], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1641 , \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1643 [4], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1644 , \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1651 , \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1652 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1652 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1652 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1652 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1652 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1652 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1653 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1653 [1], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1653 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1653 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1653 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1653 [5], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1653 [6], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1668 , \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.n1669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [8], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1674 , \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1676 [4], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1677 , \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1684 , \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1685 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1685 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1685 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1685 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1685 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1685 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1686 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1686 [1], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1686 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1686 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1686 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1686 [5], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1686 [6], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1701 , \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.n1702 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1702 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1702 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1702 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1727 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1727 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1727 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1727 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1727 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1727 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1727 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1728 [0], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1728 [1], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1728 [2], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1728 [3], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1728 [4], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1728 [5], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1728 [6], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1729 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1784 , \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.n1785 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1785 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1785 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1785 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1785 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1785 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1785 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1801 , \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.n1802 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1802 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1802 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1802 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1802 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1802 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1802 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1818 , \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.n1819 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1819 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1819 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1819 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1819 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1819 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1819 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1835 , \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.n1836 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1836 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1836 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1836 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1836 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1836 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1836 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1859 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1859 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1859 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1859 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1859 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1859 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1859 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1860 [0], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1860 [1], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1860 [2], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1860 [3], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1860 [4], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1860 [5], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1860 [6], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1861 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1916 , \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.n1917 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1917 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1917 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1917 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1917 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1917 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1917 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1933 , \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.n1934 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1934 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1934 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1934 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1934 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1934 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1934 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1950 , \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.n1951 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1951 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1951 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1951 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1951 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1951 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1951 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1967 , \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.n1968 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1968 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1968 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1968 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1968 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1968 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1968 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2065 , \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.n2066 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2066 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2066 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2066 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2066 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2066 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2066 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2082 , \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.n2083 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2083 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2083 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2083 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2083 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2083 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2083 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2099 , \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.n2100 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2100 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2100 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2100 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2100 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2100 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2116 , \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.n2117 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2117 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2117 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2117 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2117 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2117 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2117 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2121 , \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2122 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2122 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2122 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2122 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2122 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2122 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2122 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2123 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2123 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2123 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2123 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2123 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2123 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2124 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2124 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2124 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2124 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2124 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2124 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2124 [6], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2125 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2125 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2125 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2125 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2125 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2125 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2125 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2140 , \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.n2141 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2141 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2141 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2141 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2141 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2141 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2180 , \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2181 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2181 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2181 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2181 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2181 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2181 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2181 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2181 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2182 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2182 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2182 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2182 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2182 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2182 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2182 [6], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2183 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2183 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2183 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2183 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2183 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2183 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2183 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2190 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2190 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2190 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2190 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2191 , \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2192 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2192 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2192 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2192 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2192 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2192 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2193 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2193 [1], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2193 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2193 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2193 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2193 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2193 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2208 , \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.n2209 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2209 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2209 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2209 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2209 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2209 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2421 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2424 , \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2426 , \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2432 , \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2433 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2433 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2433 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2433 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2433 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2433 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2434 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2434 [1], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2434 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2434 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2434 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2434 [5], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2434 [6], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2449 , \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.n2450 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2450 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2450 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2450 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 , \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2456 , \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2462 , \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2463 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2463 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2463 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2463 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2463 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2463 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2464 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2464 [1], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2464 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2464 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2464 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2464 [5], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2464 [6], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2479 , \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.n2480 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2480 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2480 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2480 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 , \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2486 , \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2492 , \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2493 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2493 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2493 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2494 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2494 [1], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2494 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2494 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2494 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2494 [5], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2494 [6], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2509 , \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.n2510 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2510 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2510 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2510 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 , \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2516 , \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2522 , \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2523 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2523 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2523 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2523 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2523 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2523 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2524 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2524 [1], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2524 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2524 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2524 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2524 [5], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2524 [6], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2539 , \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.n2540 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2540 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2540 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2540 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2545 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2545 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2545 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2545 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2545 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2545 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2545 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2547 [6], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2548 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2548 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2548 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2552 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2552 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2552 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2552 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2552 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2552 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2552 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2552 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2552 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2558 , \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2559 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2559 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2559 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2560 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2575 , \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.n2576 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2576 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2576 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2576 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2576 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2576 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2579 , \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2581 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2581 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2581 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2581 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2581 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2581 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2581 [6], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2582 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2582 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2582 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2582 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2582 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2582 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2582 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2614 , \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2615 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2615 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2615 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2615 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2615 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2615 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2615 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2615 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2616 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2616 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2616 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2616 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2616 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2616 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2616 [6], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2617 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2617 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2617 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2617 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2617 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2617 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2617 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2622 , \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2623 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2623 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2623 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2623 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2624 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2624 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2624 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2624 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2624 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2624 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2624 [6], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2625 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2625 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2625 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2625 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2625 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2625 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2625 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2630 , \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2631 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2631 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2631 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2631 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2631 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2631 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2631 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2631 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2632 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2632 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2632 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2632 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2632 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2632 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2632 [6], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2633 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2633 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2633 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2633 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2633 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2633 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2633 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2638 , \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2639 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2639 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2639 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2640 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2640 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2640 [6], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2641 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2641 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2641 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2641 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2641 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2641 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2641 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2646 , \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2647 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2647 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2647 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2647 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2647 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2647 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2647 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2647 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2648 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2648 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2648 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2648 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2648 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2648 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2648 [6], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2649 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2649 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2649 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2649 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2649 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2649 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2649 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2674 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2674 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2674 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2674 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2674 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2674 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2675 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2675 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2675 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2675 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2675 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2675 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2675 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2676 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2676 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2676 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2676 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2676 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2676 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2676 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2676 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2677 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2677 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2677 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2677 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2678 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2678 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2678 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2678 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2678 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2678 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2679 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2680 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2681 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2682 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2683 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2684 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2685 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2686 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2693 , \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2715 [0], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2715 [1], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2715 [2], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2715 [3], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2715 [4], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2715 [5], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2715 [6], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2731 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2731 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2731 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2731 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2731 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2731 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2731 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2732 , \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2733 , \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2734 , \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2735 , \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2736 , \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2737 , \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2738 , \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2739 , \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2746 , \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.n2747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2747 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2747 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2747 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2762 , \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.n2763 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2763 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2763 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2763 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2763 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2763 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2763 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2795 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2795 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2795 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2795 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2795 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2795 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2795 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2795 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2796 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2796 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2796 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2796 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2796 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2796 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2796 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2797 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2797 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2797 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2797 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2797 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2797 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2797 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2797 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 , \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2818 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2818 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2818 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2818 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2818 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2818 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2818 [6], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2833 , \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.n2834 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2834 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2834 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2834 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2834 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2834 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2838 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2839 [0], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2839 [1], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2839 [2], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2839 [3], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2840 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2840 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2840 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2840 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2841 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2842 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2843 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2844 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2855 , \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.n2856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2874 , \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.n2875 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2875 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2875 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2875 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2875 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2875 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2875 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2891 , \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.n2892 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2892 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2892 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2892 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2892 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2892 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2892 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(ie_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(ie_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(ie_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(ie_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(ie_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(ie_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(ie_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(ie_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
