
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_acc);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1071 ;
  wire [3:0] \oc8051_golden_model_1.n1073 ;
  wire [3:0] \oc8051_golden_model_1.n1075 ;
  wire [3:0] \oc8051_golden_model_1.n1076 ;
  wire [3:0] \oc8051_golden_model_1.n1077 ;
  wire [3:0] \oc8051_golden_model_1.n1078 ;
  wire [3:0] \oc8051_golden_model_1.n1079 ;
  wire [3:0] \oc8051_golden_model_1.n1080 ;
  wire [3:0] \oc8051_golden_model_1.n1081 ;
  wire \oc8051_golden_model_1.n1118 ;
  wire \oc8051_golden_model_1.n1146 ;
  wire [8:0] \oc8051_golden_model_1.n1147 ;
  wire [8:0] \oc8051_golden_model_1.n1148 ;
  wire [7:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1150 ;
  wire \oc8051_golden_model_1.n1151 ;
  wire [2:0] \oc8051_golden_model_1.n1152 ;
  wire \oc8051_golden_model_1.n1153 ;
  wire [1:0] \oc8051_golden_model_1.n1154 ;
  wire [7:0] \oc8051_golden_model_1.n1155 ;
  wire [15:0] \oc8051_golden_model_1.n1181 ;
  wire [7:0] \oc8051_golden_model_1.n1183 ;
  wire [8:0] \oc8051_golden_model_1.n1185 ;
  wire [8:0] \oc8051_golden_model_1.n1189 ;
  wire \oc8051_golden_model_1.n1190 ;
  wire [3:0] \oc8051_golden_model_1.n1191 ;
  wire [4:0] \oc8051_golden_model_1.n1192 ;
  wire [4:0] \oc8051_golden_model_1.n1196 ;
  wire \oc8051_golden_model_1.n1197 ;
  wire [8:0] \oc8051_golden_model_1.n1198 ;
  wire \oc8051_golden_model_1.n1206 ;
  wire [7:0] \oc8051_golden_model_1.n1207 ;
  wire [8:0] \oc8051_golden_model_1.n1211 ;
  wire \oc8051_golden_model_1.n1212 ;
  wire [4:0] \oc8051_golden_model_1.n1217 ;
  wire \oc8051_golden_model_1.n1218 ;
  wire \oc8051_golden_model_1.n1226 ;
  wire [7:0] \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1229 ;
  wire [8:0] \oc8051_golden_model_1.n1231 ;
  wire \oc8051_golden_model_1.n1232 ;
  wire [3:0] \oc8051_golden_model_1.n1233 ;
  wire [4:0] \oc8051_golden_model_1.n1234 ;
  wire [4:0] \oc8051_golden_model_1.n1236 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [7:0] \oc8051_golden_model_1.n1246 ;
  wire [8:0] \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1257 ;
  wire [7:0] \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [4:0] \oc8051_golden_model_1.n1278 ;
  wire \oc8051_golden_model_1.n1279 ;
  wire [7:0] \oc8051_golden_model_1.n1280 ;
  wire [8:0] \oc8051_golden_model_1.n1282 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1290 ;
  wire [7:0] \oc8051_golden_model_1.n1291 ;
  wire [7:0] \oc8051_golden_model_1.n1292 ;
  wire [8:0] \oc8051_golden_model_1.n1295 ;
  wire [8:0] \oc8051_golden_model_1.n1296 ;
  wire [7:0] \oc8051_golden_model_1.n1297 ;
  wire \oc8051_golden_model_1.n1298 ;
  wire [7:0] \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [8:0] \oc8051_golden_model_1.n1303 ;
  wire [8:0] \oc8051_golden_model_1.n1305 ;
  wire \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1307 ;
  wire [4:0] \oc8051_golden_model_1.n1309 ;
  wire \oc8051_golden_model_1.n1310 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire [7:0] \oc8051_golden_model_1.n1318 ;
  wire [8:0] \oc8051_golden_model_1.n1322 ;
  wire \oc8051_golden_model_1.n1323 ;
  wire [4:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire [7:0] \oc8051_golden_model_1.n1334 ;
  wire [8:0] \oc8051_golden_model_1.n1338 ;
  wire \oc8051_golden_model_1.n1339 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire [7:0] \oc8051_golden_model_1.n1350 ;
  wire [8:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [4:0] \oc8051_golden_model_1.n1357 ;
  wire \oc8051_golden_model_1.n1358 ;
  wire \oc8051_golden_model_1.n1365 ;
  wire [7:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1520 ;
  wire [6:0] \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [3:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire [7:0] \oc8051_golden_model_1.n1555 ;
  wire [7:0] \oc8051_golden_model_1.n1680 ;
  wire \oc8051_golden_model_1.n1683 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire \oc8051_golden_model_1.n1691 ;
  wire [7:0] \oc8051_golden_model_1.n1692 ;
  wire \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1698 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire \oc8051_golden_model_1.n1709 ;
  wire \oc8051_golden_model_1.n1711 ;
  wire \oc8051_golden_model_1.n1717 ;
  wire [7:0] \oc8051_golden_model_1.n1718 ;
  wire \oc8051_golden_model_1.n1722 ;
  wire \oc8051_golden_model_1.n1724 ;
  wire \oc8051_golden_model_1.n1730 ;
  wire [7:0] \oc8051_golden_model_1.n1731 ;
  wire \oc8051_golden_model_1.n1733 ;
  wire [7:0] \oc8051_golden_model_1.n1734 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire [15:0] \oc8051_golden_model_1.n1739 ;
  wire \oc8051_golden_model_1.n1745 ;
  wire [7:0] \oc8051_golden_model_1.n1746 ;
  wire \oc8051_golden_model_1.n1749 ;
  wire [7:0] \oc8051_golden_model_1.n1750 ;
  wire \oc8051_golden_model_1.n1765 ;
  wire [7:0] \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1771 ;
  wire [7:0] \oc8051_golden_model_1.n1772 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire [7:0] \oc8051_golden_model_1.n1778 ;
  wire \oc8051_golden_model_1.n1783 ;
  wire [7:0] \oc8051_golden_model_1.n1784 ;
  wire \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [7:0] \oc8051_golden_model_1.n1791 ;
  wire [3:0] \oc8051_golden_model_1.n1792 ;
  wire [7:0] \oc8051_golden_model_1.n1793 ;
  wire [7:0] \oc8051_golden_model_1.n1828 ;
  wire \oc8051_golden_model_1.n1847 ;
  wire [7:0] \oc8051_golden_model_1.n1848 ;
  wire [7:0] \oc8051_golden_model_1.n1852 ;
  wire [3:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1854 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_42355_, rst);
  not (_18776_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_18787_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18798_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18787_);
  and (_18809_, _18798_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_18820_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18787_);
  and (_18831_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18787_);
  nor (_18842_, _18831_, _18820_);
  and (_18853_, _18842_, _18809_);
  nor (_18864_, _18853_, _18776_);
  and (_18875_, _18776_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18886_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_18897_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18886_);
  nor (_18908_, _18897_, _18875_);
  not (_18919_, _18908_);
  and (_18930_, _18919_, _18853_);
  or (_18941_, _18930_, _18864_);
  and (_22126_, _18941_, _42355_);
  nor (_18962_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_18973_, _18962_);
  and (_18984_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_18995_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_19006_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_19017_, _19006_);
  not (_19028_, _18897_);
  nor (_19039_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_19050_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_19061_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _19050_);
  nor (_19072_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_19082_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_19093_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _19082_);
  nor (_19104_, _19093_, _19072_);
  nor (_19115_, _19104_, _19061_);
  not (_19126_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_19137_, _19061_, _19126_);
  nor (_19148_, _19137_, _19115_);
  and (_19159_, _19148_, _19039_);
  not (_19170_, _19159_);
  and (_19181_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19192_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_19203_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_19214_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _19203_);
  and (_19225_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_19236_, _19225_, _19192_);
  and (_19247_, _19236_, _19170_);
  nor (_19258_, _19247_, _19028_);
  not (_19269_, _18875_);
  nor (_19280_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_19291_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _19082_);
  nor (_19302_, _19291_, _19280_);
  nor (_19313_, _19302_, _19061_);
  not (_19324_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_19335_, _19061_, _19324_);
  nor (_19346_, _19335_, _19313_);
  and (_19357_, _19346_, _19039_);
  not (_19368_, _19357_);
  and (_19379_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_19390_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_19401_, _19390_, _19379_);
  and (_19411_, _19401_, _19368_);
  nor (_19422_, _19411_, _19269_);
  nor (_19433_, _19422_, _19258_);
  nor (_19444_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_19455_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _19082_);
  nor (_19466_, _19455_, _19444_);
  nor (_19477_, _19466_, _19061_);
  not (_19488_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_19498_, _19061_, _19488_);
  nor (_19509_, _19498_, _19477_);
  and (_19520_, _19509_, _19039_);
  not (_19531_, _19520_);
  and (_19542_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_19553_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_19564_, _19553_, _19542_);
  and (_19574_, _19564_, _19531_);
  nor (_19585_, _19574_, _18919_);
  nor (_19596_, _19585_, _18962_);
  and (_19607_, _19596_, _19433_);
  nor (_19618_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_19629_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _19082_);
  nor (_19640_, _19629_, _19618_);
  nor (_19651_, _19640_, _19061_);
  not (_19661_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_19672_, _19061_, _19661_);
  nor (_19683_, _19672_, _19651_);
  and (_19694_, _19683_, _19039_);
  not (_19705_, _19694_);
  and (_19716_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_19727_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_19738_, _19727_, _19716_);
  and (_19748_, _19738_, _19705_);
  and (_19770_, _19748_, _18962_);
  nor (_19782_, _19770_, _19607_);
  not (_19794_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19806_, _19794_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19818_, _19806_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19830_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_19841_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19842_, _19841_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19853_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_19864_, _19853_, _19830_);
  nor (_19875_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19886_, _19875_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_19897_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_19908_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_19918_, _19806_, _19908_);
  and (_19929_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_19940_, _19929_, _19897_);
  and (_19951_, _19940_, _19864_);
  and (_19962_, _19875_, _19794_);
  and (_19973_, _19962_, _19683_);
  and (_19984_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_19995_, _19984_, _19908_);
  and (_20005_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_20016_, _19984_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_20027_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_20038_, _20027_, _20005_);
  not (_20049_, _20038_);
  nor (_20060_, _20049_, _19973_);
  and (_20071_, _20060_, _19951_);
  not (_20081_, _20071_);
  and (_20092_, _20081_, _19782_);
  not (_20103_, _20092_);
  nor (_20114_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_20125_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _19082_);
  nor (_20136_, _20125_, _20114_);
  nor (_20147_, _20136_, _19061_);
  not (_20158_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_20168_, _19061_, _20158_);
  nor (_20179_, _20168_, _20147_);
  and (_20190_, _20179_, _19039_);
  not (_20201_, _20190_);
  and (_20212_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_20223_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_20234_, _20223_, _20212_);
  and (_20245_, _20234_, _20201_);
  nor (_20255_, _20245_, _19028_);
  nor (_20266_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_20277_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _19082_);
  nor (_20288_, _20277_, _20266_);
  nor (_20299_, _20288_, _19061_);
  not (_20310_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_20321_, _19061_, _20310_);
  nor (_20332_, _20321_, _20299_);
  and (_20342_, _20332_, _19039_);
  not (_20353_, _20342_);
  and (_20364_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_20375_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_20386_, _20375_, _20364_);
  and (_20397_, _20386_, _20353_);
  nor (_20408_, _20397_, _19269_);
  nor (_20418_, _20408_, _20255_);
  nor (_20429_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_20440_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _19082_);
  nor (_20451_, _20440_, _20429_);
  nor (_20462_, _20451_, _19061_);
  not (_20473_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_20484_, _19061_, _20473_);
  nor (_20495_, _20484_, _20462_);
  and (_20505_, _20495_, _19039_);
  not (_20516_, _20505_);
  and (_20527_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_20538_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_20549_, _20538_, _20527_);
  and (_20560_, _20549_, _20516_);
  nor (_20571_, _20560_, _18919_);
  nor (_20582_, _20571_, _18962_);
  and (_20592_, _20582_, _20418_);
  nor (_20603_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_20614_, _19082_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_20625_, _20614_, _20603_);
  nor (_20636_, _20625_, _19061_);
  not (_20647_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_20658_, _19061_, _20647_);
  nor (_20678_, _20658_, _20636_);
  and (_20689_, _20678_, _19039_);
  not (_20690_, _20689_);
  and (_20701_, _19181_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20722_, _19214_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_20733_, _20722_, _20701_);
  and (_20734_, _20733_, _20690_);
  and (_20755_, _20734_, _18962_);
  nor (_20765_, _20755_, _20592_);
  and (_20766_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_20777_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_20788_, _20777_, _20766_);
  and (_20799_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_20820_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_20821_, _20820_, _20799_);
  and (_20832_, _20821_, _20788_);
  and (_20843_, _20678_, _19962_);
  and (_20854_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_20864_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_20875_, _20864_, _20854_);
  not (_20886_, _20875_);
  nor (_20897_, _20886_, _20843_);
  and (_20908_, _20897_, _20832_);
  not (_20919_, _20908_);
  and (_20930_, _20919_, _20765_);
  and (_20950_, _20930_, _20103_);
  not (_20951_, _20950_);
  and (_20962_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_20973_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_20984_, _20973_, _20962_);
  and (_20995_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_21006_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_21017_, _21006_, _20995_);
  and (_21028_, _21017_, _20984_);
  and (_21039_, _20332_, _19962_);
  and (_21049_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_21060_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_21071_, _21060_, _21049_);
  not (_21082_, _21071_);
  nor (_21093_, _21082_, _21039_);
  and (_21104_, _21093_, _21028_);
  not (_21125_, _21104_);
  and (_21126_, _21125_, _20765_);
  and (_21136_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_21147_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_21158_, _21147_, _21136_);
  and (_21169_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_21180_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_21191_, _21180_, _21169_);
  and (_21202_, _21191_, _21158_);
  and (_21213_, _19962_, _19346_);
  and (_21224_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_21234_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_21245_, _21234_, _21224_);
  not (_21256_, _21245_);
  nor (_21267_, _21256_, _21213_);
  and (_21278_, _21267_, _21202_);
  not (_21289_, _21278_);
  and (_21300_, _21289_, _19782_);
  and (_21320_, _21300_, _21126_);
  and (_21321_, _21320_, _20081_);
  nor (_21332_, _21320_, _20092_);
  nor (_21343_, _21332_, _21321_);
  and (_21354_, _21343_, _21126_);
  and (_21365_, _20930_, _20092_);
  and (_21376_, _20765_, _20081_);
  and (_21387_, _20919_, _19782_);
  nor (_21398_, _21387_, _21376_);
  nor (_21409_, _21398_, _21365_);
  and (_21419_, _21409_, _21354_);
  nor (_21430_, _21409_, _21354_);
  nor (_21441_, _21430_, _21419_);
  and (_21452_, _21441_, _21321_);
  nor (_21463_, _21452_, _21419_);
  nor (_21474_, _21463_, _20951_);
  and (_21485_, _21463_, _20951_);
  nor (_21496_, _21485_, _21474_);
  not (_21506_, _21496_);
  and (_21517_, _21289_, _20765_);
  and (_21528_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_21539_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_21550_, _21539_, _21528_);
  and (_21561_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_21572_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_21583_, _21572_, _21561_);
  and (_21594_, _21583_, _21550_);
  and (_21604_, _20179_, _19962_);
  and (_21615_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_21626_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_21637_, _21626_, _21615_);
  not (_21648_, _21637_);
  nor (_21669_, _21648_, _21604_);
  and (_21670_, _21669_, _21594_);
  not (_21681_, _21670_);
  and (_21691_, _21681_, _19782_);
  and (_21702_, _21691_, _21517_);
  and (_21713_, _21125_, _19782_);
  nor (_21724_, _21713_, _21517_);
  nor (_21735_, _21724_, _21320_);
  and (_21746_, _21735_, _21702_);
  nor (_21757_, _21126_, _20092_);
  nor (_21778_, _21757_, _21354_);
  and (_21779_, _21778_, _21746_);
  nor (_21789_, _21441_, _21321_);
  nor (_21800_, _21789_, _21452_);
  and (_21811_, _21800_, _21779_);
  nor (_21822_, _21800_, _21779_);
  nor (_21833_, _21822_, _21811_);
  not (_21844_, _21833_);
  and (_21855_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_21866_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_21876_, _21866_, _21855_);
  and (_21887_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_21898_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_21909_, _21898_, _21887_);
  and (_21920_, _21909_, _21876_);
  and (_21931_, _20495_, _19962_);
  and (_21942_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_21952_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_21963_, _21952_, _21942_);
  not (_21974_, _21963_);
  nor (_21985_, _21974_, _21931_);
  and (_21996_, _21985_, _21920_);
  not (_22007_, _21996_);
  and (_22018_, _22007_, _20765_);
  and (_22029_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_22039_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_22050_, _22039_, _22029_);
  and (_22061_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_22072_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_22083_, _22072_, _22061_);
  and (_22094_, _22083_, _22050_);
  and (_22105_, _19962_, _19148_);
  and (_22116_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_22127_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_22138_, _22127_, _22116_);
  not (_22149_, _22138_);
  nor (_22160_, _22149_, _22105_);
  and (_22171_, _22160_, _22094_);
  not (_22182_, _22171_);
  and (_22193_, _22182_, _19782_);
  and (_22204_, _22193_, _22018_);
  and (_22224_, _22007_, _19782_);
  not (_22225_, _22224_);
  and (_22236_, _22182_, _20765_);
  and (_22247_, _22236_, _22225_);
  and (_22258_, _22247_, _21691_);
  nor (_22269_, _22258_, _22204_);
  and (_22280_, _21681_, _20765_);
  nor (_22290_, _22280_, _21300_);
  nor (_22301_, _22290_, _21702_);
  not (_22312_, _22301_);
  nor (_22323_, _22312_, _22269_);
  nor (_22334_, _21735_, _21702_);
  nor (_22345_, _22334_, _21746_);
  and (_22356_, _22345_, _22323_);
  nor (_22367_, _21778_, _21746_);
  nor (_22377_, _22367_, _21779_);
  and (_22388_, _22377_, _22356_);
  and (_22399_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_22410_, _19842_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_22421_, _22410_, _22399_);
  and (_22432_, _19886_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_22443_, _19918_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_22454_, _22443_, _22432_);
  and (_22464_, _22454_, _22421_);
  and (_22475_, _19962_, _19509_);
  and (_22486_, _20016_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_22497_, _19995_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_22518_, _22497_, _22486_);
  not (_22519_, _22518_);
  nor (_22530_, _22519_, _22475_);
  and (_22540_, _22530_, _22464_);
  not (_22551_, _22540_);
  and (_22562_, _22551_, _20765_);
  and (_22573_, _22562_, _22224_);
  nor (_22584_, _22193_, _22018_);
  nor (_22595_, _22584_, _22204_);
  and (_22606_, _22595_, _22573_);
  nor (_22626_, _22247_, _21691_);
  nor (_22627_, _22626_, _22258_);
  and (_22638_, _22627_, _22606_);
  and (_22649_, _22312_, _22269_);
  nor (_22660_, _22649_, _22323_);
  and (_22671_, _22660_, _22638_);
  nor (_22682_, _22345_, _22323_);
  nor (_22693_, _22682_, _22356_);
  and (_22703_, _22693_, _22671_);
  nor (_22714_, _22377_, _22356_);
  nor (_22725_, _22714_, _22388_);
  and (_22736_, _22725_, _22703_);
  nor (_22747_, _22736_, _22388_);
  nor (_22758_, _22747_, _21844_);
  nor (_22769_, _22758_, _21811_);
  nor (_22780_, _22769_, _21506_);
  or (_22790_, _22780_, _21365_);
  nor (_22801_, _22790_, _21474_);
  nor (_22812_, _22801_, _19017_);
  and (_22823_, _22801_, _19017_);
  nor (_22844_, _22823_, _22812_);
  not (_22845_, _22844_);
  and (_22856_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_22867_, _22769_, _21506_);
  nor (_22877_, _22867_, _22780_);
  and (_22888_, _22877_, _22856_);
  and (_22899_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_22910_, _22747_, _21844_);
  nor (_22921_, _22910_, _22758_);
  and (_22932_, _22921_, _22899_);
  nor (_22943_, _22921_, _22899_);
  nor (_22953_, _22943_, _22932_);
  not (_22964_, _22953_);
  and (_22975_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_22986_, _22725_, _22703_);
  nor (_22997_, _22986_, _22736_);
  and (_23008_, _22997_, _22975_);
  nor (_23019_, _22997_, _22975_);
  nor (_23030_, _23019_, _23008_);
  and (_23040_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_23051_, _22693_, _22671_);
  nor (_23062_, _23051_, _22703_);
  and (_23073_, _23062_, _23040_);
  nor (_23084_, _23062_, _23040_);
  nor (_23105_, _23084_, _23073_);
  not (_23106_, _23105_);
  and (_23117_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_23128_, _22660_, _22638_);
  nor (_23139_, _23128_, _22671_);
  and (_23149_, _23139_, _23117_);
  and (_23160_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_23171_, _22627_, _22606_);
  nor (_23182_, _23171_, _22638_);
  and (_23193_, _23182_, _23160_);
  and (_23204_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_23215_, _22595_, _22573_);
  nor (_23226_, _23215_, _22606_);
  and (_23237_, _23226_, _23204_);
  nor (_23248_, _23182_, _23160_);
  nor (_23258_, _23248_, _23193_);
  and (_23269_, _23258_, _23237_);
  nor (_23280_, _23269_, _23193_);
  not (_23291_, _23280_);
  nor (_23302_, _23139_, _23117_);
  nor (_23313_, _23302_, _23149_);
  and (_23324_, _23313_, _23291_);
  nor (_23335_, _23324_, _23149_);
  nor (_23346_, _23335_, _23106_);
  nor (_23357_, _23346_, _23073_);
  not (_23367_, _23357_);
  and (_23388_, _23367_, _23030_);
  nor (_23389_, _23388_, _23008_);
  nor (_23400_, _23389_, _22964_);
  nor (_23411_, _23400_, _22932_);
  nor (_23422_, _22877_, _22856_);
  nor (_23433_, _23422_, _22888_);
  not (_23444_, _23433_);
  nor (_23455_, _23444_, _23411_);
  nor (_23466_, _23455_, _22888_);
  nor (_23476_, _23466_, _22845_);
  nor (_23487_, _23476_, _22812_);
  not (_23498_, _23487_);
  and (_23509_, _23498_, _18995_);
  and (_23520_, _23509_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_23531_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_23542_, _23531_, _23520_);
  and (_23553_, _23542_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_23564_, _23553_, _18984_);
  not (_23575_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_23585_, _18962_, _23575_);
  or (_23596_, _23585_, _23564_);
  nand (_23607_, _23564_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and (_23618_, _23607_, _23596_);
  and (_24284_, _23618_, _42355_);
  nor (_23639_, _18853_, _18886_);
  and (_23650_, _18853_, _18886_);
  or (_23661_, _23650_, _23639_);
  and (_02358_, _23661_, _42355_);
  and (_23682_, _22551_, _19782_);
  and (_02546_, _23682_, _42355_);
  nor (_23702_, _22562_, _22224_);
  nor (_23713_, _23702_, _22573_);
  and (_02702_, _23713_, _42355_);
  nor (_23734_, _23226_, _23204_);
  nor (_23745_, _23734_, _23237_);
  and (_02884_, _23745_, _42355_);
  nor (_23766_, _23258_, _23237_);
  nor (_23777_, _23766_, _23269_);
  and (_03126_, _23777_, _42355_);
  nor (_23797_, _23313_, _23291_);
  nor (_23818_, _23797_, _23324_);
  and (_03330_, _23818_, _42355_);
  and (_23829_, _23335_, _23106_);
  nor (_23840_, _23829_, _23346_);
  and (_03531_, _23840_, _42355_);
  nor (_23861_, _23367_, _23030_);
  nor (_23871_, _23861_, _23388_);
  and (_03732_, _23871_, _42355_);
  and (_23892_, _23389_, _22964_);
  nor (_23903_, _23892_, _23400_);
  and (_03929_, _23903_, _42355_);
  and (_23924_, _23444_, _23411_);
  nor (_23935_, _23924_, _23455_);
  and (_04027_, _23935_, _42355_);
  and (_23955_, _23466_, _22845_);
  nor (_23966_, _23955_, _23476_);
  and (_04126_, _23966_, _42355_);
  nor (_23997_, _23498_, _18995_);
  nor (_23998_, _23997_, _23509_);
  and (_04226_, _23998_, _42355_);
  and (_24019_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_24030_, _24019_, _23509_);
  nor (_24040_, _24030_, _23520_);
  and (_04325_, _24040_, _42355_);
  nor (_24061_, _23531_, _23520_);
  nor (_24072_, _24061_, _23542_);
  and (_04419_, _24072_, _42355_);
  and (_24093_, _18973_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_24104_, _24093_, _23542_);
  nor (_24115_, _24104_, _23553_);
  and (_04517_, _24115_, _42355_);
  nor (_24135_, _23553_, _18984_);
  nor (_24146_, _24135_, _23564_);
  and (_04616_, _24146_, _42355_);
  and (_24167_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18787_);
  nor (_24178_, _24167_, _18798_);
  not (_24189_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_24199_, _18820_, _24189_);
  and (_24210_, _24199_, _24178_);
  and (_24221_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24232_, _24221_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24243_, _24221_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24254_, _24243_, _24232_);
  and (_00925_, _24254_, _42355_);
  and (_00955_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _42355_);
  not (_24285_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_24296_, _20560_, _24285_);
  and (_24307_, _20245_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24318_, _24307_, _24296_);
  nor (_24329_, _24318_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24340_, _20397_, _24285_);
  and (_24351_, _20734_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24362_, _24351_, _24340_);
  and (_24372_, _24362_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24383_, _24372_, _24329_);
  nor (_24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24405_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and (_24416_, _24394_, _20908_);
  nor (_24427_, _24416_, _24405_);
  not (_24438_, _24427_);
  and (_24448_, _19574_, _24285_);
  and (_24459_, _19247_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24470_, _24459_, _24448_);
  nor (_24481_, _24470_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24492_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24503_, _19411_, _24285_);
  and (_24524_, _19748_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24525_, _24524_, _24503_);
  nor (_24535_, _24525_, _24492_);
  nor (_24546_, _24535_, _24481_);
  nor (_24557_, _24546_, _24438_);
  and (_24568_, _24546_, _24438_);
  nor (_24579_, _24568_, _24557_);
  and (_24590_, _24394_, _20071_);
  nor (_24601_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_24612_, _24601_, _24590_);
  not (_24622_, _24612_);
  nor (_24633_, _20560_, _24285_);
  nor (_24644_, _24633_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24655_, _20245_, _24285_);
  and (_24666_, _20397_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24677_, _24666_, _24655_);
  nor (_24688_, _24677_, _24492_);
  nor (_24698_, _24688_, _24644_);
  nor (_24709_, _24698_, _24622_);
  and (_24720_, _24698_, _24622_);
  nor (_24731_, _24720_, _24709_);
  not (_24742_, _24731_);
  and (_24753_, _24394_, _21104_);
  nor (_24764_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor (_24775_, _24764_, _24753_);
  not (_24785_, _24775_);
  nor (_24796_, _19574_, _24285_);
  nor (_24807_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24818_, _19247_, _24285_);
  and (_24829_, _19411_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24840_, _24829_, _24818_);
  nor (_24851_, _24840_, _24492_);
  nor (_24862_, _24851_, _24807_);
  nor (_24872_, _24862_, _24785_);
  and (_24883_, _24862_, _24785_);
  nor (_24894_, _24883_, _24872_);
  not (_24905_, _24894_);
  and (_24916_, _24318_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24927_, _24916_);
  nor (_24938_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_24948_, _24394_, _21278_);
  nor (_24959_, _24948_, _24938_);
  and (_24970_, _24959_, _24927_);
  and (_24981_, _24470_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24992_, _24981_);
  and (_25003_, _24394_, _21670_);
  nor (_25014_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_25025_, _25014_, _25003_);
  and (_25036_, _25025_, _24992_);
  nor (_25047_, _25025_, _24992_);
  nor (_25068_, _25047_, _25036_);
  not (_25069_, _25068_);
  and (_25080_, _24633_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25091_, _25080_);
  and (_25102_, _24394_, _22171_);
  nor (_25113_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_25124_, _25113_, _25102_);
  and (_25135_, _25124_, _25091_);
  and (_25146_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_25157_, _25146_);
  nor (_25168_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_25179_, _24394_, _21996_);
  nor (_25189_, _25179_, _25168_);
  nor (_25200_, _25189_, _25157_);
  not (_25211_, _25200_);
  nor (_25222_, _25124_, _25091_);
  nor (_25233_, _25222_, _25135_);
  and (_25244_, _25233_, _25211_);
  nor (_25255_, _25244_, _25135_);
  nor (_25266_, _25255_, _25069_);
  nor (_25277_, _25266_, _25036_);
  nor (_25288_, _24959_, _24927_);
  nor (_25299_, _25288_, _24970_);
  not (_25310_, _25299_);
  nor (_25331_, _25310_, _25277_);
  nor (_25332_, _25331_, _24970_);
  nor (_25343_, _25332_, _24905_);
  nor (_25354_, _25343_, _24872_);
  nor (_25365_, _25354_, _24742_);
  nor (_25376_, _25365_, _24709_);
  not (_25387_, _25376_);
  and (_25398_, _25387_, _24579_);
  or (_25409_, _25398_, _24557_);
  and (_25420_, _20734_, _19748_);
  or (_25431_, _25420_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_25442_, _24525_);
  and (_25453_, _24362_, _25442_);
  nor (_25464_, _24840_, _24677_);
  and (_25475_, _25464_, _25453_);
  or (_25486_, _25475_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_25497_, _25486_, _25431_);
  and (_25508_, _25497_, _25409_);
  and (_25519_, _25508_, _24383_);
  nor (_25530_, _25387_, _24579_);
  or (_25541_, _25530_, _25398_);
  and (_25552_, _25541_, _25519_);
  nor (_25563_, _25519_, _24427_);
  nor (_25573_, _25563_, _25552_);
  not (_25584_, _25573_);
  and (_25595_, _25573_, _24383_);
  not (_25606_, _24546_);
  and (_25617_, _25354_, _24742_);
  or (_25638_, _25617_, _25365_);
  and (_25639_, _25638_, _25519_);
  nor (_25650_, _25519_, _24612_);
  nor (_25661_, _25650_, _25639_);
  and (_25672_, _25661_, _25606_);
  nor (_25683_, _25661_, _25606_);
  nor (_25694_, _25683_, _25672_);
  not (_25705_, _25694_);
  not (_25716_, _24698_);
  nor (_25727_, _25519_, _24785_);
  and (_25738_, _25332_, _24905_);
  nor (_25749_, _25738_, _25343_);
  and (_25760_, _25749_, _25519_);
  or (_25771_, _25760_, _25727_);
  and (_25782_, _25771_, _25716_);
  nor (_25793_, _25771_, _25716_);
  not (_25804_, _24862_);
  and (_25815_, _25310_, _25277_);
  or (_25826_, _25815_, _25331_);
  and (_25837_, _25826_, _25519_);
  nor (_25848_, _25519_, _24959_);
  nor (_25859_, _25848_, _25837_);
  and (_25870_, _25859_, _25804_);
  and (_25881_, _25255_, _25069_);
  nor (_25892_, _25881_, _25266_);
  not (_25903_, _25892_);
  and (_25914_, _25903_, _25519_);
  nor (_25924_, _25519_, _25025_);
  nor (_25935_, _25924_, _25914_);
  and (_25946_, _25935_, _24927_);
  nor (_25967_, _25935_, _24927_);
  nor (_25968_, _25967_, _25946_);
  not (_25979_, _25968_);
  nor (_25990_, _25233_, _25211_);
  nor (_26001_, _25990_, _25244_);
  not (_26012_, _26001_);
  and (_26023_, _26012_, _25519_);
  nor (_26034_, _25519_, _25124_);
  nor (_26045_, _26034_, _26023_);
  and (_26056_, _26045_, _24992_);
  not (_26067_, _25189_);
  and (_26078_, _25519_, _25146_);
  or (_26089_, _26078_, _26067_);
  nand (_26100_, _25519_, _25146_);
  or (_26111_, _26100_, _25189_);
  and (_26122_, _26111_, _26089_);
  nor (_26133_, _26122_, _25080_);
  and (_26144_, _26122_, _25080_);
  nor (_26155_, _26144_, _26133_);
  and (_26166_, _24394_, _22540_);
  nor (_26177_, _24394_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_26188_, _26177_, _26166_);
  nor (_26199_, _26188_, _25157_);
  not (_26210_, _26199_);
  and (_26221_, _26210_, _26155_);
  nor (_26232_, _26221_, _26133_);
  nor (_26243_, _26045_, _24992_);
  nor (_26254_, _26243_, _26056_);
  not (_26264_, _26254_);
  nor (_26275_, _26264_, _26232_);
  nor (_26286_, _26275_, _26056_);
  nor (_26297_, _26286_, _25979_);
  nor (_26308_, _26297_, _25946_);
  nor (_26319_, _25859_, _25804_);
  nor (_26330_, _26319_, _25870_);
  not (_26341_, _26330_);
  nor (_26352_, _26341_, _26308_);
  nor (_26363_, _26352_, _25870_);
  nor (_26374_, _26363_, _25793_);
  nor (_26385_, _26374_, _25782_);
  nor (_26396_, _26385_, _25705_);
  or (_26407_, _26396_, _25672_);
  or (_26418_, _26407_, _25595_);
  and (_26429_, _26418_, _25497_);
  nor (_26450_, _26429_, _25584_);
  and (_26451_, _25595_, _25497_);
  and (_26462_, _26451_, _26407_);
  or (_26473_, _26462_, _26450_);
  and (_00974_, _26473_, _42355_);
  or (_26494_, _25573_, _24383_);
  and (_26505_, _26494_, _26429_);
  and (_02839_, _26505_, _42355_);
  and (_02851_, _25519_, _42355_);
  and (_02873_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _42355_);
  and (_02897_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _42355_);
  and (_02919_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _42355_);
  or (_26566_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_26577_, _24221_, rst);
  and (_02931_, _26577_, _26566_);
  not (_26597_, _26188_);
  and (_26608_, _26505_, _25146_);
  nor (_26619_, _26608_, _26597_);
  and (_26630_, _26608_, _26597_);
  or (_26641_, _26630_, _26619_);
  and (_02943_, _26641_, _42355_);
  nor (_26672_, _26505_, _26122_);
  nor (_26673_, _26210_, _26155_);
  nor (_26684_, _26673_, _26221_);
  and (_26695_, _26684_, _26505_);
  or (_26706_, _26695_, _26672_);
  and (_02957_, _26706_, _42355_);
  and (_26727_, _26264_, _26232_);
  or (_26738_, _26727_, _26275_);
  nand (_26749_, _26738_, _26505_);
  or (_26760_, _26505_, _26045_);
  and (_26771_, _26760_, _26749_);
  and (_02971_, _26771_, _42355_);
  and (_26792_, _26286_, _25979_);
  or (_26803_, _26792_, _26297_);
  nand (_26814_, _26803_, _26505_);
  or (_26825_, _26505_, _25935_);
  and (_26836_, _26825_, _26814_);
  and (_02984_, _26836_, _42355_);
  and (_26857_, _26341_, _26308_);
  or (_26868_, _26857_, _26352_);
  nand (_26879_, _26868_, _26505_);
  or (_26890_, _26505_, _25859_);
  and (_26901_, _26890_, _26879_);
  and (_02998_, _26901_, _42355_);
  or (_26922_, _25793_, _25782_);
  and (_26933_, _26922_, _26363_);
  nor (_26943_, _26922_, _26363_);
  or (_26954_, _26943_, _26933_);
  nand (_26965_, _26954_, _26505_);
  or (_26976_, _26505_, _25771_);
  and (_26987_, _26976_, _26965_);
  and (_03011_, _26987_, _42355_);
  and (_27008_, _26385_, _25705_);
  or (_27019_, _27008_, _26396_);
  nand (_27030_, _27019_, _26505_);
  or (_27041_, _26505_, _25661_);
  and (_27052_, _27041_, _27030_);
  and (_03023_, _27052_, _42355_);
  not (_27073_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27084_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18787_);
  and (_27095_, _27084_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_27106_, _27095_, _27073_);
  and (_27117_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27128_, _27117_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_27139_, _27117_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_27150_, _27139_, _27128_);
  and (_27161_, _27150_, _27106_);
  not (_27172_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_27183_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18787_);
  and (_27194_, _27183_, _27073_);
  and (_27205_, _27194_, _27172_);
  and (_27216_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_27227_, _27216_, _27161_);
  not (_27248_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_27249_, _27084_, _27248_);
  and (_27260_, _27249_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27271_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_27282_, _27249_, _27073_);
  and (_27292_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_27303_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27314_, _27303_, _18787_);
  nor (_27325_, _27314_, _27084_);
  and (_27336_, _27325_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_27347_, _27336_, _27292_);
  nor (_27358_, _27347_, _27271_);
  and (_27369_, _27358_, _27227_);
  nor (_27380_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_27391_, _27380_, _27117_);
  and (_27402_, _27391_, _27106_);
  and (_27413_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_27424_, _27413_, _27402_);
  and (_27435_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_27446_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_27457_, _27325_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_27468_, _27457_, _27446_);
  nor (_27479_, _27468_, _27435_);
  and (_27490_, _27479_, _27424_);
  and (_27501_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_27512_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_27523_, _27512_, _27501_);
  and (_27534_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_27545_, _27534_);
  not (_27556_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_27567_, _27106_, _27556_);
  and (_27578_, _27325_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_27589_, _27578_, _27567_);
  and (_27600_, _27589_, _27545_);
  and (_27611_, _27600_, _27523_);
  and (_27622_, _27611_, _27490_);
  and (_27633_, _27622_, _27369_);
  and (_27643_, _27128_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_27654_, _27643_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_27665_, _27654_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_27676_, _27665_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_27687_, _27676_);
  not (_27698_, _27106_);
  nor (_27709_, _27665_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_27720_, _27709_, _27698_);
  and (_27731_, _27720_, _27687_);
  not (_27742_, _27731_);
  and (_27753_, _27095_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_27764_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_27775_, _27764_, _27753_);
  and (_27786_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_27797_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_27808_, _27797_, _27786_);
  and (_27819_, _27808_, _27775_);
  and (_27830_, _27819_, _27742_);
  nor (_27841_, _27654_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_27852_, _27841_);
  nor (_27863_, _27665_, _27698_);
  and (_27884_, _27863_, _27852_);
  not (_27885_, _27884_);
  and (_27896_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_27907_, _27896_, _27753_);
  and (_27918_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_27929_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_27940_, _27929_, _27918_);
  and (_27950_, _27940_, _27907_);
  and (_27961_, _27950_, _27885_);
  nor (_27972_, _27961_, _27830_);
  not (_27983_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_27994_, _27676_, _27983_);
  and (_28005_, _27676_, _27983_);
  nor (_28016_, _28005_, _27994_);
  nor (_28027_, _28016_, _27698_);
  not (_28038_, _28027_);
  and (_28049_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_28060_, _28049_);
  not (_28071_, _27753_);
  and (_28082_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_28093_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_28104_, _28093_, _28082_);
  and (_28115_, _28104_, _28071_);
  and (_28126_, _28115_, _28060_);
  and (_28137_, _28126_, _28038_);
  not (_28148_, _28137_);
  and (_28159_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_28170_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_28191_, _28170_, _28159_);
  not (_28192_, _27643_);
  nor (_28203_, _27128_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_28214_, _28203_, _27698_);
  and (_28225_, _28214_, _28192_);
  and (_28236_, _27325_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_28247_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_28258_, _28247_, _28236_);
  not (_28268_, _28258_);
  nor (_28279_, _28268_, _28225_);
  and (_28290_, _28279_, _28191_);
  not (_28301_, _28290_);
  and (_28312_, _27260_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_28323_, _28312_, _27753_);
  nor (_28334_, _27643_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_28345_, _28334_, _27698_);
  nor (_28356_, _28345_, _27654_);
  and (_28367_, _27282_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_28378_, _28367_, _28356_);
  and (_28389_, _28378_, _28323_);
  and (_28400_, _27325_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_28411_, _27205_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_28422_, _28411_, _28400_);
  and (_28433_, _28422_, _28389_);
  nor (_28444_, _28433_, _28301_);
  and (_28455_, _28444_, _28148_);
  and (_28466_, _28455_, _27972_);
  nand (_28477_, _28466_, _27633_);
  and (_28488_, _26473_, _24210_);
  not (_28499_, _28488_);
  and (_28510_, _23618_, _18853_);
  not (_28521_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_28542_, _18798_, _28521_);
  and (_28543_, _28542_, _18842_);
  not (_28554_, _28543_);
  nor (_28565_, _20908_, _20734_);
  and (_28575_, _20908_, _20734_);
  nor (_28586_, _28575_, _28565_);
  not (_28597_, _19748_);
  nor (_28608_, _20071_, _28597_);
  nor (_28619_, _20071_, _19748_);
  and (_28630_, _20071_, _19748_);
  nor (_28641_, _28630_, _28619_);
  not (_28652_, _20397_);
  nor (_28663_, _21104_, _28652_);
  nor (_28674_, _21104_, _20397_);
  and (_28685_, _21104_, _20397_);
  nor (_28696_, _28685_, _28674_);
  not (_28707_, _19411_);
  and (_28718_, _21278_, _28707_);
  nor (_28729_, _28718_, _28696_);
  nor (_28740_, _28729_, _28663_);
  nor (_28751_, _28740_, _28641_);
  nor (_28762_, _28751_, _28608_);
  and (_28773_, _28740_, _28641_);
  nor (_28784_, _28773_, _28751_);
  not (_28795_, _28784_);
  and (_28806_, _28718_, _28696_);
  nor (_28817_, _28806_, _28729_);
  not (_28828_, _28817_);
  nor (_28839_, _21278_, _19411_);
  and (_28850_, _21278_, _19411_);
  nor (_28861_, _28850_, _28839_);
  not (_28872_, _28861_);
  and (_28882_, _21670_, _20245_);
  nor (_28893_, _21670_, _20245_);
  nor (_28914_, _28893_, _28882_);
  not (_28915_, _28914_);
  nor (_28926_, _22171_, _19247_);
  and (_28937_, _22171_, _19247_);
  nor (_28948_, _28937_, _28926_);
  nor (_28959_, _21996_, _20560_);
  and (_28970_, _21996_, _20560_);
  nor (_28981_, _28970_, _28959_);
  not (_28992_, _19574_);
  and (_29003_, _22540_, _28992_);
  nor (_29014_, _29003_, _28981_);
  not (_29025_, _20560_);
  nor (_29036_, _21996_, _29025_);
  nor (_29047_, _29036_, _29014_);
  nor (_29058_, _29047_, _28948_);
  not (_29069_, _19247_);
  nor (_29080_, _22171_, _29069_);
  nor (_29091_, _29080_, _29058_);
  nor (_29102_, _29091_, _28915_);
  and (_29113_, _29091_, _28915_);
  nor (_29124_, _29113_, _29102_);
  and (_29135_, _29047_, _28948_);
  nor (_29146_, _29135_, _29058_);
  not (_29157_, _29146_);
  nor (_29168_, _22540_, _19574_);
  and (_29178_, _22540_, _19574_);
  nor (_29189_, _29178_, _29168_);
  not (_29200_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_29211_, _19061_, _29200_);
  not (_29222_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_29233_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29244_, _29233_, _20625_);
  nor (_29255_, _29244_, _29222_);
  nor (_29266_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29277_, _29266_, _19302_);
  not (_29288_, _29277_);
  not (_29299_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29310_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _29299_);
  and (_29321_, _29310_, _20288_);
  not (_29332_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_29343_, _29332_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_29354_, _29343_, _19640_);
  nor (_29365_, _29354_, _29321_);
  and (_29376_, _29365_, _29288_);
  and (_29387_, _29376_, _29255_);
  and (_29398_, _29233_, _20136_);
  nor (_29409_, _29398_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_29420_, _29343_, _19104_);
  not (_29441_, _29420_);
  and (_29442_, _29310_, _20451_);
  and (_29453_, _29266_, _19466_);
  nor (_29464_, _29453_, _29442_);
  and (_29475_, _29464_, _29441_);
  and (_29485_, _29475_, _29409_);
  nor (_29496_, _29485_, _29387_);
  nor (_29507_, _29496_, _19061_);
  nor (_29518_, _29507_, _29211_);
  and (_29529_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_29540_, _29529_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_29551_, _29540_);
  and (_29562_, _29551_, _29518_);
  and (_29573_, _29551_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_29584_, _29573_, _29562_);
  nor (_29595_, _29584_, _29189_);
  and (_29606_, _29003_, _28981_);
  nor (_29617_, _29606_, _29014_);
  not (_29628_, _29617_);
  and (_29639_, _29628_, _29595_);
  and (_29650_, _29639_, _29157_);
  and (_29661_, _29650_, _29124_);
  not (_29672_, _20245_);
  or (_29683_, _21670_, _29672_);
  and (_29694_, _21670_, _29672_);
  or (_29715_, _29091_, _29694_);
  and (_29716_, _29715_, _29683_);
  or (_29727_, _29716_, _29661_);
  and (_29738_, _29727_, _28872_);
  and (_29749_, _29738_, _28828_);
  and (_29760_, _29749_, _28795_);
  nor (_29771_, _29760_, _28762_);
  nor (_29781_, _29771_, _28586_);
  and (_29792_, _29771_, _28586_);
  nor (_29803_, _29792_, _29781_);
  nor (_29814_, _29803_, _28554_);
  not (_29825_, _29814_);
  not (_29836_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_29847_, _24167_, _29836_);
  and (_29858_, _29847_, _18842_);
  not (_29869_, _28586_);
  not (_29879_, _28641_);
  and (_29890_, _28839_, _28696_);
  nor (_29901_, _29890_, _28674_);
  nor (_29912_, _29901_, _29879_);
  not (_29923_, _28948_);
  and (_29934_, _29168_, _28981_);
  nor (_29945_, _29934_, _28959_);
  nor (_29956_, _29945_, _29923_);
  nor (_29967_, _29956_, _28926_);
  nor (_29978_, _29967_, _28914_);
  and (_29989_, _29967_, _28914_);
  nor (_29999_, _29989_, _29978_);
  not (_30010_, _29189_);
  nor (_30021_, _29584_, _30010_);
  and (_30032_, _30021_, _28981_);
  and (_30043_, _29945_, _29923_);
  nor (_30054_, _30043_, _29956_);
  and (_30065_, _30054_, _30032_);
  not (_30076_, _30065_);
  nor (_30087_, _30076_, _29999_);
  nor (_30098_, _29967_, _28882_);
  or (_30108_, _30098_, _28893_);
  or (_30119_, _30108_, _30087_);
  and (_30130_, _30119_, _28861_);
  nor (_30141_, _28839_, _28696_);
  nor (_30152_, _30141_, _29890_);
  and (_30163_, _30152_, _30130_);
  and (_30174_, _29901_, _29879_);
  nor (_30185_, _30174_, _29912_);
  and (_30196_, _30185_, _30163_);
  or (_30207_, _30196_, _29912_);
  nor (_30217_, _30207_, _28619_);
  nor (_30228_, _30217_, _29869_);
  and (_30239_, _30217_, _29869_);
  nor (_30250_, _30239_, _30228_);
  and (_30261_, _30250_, _29858_);
  and (_30272_, _18831_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30283_, _30272_, _28542_);
  nor (_30294_, _22540_, _21996_);
  and (_30305_, _30294_, _22182_);
  and (_30316_, _30305_, _21681_);
  and (_30336_, _30316_, _21289_);
  and (_30337_, _30336_, _21125_);
  and (_30348_, _30337_, _20081_);
  and (_30359_, _30348_, _29584_);
  not (_30370_, _29584_);
  and (_30381_, _21104_, _20071_);
  and (_30392_, _22540_, _21996_);
  and (_30403_, _30392_, _22171_);
  and (_30414_, _30403_, _21670_);
  and (_30425_, _30414_, _21278_);
  and (_30435_, _30425_, _30381_);
  and (_30446_, _30435_, _30370_);
  nor (_30457_, _30446_, _30359_);
  and (_30468_, _30457_, _20908_);
  nor (_30479_, _30457_, _20908_);
  nor (_30490_, _30479_, _30468_);
  and (_30501_, _30490_, _30283_);
  not (_30512_, _20734_);
  nor (_30523_, _29584_, _30512_);
  not (_30534_, _30523_);
  and (_30544_, _29584_, _20908_);
  and (_30555_, _30272_, _18809_);
  not (_30566_, _30555_);
  nor (_30577_, _30566_, _30544_);
  and (_30588_, _30577_, _30534_);
  nor (_30599_, _30588_, _30501_);
  and (_30610_, _29847_, _24199_);
  not (_30621_, _30610_);
  and (_30632_, _22171_, _21996_);
  nor (_30642_, _30632_, _21670_);
  and (_30653_, _30642_, _30610_);
  and (_30664_, _30653_, _21289_);
  nor (_30675_, _30664_, _21125_);
  and (_30686_, _30675_, _20071_);
  nor (_30697_, _30381_, _20908_);
  nor (_30708_, _30697_, _30653_);
  and (_30719_, _30708_, _29584_);
  nor (_30730_, _30719_, _30686_);
  and (_30741_, _30730_, _20908_);
  nor (_30752_, _30730_, _20908_);
  nor (_30762_, _30752_, _30741_);
  nor (_30773_, _30762_, _30621_);
  and (_30784_, _30272_, _29847_);
  not (_30795_, _30784_);
  nor (_30806_, _30795_, _29584_);
  not (_30817_, _30806_);
  not (_30828_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_30839_, _18831_, _30828_);
  and (_30850_, _30839_, _29847_);
  not (_30861_, _30850_);
  nor (_30871_, _30861_, _28575_);
  and (_30882_, _30839_, _24178_);
  and (_30893_, _30882_, _28586_);
  nor (_30904_, _30893_, _30871_);
  and (_30915_, _24199_, _18809_);
  and (_30926_, _30915_, _28565_);
  and (_30937_, _28542_, _24199_);
  and (_30948_, _30937_, _20908_);
  nor (_30959_, _30948_, _30926_);
  and (_30970_, _24178_, _18842_);
  not (_30980_, _30970_);
  nor (_30991_, _30980_, _20908_);
  not (_31002_, _30991_);
  and (_31013_, _30272_, _24178_);
  not (_31024_, _31013_);
  nor (_31046_, _31024_, _22540_);
  and (_31047_, _30839_, _18798_);
  not (_31069_, _31047_);
  nor (_31070_, _31069_, _20071_);
  nor (_31091_, _31070_, _31046_);
  and (_31092_, _31091_, _31002_);
  and (_31114_, _31092_, _30959_);
  and (_31115_, _31114_, _30904_);
  and (_31126_, _31115_, _30817_);
  not (_31137_, _31126_);
  nor (_31148_, _31137_, _30773_);
  and (_31169_, _31148_, _30599_);
  not (_31170_, _31169_);
  nor (_31191_, _31170_, _30261_);
  and (_31192_, _31191_, _29825_);
  not (_31212_, _31192_);
  nor (_31213_, _31212_, _28510_);
  and (_31234_, _31213_, _28499_);
  not (_31235_, _31234_);
  or (_31256_, _31235_, _28477_);
  not (_31257_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31278_, \oc8051_top_1.oc8051_decoder1.wr , _18787_);
  not (_31279_, _31278_);
  nor (_31300_, _31279_, _27194_);
  and (_31301_, _31300_, _31257_);
  not (_31321_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_31322_, _28477_, _31321_);
  and (_31343_, _31322_, _31301_);
  and (_31344_, _31343_, _31256_);
  nor (_31365_, _31300_, _31321_);
  not (_31366_, _29858_);
  nor (_31387_, _30228_, _28565_);
  nor (_31388_, _31387_, _31366_);
  not (_31409_, _31388_);
  and (_31410_, _20908_, _30512_);
  nor (_31430_, _31410_, _29781_);
  nor (_31431_, _31430_, _28554_);
  and (_31452_, _29584_, _20071_);
  and (_31453_, _31452_, _30675_);
  nor (_31474_, _31453_, _30544_);
  nor (_31475_, _29584_, _20908_);
  not (_31496_, _31475_);
  nor (_31497_, _31496_, _30686_);
  nor (_31518_, _31497_, _30621_);
  and (_31519_, _31518_, _31474_);
  or (_31539_, _31519_, _30653_);
  nor (_31540_, _29573_, _29518_);
  not (_31561_, _29562_);
  and (_31562_, _30882_, _31561_);
  nor (_31583_, _31562_, _30850_);
  nor (_31584_, _31583_, _31540_);
  not (_31605_, _31584_);
  nor (_31606_, _30980_, _29584_);
  not (_31627_, _31606_);
  and (_31628_, _29540_, _29518_);
  and (_31648_, _30839_, _28542_);
  and (_31649_, _30915_, _29518_);
  nor (_31670_, _31649_, _31648_);
  nor (_31671_, _31670_, _31628_);
  not (_31692_, _31671_);
  and (_31693_, _31024_, _29573_);
  nor (_31714_, _30937_, _29573_);
  nor (_31715_, _31714_, _31693_);
  and (_31736_, _31715_, _31561_);
  nor (_31737_, _30795_, _22540_);
  and (_31757_, _30839_, _18809_);
  not (_31758_, _31757_);
  nor (_31769_, _31758_, _20908_);
  nor (_31780_, _31769_, _31737_);
  not (_31791_, _31780_);
  nor (_31802_, _31791_, _31736_);
  and (_31813_, _31802_, _31692_);
  and (_31824_, _31813_, _31627_);
  and (_31835_, _31824_, _31605_);
  not (_31846_, _31835_);
  nor (_31856_, _31846_, _31539_);
  not (_31867_, _31856_);
  nor (_31878_, _31867_, _31431_);
  and (_31889_, _31878_, _31409_);
  not (_31900_, _27369_);
  nor (_31911_, _27611_, _27490_);
  and (_31922_, _31911_, _31900_);
  and (_31933_, _31922_, _28466_);
  nand (_31944_, _31933_, _31889_);
  or (_31955_, _31933_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_31965_, _31300_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_31976_, _31965_, _31955_);
  and (_31987_, _31976_, _31944_);
  or (_31998_, _31987_, _31365_);
  or (_32009_, _31998_, _31344_);
  and (_06631_, _32009_, _42355_);
  and (_32030_, _26641_, _24210_);
  not (_32041_, _32030_);
  and (_32052_, _23935_, _18853_);
  and (_32063_, _29584_, _30010_);
  nor (_32073_, _32063_, _30021_);
  not (_32084_, _32073_);
  nor (_32095_, _29858_, _28543_);
  nor (_32106_, _32095_, _32084_);
  not (_32117_, _32106_);
  and (_32128_, _30882_, _29189_);
  not (_32139_, _32128_);
  and (_32150_, _30915_, _29168_);
  not (_32161_, _32150_);
  nor (_32172_, _30861_, _29178_);
  and (_32182_, _30937_, _22540_);
  nor (_32193_, _32182_, _32172_);
  and (_32204_, _32193_, _32161_);
  and (_32215_, _32204_, _32139_);
  nor (_32226_, _31758_, _29584_);
  not (_32237_, _32226_);
  nor (_32248_, _30566_, _19574_);
  and (_32259_, _30283_, _22540_);
  nor (_32270_, _32259_, _32248_);
  and (_32281_, _30272_, _29836_);
  not (_32291_, _32281_);
  nor (_32302_, _32291_, _21996_);
  not (_32313_, _32302_);
  and (_32324_, _31648_, _20919_);
  nor (_32335_, _30970_, _30610_);
  nor (_32346_, _32335_, _22540_);
  nor (_32357_, _32346_, _32324_);
  and (_32368_, _32357_, _32313_);
  and (_32379_, _32368_, _32270_);
  and (_32390_, _32379_, _32237_);
  and (_32400_, _32390_, _32215_);
  and (_32411_, _32400_, _32117_);
  not (_32422_, _32411_);
  nor (_32433_, _32422_, _32052_);
  and (_32444_, _32433_, _32041_);
  not (_32455_, _32444_);
  or (_32466_, _32455_, _28477_);
  not (_32477_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_32488_, _28477_, _32477_);
  and (_32499_, _32488_, _31301_);
  and (_32509_, _32499_, _32466_);
  nor (_32520_, _31300_, _32477_);
  not (_32531_, _31889_);
  or (_32542_, _32531_, _28477_);
  and (_32553_, _32488_, _31965_);
  and (_32564_, _32553_, _32542_);
  or (_32575_, _32564_, _32520_);
  or (_32586_, _32575_, _32509_);
  and (_08872_, _32586_, _42355_);
  and (_32607_, _26706_, _24210_);
  not (_32617_, _32607_);
  and (_32628_, _23966_, _18853_);
  nor (_32639_, _30566_, _20560_);
  nor (_32650_, _30392_, _30294_);
  not (_32661_, _32650_);
  nor (_32672_, _32661_, _29584_);
  and (_32683_, _32661_, _29584_);
  nor (_32694_, _32683_, _32672_);
  and (_32705_, _32694_, _30283_);
  nor (_32716_, _32705_, _32639_);
  nor (_32726_, _30642_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_32737_, _32726_, _22007_);
  nor (_32748_, _32726_, _22007_);
  nor (_32759_, _32748_, _32737_);
  nor (_32770_, _32759_, _30621_);
  not (_32781_, _32770_);
  and (_32792_, _30882_, _28981_);
  nor (_32803_, _30861_, _28970_);
  not (_32814_, _32803_);
  and (_32825_, _30915_, _28959_);
  and (_32836_, _30937_, _21996_);
  nor (_32846_, _32836_, _32825_);
  nand (_32857_, _32846_, _32814_);
  nor (_32868_, _32857_, _32792_);
  nor (_32879_, _31069_, _22540_);
  not (_32890_, _32879_);
  nor (_32901_, _30980_, _21996_);
  nor (_32912_, _32291_, _22171_);
  nor (_32923_, _32912_, _32901_);
  and (_32934_, _32923_, _32890_);
  and (_32944_, _32934_, _32868_);
  and (_32955_, _32944_, _32781_);
  and (_32966_, _32955_, _32716_);
  nor (_32977_, _29168_, _28981_);
  or (_32988_, _32977_, _29934_);
  and (_32999_, _32988_, _30021_);
  nor (_33010_, _32988_, _30021_);
  or (_33021_, _33010_, _32999_);
  and (_33032_, _33021_, _29858_);
  nor (_33043_, _29628_, _29595_);
  nor (_33053_, _33043_, _29639_);
  nor (_33064_, _33053_, _28554_);
  nor (_33075_, _33064_, _33032_);
  and (_33086_, _33075_, _32966_);
  not (_33097_, _33086_);
  nor (_33108_, _33097_, _32628_);
  and (_33119_, _33108_, _32617_);
  not (_33130_, _33119_);
  or (_33141_, _33130_, _28477_);
  not (_33152_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_33162_, _28477_, _33152_);
  and (_33173_, _33162_, _31301_);
  and (_33184_, _33173_, _33141_);
  nor (_33195_, _31300_, _33152_);
  not (_33206_, _27611_);
  and (_33217_, _33206_, _27490_);
  and (_33228_, _33217_, _27369_);
  and (_33239_, _33228_, _28466_);
  nand (_33250_, _33239_, _31889_);
  or (_33261_, _33239_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_33271_, _33261_, _31965_);
  and (_33282_, _33271_, _33250_);
  or (_33293_, _33282_, _33195_);
  or (_33304_, _33293_, _33184_);
  and (_08883_, _33304_, _42355_);
  and (_33325_, _26771_, _24210_);
  not (_33336_, _33325_);
  and (_33347_, _23998_, _18853_);
  nor (_33358_, _30566_, _19247_);
  and (_33369_, _30294_, _29584_);
  and (_33380_, _30392_, _30370_);
  nor (_33390_, _33380_, _33369_);
  and (_33401_, _33390_, _22171_);
  nor (_33412_, _33390_, _22171_);
  nor (_33423_, _33412_, _33401_);
  and (_33434_, _33423_, _30283_);
  nor (_33445_, _33434_, _33358_);
  nor (_33456_, _29639_, _29157_);
  nor (_33467_, _33456_, _29650_);
  nor (_33478_, _33467_, _28554_);
  not (_33489_, _33478_);
  nor (_33499_, _30054_, _30032_);
  nor (_33510_, _33499_, _31366_);
  and (_33521_, _33510_, _30076_);
  and (_33532_, _30632_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_33543_, _32748_, _22171_);
  nor (_33554_, _33543_, _33532_);
  nor (_33565_, _33554_, _30621_);
  and (_33576_, _30882_, _28948_);
  not (_33587_, _33576_);
  nor (_33598_, _30861_, _28937_);
  not (_33608_, _33598_);
  and (_33619_, _30915_, _28926_);
  and (_33630_, _30937_, _22171_);
  nor (_33641_, _33630_, _33619_);
  and (_33652_, _33641_, _33608_);
  and (_33663_, _33652_, _33587_);
  nor (_33674_, _30980_, _22171_);
  not (_33685_, _33674_);
  nor (_33696_, _32291_, _21670_);
  nor (_33706_, _31069_, _21996_);
  nor (_33717_, _33706_, _33696_);
  and (_33728_, _33717_, _33685_);
  and (_33739_, _33728_, _33663_);
  not (_33750_, _33739_);
  nor (_33761_, _33750_, _33565_);
  not (_33772_, _33761_);
  nor (_33783_, _33772_, _33521_);
  and (_33794_, _33783_, _33489_);
  and (_33805_, _33794_, _33445_);
  not (_33815_, _33805_);
  nor (_33826_, _33815_, _33347_);
  and (_33837_, _33826_, _33336_);
  not (_33848_, _33837_);
  or (_33859_, _33848_, _28477_);
  not (_33870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_33881_, _28477_, _33870_);
  and (_33892_, _33881_, _31301_);
  and (_33903_, _33892_, _33859_);
  nor (_33914_, _31300_, _33870_);
  nand (_33925_, _28466_, _27369_);
  or (_33935_, _31911_, _33925_);
  and (_33946_, _33935_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_33957_, _27490_);
  and (_33968_, _27369_, _27611_);
  and (_33979_, _33968_, _33957_);
  not (_33990_, _33979_);
  nor (_34001_, _33990_, _31889_);
  and (_34012_, _27369_, _27490_);
  and (_34023_, _34012_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_34034_, _34023_, _34001_);
  and (_34044_, _34034_, _28466_);
  or (_34055_, _34044_, _33946_);
  and (_34066_, _34055_, _31965_);
  or (_34077_, _34066_, _33914_);
  or (_34088_, _34077_, _33903_);
  and (_08894_, _34088_, _42355_);
  and (_34109_, _26836_, _24210_);
  and (_34120_, _24040_, _18853_);
  nand (_34131_, _30076_, _29999_);
  nor (_34142_, _31366_, _30087_);
  and (_34152_, _34142_, _34131_);
  nor (_34163_, _29650_, _29124_);
  or (_34174_, _34163_, _29661_);
  and (_34187_, _34174_, _28543_);
  nor (_34206_, _30566_, _20245_);
  and (_34217_, _30305_, _29584_);
  and (_34228_, _30403_, _30370_);
  nor (_34239_, _34228_, _34217_);
  nor (_34250_, _34239_, _21670_);
  not (_34261_, _30283_);
  and (_34271_, _34239_, _21670_);
  or (_34282_, _34271_, _34261_);
  nor (_34293_, _34282_, _34250_);
  nor (_34304_, _34293_, _34206_);
  not (_34315_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_34326_, _30632_, _34315_);
  or (_34337_, _34326_, _21681_);
  nor (_34348_, _30980_, _21670_);
  nor (_34359_, _30642_, _30621_);
  or (_34370_, _34359_, _34348_);
  and (_34380_, _34370_, _34337_);
  nor (_34391_, _30861_, _28882_);
  and (_34402_, _30882_, _28914_);
  nor (_34413_, _34402_, _34391_);
  and (_34424_, _30915_, _28893_);
  and (_34435_, _30937_, _21670_);
  nor (_34446_, _34435_, _34424_);
  nor (_34457_, _32291_, _21278_);
  nor (_34468_, _31069_, _22171_);
  nor (_34478_, _34468_, _34457_);
  and (_34489_, _34478_, _34446_);
  nand (_34500_, _34489_, _34413_);
  nor (_34511_, _34500_, _34380_);
  nand (_34522_, _34511_, _34304_);
  or (_34533_, _34522_, _34187_);
  or (_34544_, _34533_, _34152_);
  or (_34555_, _34544_, _34120_);
  or (_34566_, _34555_, _34109_);
  or (_34577_, _34566_, _28477_);
  not (_34588_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_34598_, _28477_, _34588_);
  and (_34609_, _34598_, _31301_);
  and (_34620_, _34609_, _34577_);
  nor (_34631_, _31300_, _34588_);
  and (_34642_, _33925_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_34653_, _31911_, _27369_);
  and (_34664_, _34653_, _32531_);
  or (_34675_, _31911_, _31900_);
  nor (_34686_, _34675_, _34588_);
  or (_34697_, _34686_, _34664_);
  and (_34707_, _34697_, _28466_);
  or (_34718_, _34707_, _34642_);
  and (_34729_, _34718_, _31965_);
  or (_34740_, _34729_, _34631_);
  or (_34751_, _34740_, _34620_);
  and (_08905_, _34751_, _42355_);
  and (_34772_, _26901_, _24210_);
  and (_34783_, _24072_, _18853_);
  nor (_34794_, _29727_, _28861_);
  and (_34805_, _29727_, _28861_);
  nor (_34815_, _34805_, _34794_);
  and (_34826_, _34815_, _28543_);
  or (_34837_, _30119_, _28861_);
  nor (_34848_, _31366_, _30130_);
  and (_34859_, _34848_, _34837_);
  nor (_34870_, _29584_, _19411_);
  and (_34881_, _29584_, _21289_);
  nor (_34892_, _34881_, _34870_);
  nor (_34903_, _34892_, _30566_);
  and (_34914_, _30316_, _29584_);
  and (_34924_, _30414_, _30370_);
  nor (_34935_, _34924_, _34914_);
  and (_34946_, _34935_, _21278_);
  nor (_34957_, _34935_, _21278_);
  nor (_34968_, _34957_, _34946_);
  and (_34979_, _34968_, _30283_);
  nor (_34990_, _34979_, _34903_);
  or (_35001_, _30653_, _21289_);
  nor (_35012_, _30664_, _30621_);
  and (_35023_, _35012_, _35001_);
  nor (_35033_, _30861_, _28850_);
  and (_35044_, _30882_, _28861_);
  nor (_35055_, _35044_, _35033_);
  and (_35066_, _30915_, _28839_);
  and (_35077_, _30937_, _21278_);
  nor (_35088_, _35077_, _35066_);
  nor (_35099_, _32291_, _21104_);
  nor (_35110_, _30980_, _21278_);
  nor (_35121_, _31069_, _21670_);
  or (_35132_, _35121_, _35110_);
  nor (_35142_, _35132_, _35099_);
  and (_35153_, _35142_, _35088_);
  nand (_35164_, _35153_, _35055_);
  nor (_35175_, _35164_, _35023_);
  nand (_35186_, _35175_, _34990_);
  or (_35197_, _35186_, _34859_);
  or (_35208_, _35197_, _34826_);
  or (_35218_, _35208_, _34783_);
  or (_35229_, _35218_, _34772_);
  or (_35240_, _35229_, _28477_);
  not (_35251_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_35262_, _28477_, _35251_);
  and (_35273_, _35262_, _31301_);
  and (_35284_, _35273_, _35240_);
  nor (_35295_, _31300_, _35251_);
  not (_35306_, _28466_);
  and (_35317_, _27622_, _31900_);
  nor (_35328_, _27622_, _31900_);
  nor (_35338_, _35328_, _35317_);
  or (_35349_, _35338_, _35306_);
  and (_35360_, _35349_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_35371_, _35317_, _32531_);
  and (_35382_, _35328_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_35393_, _35382_, _35371_);
  and (_35404_, _35393_, _28466_);
  or (_35415_, _35404_, _35360_);
  and (_35426_, _35415_, _31965_);
  or (_35437_, _35426_, _35295_);
  or (_35448_, _35437_, _35284_);
  and (_08916_, _35448_, _42355_);
  and (_35468_, _26987_, _24210_);
  not (_35479_, _35468_);
  and (_35490_, _24115_, _18853_);
  nor (_35501_, _30152_, _30130_);
  not (_35512_, _35501_);
  nor (_35523_, _31366_, _30163_);
  and (_35534_, _35523_, _35512_);
  not (_35545_, _35534_);
  nor (_35556_, _29738_, _28828_);
  nor (_35567_, _35556_, _29749_);
  nor (_35577_, _35567_, _28554_);
  nor (_35588_, _29584_, _20397_);
  and (_35599_, _29584_, _21125_);
  nor (_35610_, _35599_, _35588_);
  nor (_35621_, _35610_, _30566_);
  and (_35632_, _30336_, _29584_);
  and (_35643_, _30425_, _30370_);
  nor (_35654_, _35643_, _35632_);
  and (_35665_, _35654_, _21104_);
  nor (_35676_, _35654_, _21104_);
  or (_35687_, _35676_, _34261_);
  nor (_35698_, _35687_, _35665_);
  nor (_35708_, _35698_, _35621_);
  not (_35719_, _30719_);
  and (_35730_, _35719_, _30675_);
  nor (_35741_, _30719_, _30664_);
  nor (_35752_, _35741_, _21104_);
  nor (_35763_, _35752_, _35730_);
  nor (_35774_, _35763_, _30621_);
  nor (_35785_, _30861_, _28685_);
  and (_35796_, _30882_, _28696_);
  nor (_35807_, _35796_, _35785_);
  and (_35818_, _30915_, _28674_);
  and (_35828_, _30937_, _21104_);
  nor (_35839_, _35828_, _35818_);
  nor (_35850_, _30980_, _21104_);
  not (_35861_, _35850_);
  nor (_35872_, _32291_, _20071_);
  nor (_35883_, _31069_, _21278_);
  nor (_35894_, _35883_, _35872_);
  and (_35905_, _35894_, _35861_);
  and (_35916_, _35905_, _35839_);
  and (_35927_, _35916_, _35807_);
  not (_35938_, _35927_);
  nor (_35949_, _35938_, _35774_);
  and (_35959_, _35949_, _35708_);
  not (_35970_, _35959_);
  nor (_35981_, _35970_, _35577_);
  and (_35992_, _35981_, _35545_);
  not (_36003_, _35992_);
  nor (_36014_, _36003_, _35490_);
  and (_36025_, _36014_, _35479_);
  not (_36035_, _36025_);
  or (_36046_, _36035_, _28477_);
  not (_36057_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_36068_, _28477_, _36057_);
  and (_36079_, _36068_, _31301_);
  and (_36090_, _36079_, _36046_);
  nor (_36101_, _31300_, _36057_);
  and (_36112_, _33217_, _31900_);
  and (_36122_, _36112_, _28466_);
  nand (_36133_, _36122_, _31889_);
  or (_36144_, _36122_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_36155_, _36144_, _31965_);
  and (_36166_, _36155_, _36133_);
  or (_36177_, _36166_, _36101_);
  or (_36188_, _36177_, _36090_);
  and (_08927_, _36188_, _42355_);
  and (_36208_, _27052_, _24210_);
  not (_36219_, _36208_);
  and (_36230_, _24146_, _18853_);
  nor (_36241_, _30185_, _30163_);
  not (_36252_, _36241_);
  nor (_36263_, _31366_, _30196_);
  and (_36274_, _36263_, _36252_);
  not (_36284_, _36274_);
  nor (_36295_, _29749_, _28795_);
  nor (_36306_, _36295_, _29760_);
  nor (_36317_, _36306_, _28554_);
  nor (_36328_, _29584_, _28597_);
  or (_36339_, _36328_, _30566_);
  nor (_36350_, _36339_, _31452_);
  or (_36361_, _29584_, _21104_);
  or (_36371_, _35643_, _30337_);
  and (_36382_, _36371_, _36361_);
  nor (_36393_, _36382_, _20081_);
  not (_36404_, _36393_);
  and (_36415_, _36382_, _20081_);
  nor (_36426_, _36415_, _34261_);
  and (_36437_, _36426_, _36404_);
  nor (_36448_, _36437_, _36350_);
  nor (_36458_, _35730_, _20071_);
  and (_36469_, _35730_, _20071_);
  nor (_36480_, _36469_, _36458_);
  nor (_36491_, _36480_, _30621_);
  and (_36502_, _30882_, _28641_);
  nor (_36513_, _30861_, _28630_);
  not (_36524_, _36513_);
  and (_36534_, _30915_, _28619_);
  and (_36545_, _30937_, _20071_);
  nor (_36556_, _36545_, _36534_);
  nand (_36567_, _36556_, _36524_);
  nor (_36578_, _36567_, _36502_);
  nor (_36589_, _30980_, _20071_);
  not (_36600_, _36589_);
  nor (_36611_, _32291_, _20908_);
  nor (_36622_, _31069_, _21104_);
  nor (_36633_, _36622_, _36611_);
  and (_36643_, _36633_, _36600_);
  and (_36654_, _36643_, _36578_);
  not (_36665_, _36654_);
  nor (_36676_, _36665_, _36491_);
  and (_36687_, _36676_, _36448_);
  not (_36698_, _36687_);
  nor (_36709_, _36698_, _36317_);
  and (_36720_, _36709_, _36284_);
  not (_36731_, _36720_);
  nor (_36742_, _36731_, _36230_);
  and (_36752_, _36742_, _36219_);
  not (_36763_, _36752_);
  or (_36774_, _36763_, _28477_);
  not (_36785_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_36796_, _28477_, _36785_);
  and (_36807_, _36796_, _31301_);
  and (_36818_, _36807_, _36774_);
  nor (_36829_, _31300_, _36785_);
  nor (_36840_, _27369_, _27490_);
  and (_36851_, _36840_, _27611_);
  and (_36862_, _36851_, _28466_);
  nand (_36873_, _36862_, _31889_);
  or (_36884_, _36862_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_36895_, _36884_, _31965_);
  and (_36906_, _36895_, _36873_);
  or (_36917_, _36906_, _36829_);
  or (_36928_, _36917_, _36818_);
  and (_08938_, _36928_, _42355_);
  and (_36949_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_36960_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_36971_, _36960_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_36982_, _36971_);
  not (_36993_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_37003_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_37014_, _37003_, _36993_);
  and (_37025_, _36960_, _18787_);
  and (_37036_, _37025_, _37014_);
  not (_37047_, _37036_);
  not (_37058_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_37069_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_37080_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37091_, _37080_, _37069_);
  and (_37102_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_37112_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37123_, _37112_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_37134_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_37145_, _37134_, _37102_);
  and (_37156_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_37167_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37178_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _37167_);
  and (_37189_, _37178_, _37069_);
  and (_37200_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_37211_, _37200_, _37156_);
  and (_37222_, _37211_, _37145_);
  not (_37232_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_37243_, _37232_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_37254_, _37243_, _37069_);
  and (_37265_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_37276_, _37265_);
  and (_37287_, _37112_, _37069_);
  and (_37298_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_37309_, _37112_, _37069_);
  and (_37320_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_37331_, _37320_, _37298_);
  and (_37341_, _37331_, _37276_);
  and (_37352_, _37341_, _37222_);
  and (_37363_, _37352_, _37058_);
  nor (_37374_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _37058_);
  nor (_37385_, _37374_, _37363_);
  nor (_37396_, _37385_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_37407_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37418_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _37407_);
  nor (_37429_, _37418_, _37396_);
  nor (_37440_, _37429_, _37047_);
  not (_37451_, _37440_);
  not (_37462_, _37014_);
  nor (_37473_, _37025_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_37484_, _37473_, _37462_);
  and (_37495_, _37484_, _37451_);
  not (_37505_, _37495_);
  and (_37516_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_37527_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_37538_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_37542_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_37543_, _37542_, _37538_);
  and (_37544_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_37545_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_37546_, _37545_, _37544_);
  and (_37547_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_37548_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_37549_, _37548_, _37547_);
  and (_37550_, _37549_, _37546_);
  and (_37551_, _37550_, _37543_);
  nor (_37552_, _37551_, _37156_);
  and (_37553_, _37552_, _37058_);
  or (_37554_, _37553_, _37527_);
  and (_37555_, _37554_, _37407_);
  nor (_37556_, _37555_, _37516_);
  and (_37557_, _37556_, _37036_);
  not (_37558_, _37557_);
  nor (_37559_, _37025_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_37560_, _37559_, _37462_);
  and (_37561_, _37560_, _37558_);
  and (_37562_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37563_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37564_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_37565_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_37566_, _37565_, _37564_);
  and (_37567_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37568_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_37569_, _37568_, _37567_);
  and (_37570_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_37571_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_37572_, _37571_, _37570_);
  and (_37573_, _37572_, _37569_);
  and (_37574_, _37573_, _37566_);
  nor (_37575_, _37574_, _37156_);
  and (_37576_, _37575_, _37058_);
  or (_37577_, _37576_, _37563_);
  and (_37578_, _37577_, _37407_);
  nor (_37579_, _37578_, _37562_);
  and (_37580_, _37579_, _37036_);
  not (_37581_, _37580_);
  nor (_37582_, _37025_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_37583_, _37582_, _37462_);
  and (_37584_, _37583_, _37581_);
  not (_37585_, _37584_);
  and (_37586_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37587_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37588_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_37589_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_37590_, _37589_, _37588_);
  and (_37591_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_37592_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_37593_, _37592_, _37591_);
  and (_37594_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_37595_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_37596_, _37595_, _37594_);
  and (_37597_, _37596_, _37593_);
  and (_37598_, _37597_, _37590_);
  nor (_37599_, _37598_, _37156_);
  and (_37600_, _37599_, _37058_);
  or (_37601_, _37600_, _37587_);
  and (_37602_, _37601_, _37407_);
  nor (_37603_, _37602_, _37586_);
  nor (_37604_, _37603_, _37047_);
  and (_37605_, _37047_, \oc8051_top_1.oc8051_decoder1.op [6]);
  or (_37606_, _37605_, _37604_);
  and (_37607_, _37606_, _37014_);
  nor (_37608_, _37607_, _37585_);
  and (_37609_, _37608_, _37561_);
  and (_37610_, _37609_, _37505_);
  and (_37611_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37612_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37613_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_37614_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_37615_, _37614_, _37613_);
  and (_37616_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_37617_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_37618_, _37617_, _37616_);
  and (_37619_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_37620_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_37621_, _37620_, _37619_);
  and (_37622_, _37621_, _37618_);
  and (_37623_, _37622_, _37615_);
  nor (_37624_, _37623_, _37156_);
  and (_37625_, _37624_, _37058_);
  or (_37626_, _37625_, _37612_);
  and (_37627_, _37626_, _37407_);
  nor (_37628_, _37627_, _37611_);
  and (_37629_, _37628_, _37036_);
  not (_37630_, _37629_);
  nor (_37631_, _37025_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_37632_, _37631_, _37462_);
  and (_37633_, _37632_, _37630_);
  and (_37634_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_37635_, _37634_);
  and (_37636_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_37637_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_37638_, _37637_, _37636_);
  and (_37639_, _37638_, _37635_);
  and (_37640_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_37641_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_37642_, _37641_, _37640_);
  and (_37643_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_37644_, _37643_, _37156_);
  and (_37645_, _37644_, _37642_);
  and (_37646_, _37645_, _37639_);
  and (_37647_, _37646_, _37058_);
  nor (_37648_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _37058_);
  or (_37649_, _37648_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_37650_, _37649_, _37647_);
  and (_37651_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_37652_, _37651_, _37650_);
  nor (_37653_, _37652_, _37047_);
  not (_37654_, _37653_);
  nor (_37655_, _37025_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_37656_, _37655_, _37462_);
  and (_37657_, _37656_, _37654_);
  and (_37658_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37659_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37660_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_37661_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_37662_, _37661_, _37660_);
  and (_37663_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_37664_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_37665_, _37664_, _37663_);
  and (_37666_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_37667_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_37668_, _37667_, _37666_);
  and (_37669_, _37668_, _37665_);
  and (_37670_, _37669_, _37662_);
  nor (_37671_, _37670_, _37156_);
  and (_37672_, _37671_, _37058_);
  or (_37673_, _37672_, _37659_);
  and (_37674_, _37673_, _37407_);
  nor (_37675_, _37674_, _37658_);
  nor (_37676_, _37675_, _37047_);
  and (_37677_, _37047_, \oc8051_top_1.oc8051_decoder1.op [2]);
  or (_37678_, _37677_, _37676_);
  and (_37679_, _37678_, _37014_);
  and (_37680_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_37681_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_37682_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_37683_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_37684_, _37683_, _37682_);
  and (_37685_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_37686_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_37687_, _37686_, _37685_);
  and (_37688_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_37689_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_37690_, _37689_, _37688_);
  and (_37691_, _37690_, _37687_);
  and (_37692_, _37691_, _37684_);
  nor (_37693_, _37692_, _37156_);
  and (_37694_, _37693_, _37058_);
  or (_37695_, _37694_, _37681_);
  and (_37696_, _37695_, _37407_);
  nor (_37697_, _37696_, _37680_);
  and (_37698_, _37697_, _37036_);
  not (_37699_, _37698_);
  nor (_37700_, _37025_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_37701_, _37700_, _37462_);
  and (_37702_, _37701_, _37699_);
  nor (_37703_, _37702_, _37679_);
  and (_37704_, _37703_, _37657_);
  and (_37705_, _37704_, _37633_);
  and (_37706_, _37705_, _37610_);
  not (_37707_, _37706_);
  not (_37708_, _37561_);
  and (_37709_, _37607_, _37584_);
  and (_37710_, _37709_, _37708_);
  and (_37711_, _37710_, _37495_);
  and (_37712_, _37705_, _37711_);
  nor (_37713_, _37607_, _37584_);
  and (_37714_, _37713_, _37561_);
  and (_37715_, _37714_, _37495_);
  and (_37716_, _37705_, _37715_);
  nor (_37717_, _37716_, _37712_);
  and (_37718_, _37717_, _37707_);
  nor (_37719_, _37718_, _36982_);
  not (_37720_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_37721_, _18787_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_37722_, _37721_, _37720_);
  nor (_37723_, _37633_, _37657_);
  and (_37724_, _37723_, _37703_);
  and (_37725_, _37607_, _37708_);
  and (_37726_, _37725_, _37724_);
  and (_37727_, _37726_, _37722_);
  not (_37728_, _37727_);
  and (_37729_, _37714_, _37505_);
  not (_37730_, _37702_);
  and (_37731_, _37730_, _37679_);
  and (_37732_, _37723_, _37731_);
  and (_37733_, _37732_, _37729_);
  and (_37734_, _37732_, _37610_);
  nor (_37735_, _37734_, _37733_);
  and (_37736_, _37735_, _37728_);
  not (_37737_, _37736_);
  nor (_37738_, _37737_, _37719_);
  nor (_37739_, _37738_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37740_, _37739_, _36949_);
  and (_37741_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_37742_, _37657_);
  and (_37743_, _37633_, _37742_);
  and (_37744_, _37743_, _37731_);
  nor (_37745_, _37607_, _37561_);
  and (_37746_, _37745_, _37585_);
  and (_37747_, _37746_, _37495_);
  and (_37748_, _37747_, _37744_);
  not (_37749_, _37748_);
  not (_37750_, _37633_);
  and (_37751_, _37704_, _37750_);
  and (_37752_, _37609_, _37495_);
  and (_37753_, _37752_, _37751_);
  and (_37754_, _37607_, _37585_);
  and (_37755_, _37754_, _37561_);
  and (_37756_, _37755_, _37505_);
  and (_37757_, _37756_, _37751_);
  nor (_37758_, _37757_, _37753_);
  nand (_37759_, _37758_, _37749_);
  and (_37760_, _37724_, _37609_);
  and (_37761_, _37754_, _37708_);
  and (_37762_, _37761_, _37505_);
  and (_37763_, _37762_, _37744_);
  nor (_37764_, _37763_, _37760_);
  and (_37765_, _37755_, _37495_);
  and (_37766_, _37765_, _37744_);
  not (_37767_, _37766_);
  and (_37768_, _37711_, _37751_);
  and (_37769_, _37762_, _37704_);
  nor (_37770_, _37769_, _37768_);
  and (_37771_, _37770_, _37767_);
  nand (_37772_, _37771_, _37764_);
  nor (_37773_, _37772_, _37759_);
  and (_37774_, _37729_, _37751_);
  and (_37775_, _37761_, _37495_);
  and (_37776_, _37775_, _37704_);
  nor (_37777_, _37776_, _37774_);
  and (_37778_, _37715_, _37751_);
  and (_37779_, _37729_, _37744_);
  nor (_37780_, _37779_, _37778_);
  and (_37781_, _37780_, _37777_);
  and (_37782_, _37745_, _37584_);
  and (_37783_, _37782_, _37495_);
  and (_37784_, _37783_, _37724_);
  not (_37785_, _37784_);
  and (_37786_, _37782_, _37505_);
  and (_37787_, _37786_, _37724_);
  and (_37788_, _37724_, _37747_);
  nor (_37789_, _37788_, _37787_);
  and (_37790_, _37789_, _37785_);
  and (_37791_, _37724_, _37755_);
  and (_37792_, _37710_, _37505_);
  and (_37793_, _37792_, _37704_);
  nor (_37794_, _37793_, _37791_);
  and (_37795_, _37794_, _37790_);
  and (_37796_, _37795_, _37781_);
  and (_37797_, _37709_, _37561_);
  and (_37798_, _37797_, _37505_);
  and (_37799_, _37798_, _37744_);
  not (_37800_, _37799_);
  and (_37801_, _37657_, _37679_);
  and (_37802_, _37801_, _37730_);
  and (_37803_, _37802_, _37505_);
  and (_37804_, _37803_, _37609_);
  or (_37805_, _37715_, _37752_);
  and (_37806_, _37805_, _37744_);
  nor (_37807_, _37806_, _37804_);
  and (_37808_, _37807_, _37800_);
  not (_37809_, _37744_);
  nor (_37810_, _37782_, _37775_);
  nor (_37811_, _37810_, _37809_);
  not (_37812_, _37811_);
  and (_37813_, _37782_, _37751_);
  not (_37814_, _37813_);
  and (_37815_, _37746_, _37505_);
  and (_37816_, _37815_, _37744_);
  and (_37817_, _37610_, _37702_);
  nor (_37818_, _37817_, _37816_);
  and (_37819_, _37818_, _37814_);
  and (_37820_, _37819_, _37812_);
  and (_37821_, _37792_, _37744_);
  and (_37822_, _37756_, _37744_);
  nor (_37823_, _37822_, _37821_);
  and (_37824_, _37765_, _37751_);
  and (_37825_, _37610_, _37751_);
  nor (_37826_, _37825_, _37824_);
  and (_37827_, _37826_, _37823_);
  and (_37828_, _37827_, _37820_);
  and (_37829_, _37828_, _37808_);
  and (_37830_, _37829_, _37796_);
  and (_37831_, _37830_, _37773_);
  nor (_37832_, _37831_, _36982_);
  and (_37833_, \oc8051_top_1.oc8051_decoder1.state [0], _18787_);
  and (_37834_, _37833_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_37835_, _37834_, _37813_);
  nor (_37836_, _37835_, _37832_);
  and (_37837_, _37836_, _37728_);
  nor (_37838_, _37837_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37839_, _37838_, _37741_);
  and (_37840_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37841_, _37505_, _37702_);
  and (_37842_, _37841_, _37801_);
  and (_37843_, _37842_, _37761_);
  and (_37844_, _37802_, _37782_);
  or (_37845_, _37844_, _37843_);
  not (_37846_, _37845_);
  and (_37847_, _37802_, _37729_);
  nor (_37848_, _37847_, _37813_);
  and (_37849_, _37842_, _37609_);
  and (_37850_, _37802_, _37746_);
  or (_37851_, _37850_, _37849_);
  or (_37852_, _37797_, _37761_);
  and (_37853_, _37852_, _37803_);
  nor (_37854_, _37853_, _37851_);
  and (_37855_, _37854_, _37848_);
  and (_37856_, _37855_, _37846_);
  and (_37857_, _37765_, _37724_);
  not (_37858_, _37857_);
  and (_37859_, _37802_, _37755_);
  and (_37860_, _37842_, _37714_);
  nor (_37861_, _37860_, _37859_);
  not (_37862_, _37861_);
  and (_37863_, _37802_, _37792_);
  nor (_37864_, _37863_, _37862_);
  and (_37865_, _37864_, _37858_);
  and (_37866_, _37865_, _37718_);
  and (_37867_, _37866_, _37856_);
  nor (_37868_, _37867_, _36982_);
  and (_37869_, _37722_, _37724_);
  and (_37870_, _37869_, _37710_);
  or (_37871_, _37870_, _37835_);
  nor (_37872_, _37871_, _37868_);
  nor (_37873_, _37872_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_37874_, _37873_, _37840_);
  nor (_37875_, _37874_, _37839_);
  and (_37876_, _37875_, _37740_);
  and (_09488_, _37876_, _42355_);
  and (_37877_, _31301_, _28290_);
  and (_37878_, _37877_, _27369_);
  and (_37879_, _28433_, _27961_);
  not (_37880_, _27830_);
  nor (_37881_, _37880_, _28137_);
  and (_37882_, _37881_, _37879_);
  and (_37883_, _37882_, _33217_);
  and (_37884_, _37883_, _37878_);
  not (_37885_, _37884_);
  and (_37886_, _37885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_37887_, _24210_, _18853_);
  and (_37888_, _29847_, _24189_);
  nor (_37889_, _31047_, _37888_);
  and (_37890_, _37889_, _30980_);
  and (_37891_, _37890_, _37887_);
  and (_37892_, _37891_, _32291_);
  nor (_37893_, _37892_, _20071_);
  not (_37894_, _37893_);
  and (_37895_, _37894_, _36578_);
  and (_37896_, _37895_, _36448_);
  nor (_37897_, _37896_, _37885_);
  nor (_37898_, _37897_, _37886_);
  and (_37899_, _37885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_37900_, _37892_, _21104_);
  not (_37901_, _37900_);
  and (_37902_, _37901_, _35839_);
  and (_37903_, _37902_, _35807_);
  and (_37904_, _37903_, _35708_);
  nor (_37905_, _37904_, _37885_);
  nor (_37906_, _37905_, _37899_);
  and (_37907_, _37885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_37908_, _37892_, _21278_);
  not (_37909_, _37908_);
  and (_37910_, _37909_, _35088_);
  and (_37911_, _37910_, _35055_);
  and (_37912_, _37911_, _34990_);
  nor (_37913_, _37912_, _37885_);
  nor (_37914_, _37913_, _37907_);
  and (_37915_, _37885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_37916_, _37892_, _21670_);
  not (_37917_, _37916_);
  and (_37918_, _37917_, _34446_);
  and (_37919_, _37918_, _34413_);
  and (_37920_, _37919_, _34304_);
  nor (_37921_, _37920_, _37885_);
  nor (_37922_, _37921_, _37915_);
  and (_37923_, _37885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_37924_, _37892_, _22171_);
  not (_37925_, _37924_);
  and (_37926_, _37925_, _33663_);
  and (_37927_, _37926_, _33445_);
  nor (_37928_, _37927_, _37885_);
  nor (_37929_, _37928_, _37923_);
  and (_37930_, _37885_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_37931_, _37892_, _21996_);
  not (_37932_, _37931_);
  and (_37933_, _37932_, _32868_);
  and (_37934_, _37933_, _32716_);
  nor (_37935_, _37934_, _37885_);
  nor (_37936_, _37935_, _37930_);
  nor (_37937_, _37884_, _27556_);
  nor (_37938_, _37892_, _22540_);
  not (_37939_, _37938_);
  and (_37940_, _37939_, _32270_);
  and (_37941_, _37940_, _32215_);
  not (_37942_, _37941_);
  and (_37943_, _37942_, _37884_);
  nor (_37944_, _37943_, _37937_);
  and (_37945_, _37944_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_37946_, _37945_, _37936_);
  and (_37947_, _37946_, _37929_);
  and (_37948_, _37947_, _37922_);
  and (_37949_, _37948_, _37914_);
  and (_37950_, _37949_, _37906_);
  and (_37951_, _37950_, _37898_);
  nor (_37952_, _37884_, _27983_);
  nand (_37953_, _37952_, _37951_);
  or (_37954_, _37952_, _37951_);
  and (_37955_, _37954_, _27698_);
  and (_37956_, _37955_, _37953_);
  or (_37957_, _37884_, _28027_);
  or (_37958_, _37957_, _37956_);
  nor (_37959_, _37892_, _20908_);
  not (_37960_, _37959_);
  and (_37961_, _37960_, _30959_);
  and (_37962_, _37961_, _30904_);
  and (_37963_, _37962_, _30599_);
  nand (_37964_, _37963_, _37884_);
  and (_37965_, _37964_, _37958_);
  and (_09509_, _37965_, _42355_);
  not (_37966_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_37967_, _37944_, _37966_);
  nor (_37968_, _37944_, _37966_);
  nor (_37969_, _37968_, _37967_);
  and (_37970_, _37969_, _27698_);
  nor (_37971_, _37970_, _27567_);
  nor (_37972_, _37971_, _37884_);
  nor (_37973_, _37972_, _37943_);
  nand (_10665_, _37973_, _42355_);
  nor (_37974_, _37945_, _37936_);
  nor (_37975_, _37974_, _37946_);
  nor (_37976_, _37975_, _27106_);
  nor (_37977_, _37976_, _27402_);
  nor (_37978_, _37977_, _37884_);
  nor (_37979_, _37978_, _37935_);
  nand (_10676_, _37979_, _42355_);
  nor (_37980_, _37946_, _37929_);
  nor (_37981_, _37980_, _37947_);
  nor (_37982_, _37981_, _27106_);
  nor (_37983_, _37982_, _27161_);
  nor (_37984_, _37983_, _37884_);
  nor (_37985_, _37984_, _37928_);
  nand (_10687_, _37985_, _42355_);
  nor (_37986_, _37947_, _37922_);
  nor (_37987_, _37986_, _37948_);
  nor (_37988_, _37987_, _27106_);
  nor (_37989_, _37988_, _28225_);
  nor (_37990_, _37989_, _37884_);
  nor (_37991_, _37990_, _37921_);
  nor (_10698_, _37991_, rst);
  nor (_37992_, _37948_, _37914_);
  nor (_37993_, _37992_, _37949_);
  nor (_37994_, _37993_, _27106_);
  nor (_37995_, _37994_, _28356_);
  nor (_37996_, _37995_, _37884_);
  nor (_37997_, _37996_, _37913_);
  nor (_10709_, _37997_, rst);
  nor (_37998_, _37949_, _37906_);
  nor (_37999_, _37998_, _37950_);
  nor (_38000_, _37999_, _27106_);
  nor (_38001_, _38000_, _27884_);
  nor (_38002_, _38001_, _37884_);
  nor (_38003_, _38002_, _37905_);
  nor (_10720_, _38003_, rst);
  nor (_38004_, _37950_, _37898_);
  nor (_38005_, _38004_, _37951_);
  nor (_38006_, _38005_, _27106_);
  nor (_38007_, _38006_, _27731_);
  nor (_38008_, _38007_, _37884_);
  nor (_38009_, _38008_, _37897_);
  nor (_10731_, _38009_, rst);
  and (_38010_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18787_);
  and (_38011_, _38010_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_38012_, _38011_);
  nor (_38013_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_38014_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_38015_, _38014_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38016_, _38015_, _38013_);
  nor (_38017_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_38018_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_38019_, _38018_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38020_, _38019_, _38017_);
  not (_38021_, _38020_);
  nor (_38022_, _38021_, _31387_);
  nor (_38023_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_38024_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_38025_, _38024_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38026_, _38025_, _38023_);
  and (_38027_, _38026_, _38022_);
  nor (_38028_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_38029_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_38030_, _38029_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38031_, _38030_, _38028_);
  and (_38032_, _38031_, _38027_);
  and (_38033_, _38032_, _38016_);
  nor (_38034_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_38035_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_38036_, _38035_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38037_, _38036_, _38034_);
  and (_38038_, _38037_, _38033_);
  nor (_38039_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_38040_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_38041_, _38040_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38042_, _38041_, _38039_);
  and (_38043_, _38042_, _38038_);
  nor (_38044_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_38045_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_38046_, _38045_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38047_, _38046_, _38044_);
  and (_38048_, _38047_, _38043_);
  nor (_38049_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_38050_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_38051_, _38050_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_38052_, _38051_, _38049_);
  or (_38053_, _38052_, _38048_);
  nand (_38054_, _38052_, _38048_);
  and (_38055_, _38054_, _29858_);
  and (_38056_, _38055_, _38053_);
  not (_38057_, _38056_);
  and (_38058_, _23903_, _18853_);
  and (_38059_, _30348_, _20919_);
  and (_38060_, _38059_, _28992_);
  and (_38061_, _38060_, _29025_);
  and (_38062_, _38061_, _29069_);
  and (_38063_, _38062_, _29672_);
  and (_38064_, _38063_, _28707_);
  or (_38065_, _38064_, _30370_);
  and (_38066_, _30435_, _20908_);
  and (_38067_, _20245_, _19247_);
  and (_38068_, _20560_, _19574_);
  and (_38069_, _38068_, _38067_);
  and (_38070_, _38069_, _38066_);
  and (_38071_, _20397_, _19411_);
  and (_38072_, _38071_, _38070_);
  nor (_38073_, _38072_, _29584_);
  and (_38074_, _29584_, _20397_);
  nor (_38075_, _38074_, _38073_);
  and (_38076_, _38075_, _38065_);
  nor (_38077_, _29584_, _19748_);
  and (_38078_, _29584_, _19748_);
  nor (_38079_, _38078_, _38077_);
  and (_38080_, _38079_, _38076_);
  nor (_38081_, _38080_, _30512_);
  and (_38082_, _38080_, _30512_);
  nor (_38083_, _38082_, _38081_);
  and (_38084_, _38083_, _30283_);
  and (_38085_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_38086_, _29584_, _30512_);
  nor (_38087_, _38086_, _31475_);
  nor (_38088_, _38087_, _30566_);
  nor (_38089_, _31758_, _21670_);
  nor (_38090_, _30980_, _20734_);
  or (_38091_, _38090_, _38089_);
  or (_38092_, _38091_, _38088_);
  nor (_38093_, _38092_, _38085_);
  not (_38094_, _38093_);
  nor (_38095_, _38094_, _38084_);
  not (_38096_, _38095_);
  nor (_38097_, _38096_, _38058_);
  and (_38098_, _38097_, _38057_);
  nor (_38099_, _38098_, _38012_);
  and (_38100_, _37882_, _34653_);
  and (_38101_, _38100_, _37877_);
  or (_38102_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_38103_, _38102_, _38012_);
  nand (_38104_, _38101_, _31234_);
  and (_38105_, _38104_, _38103_);
  or (_38106_, _38105_, _38099_);
  and (_12682_, _38106_, _42355_);
  and (_38107_, _37882_, _33979_);
  and (_38108_, _38107_, _37877_);
  nor (_38109_, _38108_, _38011_);
  not (_38110_, _38109_);
  nand (_38111_, _38110_, _31234_);
  or (_38112_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_38113_, _38112_, _42355_);
  and (_12703_, _38113_, _38111_);
  and (_38114_, _26505_, _24210_);
  not (_38115_, _38114_);
  and (_38116_, _38021_, _31387_);
  nor (_38117_, _38116_, _38022_);
  and (_38118_, _38117_, _29858_);
  nor (_38119_, _31475_, _30544_);
  not (_38120_, _38119_);
  nor (_38121_, _38120_, _30457_);
  nor (_38122_, _38121_, _28992_);
  and (_38123_, _38121_, _28992_);
  nor (_38124_, _38123_, _38122_);
  and (_38125_, _38124_, _30283_);
  nor (_38126_, _30980_, _19574_);
  and (_38127_, _23682_, _18853_);
  nor (_38128_, _31758_, _21278_);
  nor (_38129_, _30566_, _22540_);
  or (_38130_, _38129_, _38128_);
  or (_38131_, _38130_, _38127_);
  nor (_38132_, _38131_, _38126_);
  not (_38133_, _38132_);
  nor (_38134_, _38133_, _38125_);
  not (_38135_, _38134_);
  nor (_38136_, _38135_, _38118_);
  and (_38137_, _38136_, _38115_);
  nor (_38138_, _38137_, _38012_);
  or (_38139_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_38140_, _38139_, _38012_);
  nand (_38141_, _38101_, _32444_);
  and (_38142_, _38141_, _38140_);
  or (_38143_, _38142_, _38138_);
  and (_13618_, _38143_, _42355_);
  nor (_38144_, _38026_, _38022_);
  nor (_38145_, _38144_, _38027_);
  and (_38146_, _38145_, _29858_);
  not (_38147_, _38146_);
  and (_38148_, _25519_, _24210_);
  nor (_38149_, _38060_, _30370_);
  and (_38150_, _38066_, _19574_);
  nor (_38151_, _38150_, _29584_);
  or (_38152_, _38151_, _38149_);
  and (_38153_, _38152_, _20560_);
  nor (_38154_, _38152_, _20560_);
  or (_38155_, _38154_, _34261_);
  nor (_38156_, _38155_, _38153_);
  nor (_38157_, _30980_, _20560_);
  and (_38158_, _23713_, _18853_);
  nor (_38159_, _31758_, _21104_);
  nor (_38160_, _30566_, _21996_);
  or (_38161_, _38160_, _38159_);
  or (_38162_, _38161_, _38158_);
  nor (_38163_, _38162_, _38157_);
  not (_38164_, _38163_);
  nor (_38165_, _38164_, _38156_);
  not (_38166_, _38165_);
  nor (_38167_, _38166_, _38148_);
  and (_38168_, _38167_, _38147_);
  nor (_38169_, _38168_, _38012_);
  or (_38170_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_38171_, _38170_, _38012_);
  nand (_38172_, _38101_, _33119_);
  and (_38173_, _38172_, _38171_);
  or (_38174_, _38173_, _38169_);
  and (_13629_, _38174_, _42355_);
  nor (_38175_, _38031_, _38027_);
  nor (_38176_, _38175_, _38032_);
  and (_38177_, _38176_, _29858_);
  not (_38178_, _38177_);
  and (_38179_, _38150_, _20560_);
  and (_38180_, _38179_, _30370_);
  and (_38181_, _38061_, _29584_);
  nor (_38182_, _38181_, _38180_);
  and (_38183_, _38182_, _19247_);
  nor (_38184_, _38182_, _19247_);
  nor (_38185_, _38184_, _38183_);
  and (_38186_, _38185_, _30283_);
  not (_38187_, _38186_);
  nor (_38188_, _30566_, _22171_);
  and (_38189_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_38190_, _38189_, _38188_);
  and (_38191_, _23745_, _18853_);
  nor (_38192_, _31758_, _20071_);
  nor (_38193_, _30980_, _19247_);
  or (_38194_, _38193_, _38192_);
  nor (_38195_, _38194_, _38191_);
  and (_38196_, _38195_, _38190_);
  and (_38197_, _38196_, _38187_);
  and (_38198_, _38197_, _38178_);
  nor (_38199_, _38198_, _38012_);
  or (_38200_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_38201_, _38200_, _38012_);
  nand (_38202_, _38101_, _33837_);
  and (_38203_, _38202_, _38201_);
  or (_38204_, _38203_, _38199_);
  and (_13640_, _38204_, _42355_);
  or (_38205_, _38032_, _38016_);
  nor (_38206_, _38033_, _31366_);
  and (_38207_, _38206_, _38205_);
  and (_38208_, _23777_, _18853_);
  nor (_38209_, _38063_, _30370_);
  or (_38210_, _38062_, _29672_);
  and (_38211_, _38210_, _38209_);
  nand (_38212_, _38179_, _19247_);
  and (_38213_, _38212_, _29672_);
  or (_38214_, _38213_, _38070_);
  and (_38215_, _38214_, _30370_);
  or (_38216_, _38215_, _38211_);
  and (_38217_, _38216_, _30283_);
  nor (_38218_, _30566_, _21670_);
  nor (_38219_, _30980_, _20245_);
  and (_38220_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_38221_, _38220_, _38219_);
  or (_38222_, _38221_, _31769_);
  or (_38223_, _38222_, _38218_);
  or (_38224_, _38223_, _38217_);
  or (_38225_, _38224_, _38208_);
  or (_38226_, _38225_, _38207_);
  and (_38227_, _38226_, _38011_);
  or (_38228_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_38229_, _38228_, _38012_);
  not (_38230_, _38101_);
  or (_38231_, _38230_, _34566_);
  and (_38232_, _38231_, _38229_);
  or (_38233_, _38232_, _38227_);
  and (_13651_, _38233_, _42355_);
  or (_38234_, _38037_, _38033_);
  nor (_38235_, _38038_, _31366_);
  and (_38236_, _38235_, _38234_);
  and (_38237_, _23818_, _18853_);
  nor (_38238_, _38070_, _29584_);
  nor (_38239_, _38238_, _38209_);
  or (_38240_, _38239_, _28707_);
  nand (_38241_, _38239_, _28707_);
  and (_38242_, _38241_, _38240_);
  and (_38243_, _38242_, _30283_);
  or (_38244_, _29584_, _21289_);
  nand (_38245_, _29584_, _19411_);
  and (_38246_, _38245_, _30555_);
  and (_38247_, _38246_, _38244_);
  nor (_38248_, _31758_, _22540_);
  nor (_38249_, _30980_, _19411_);
  and (_38250_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_38251_, _38250_, _38249_);
  or (_38252_, _38251_, _38248_);
  or (_38253_, _38252_, _38247_);
  or (_38254_, _38253_, _38243_);
  or (_38255_, _38254_, _38237_);
  or (_38256_, _38255_, _38236_);
  and (_38257_, _38256_, _38011_);
  or (_38258_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_38259_, _38258_, _38012_);
  or (_38260_, _38230_, _35229_);
  and (_38261_, _38260_, _38259_);
  or (_38262_, _38261_, _38257_);
  and (_13662_, _38262_, _42355_);
  nor (_38263_, _38042_, _38038_);
  not (_38264_, _38263_);
  nor (_38265_, _38043_, _31366_);
  and (_38266_, _38265_, _38264_);
  not (_38267_, _38266_);
  and (_38268_, _23840_, _18853_);
  and (_38269_, _38070_, _19411_);
  nor (_38270_, _38269_, _29584_);
  not (_38271_, _38270_);
  and (_38272_, _38271_, _38065_);
  and (_38273_, _38272_, _20397_);
  nor (_38274_, _38272_, _20397_);
  nor (_38275_, _38274_, _38273_);
  nor (_38276_, _38275_, _34261_);
  nor (_38277_, _29584_, _21125_);
  or (_38278_, _38277_, _30566_);
  nor (_38279_, _38278_, _38074_);
  nor (_38280_, _30980_, _20397_);
  nor (_38281_, _31758_, _21996_);
  and (_38282_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_38283_, _38282_, _38281_);
  nor (_38284_, _38283_, _38280_);
  not (_38285_, _38284_);
  nor (_38286_, _38285_, _38279_);
  not (_38287_, _38286_);
  nor (_38288_, _38287_, _38276_);
  not (_38289_, _38288_);
  nor (_38290_, _38289_, _38268_);
  and (_38291_, _38290_, _38267_);
  nor (_38292_, _38291_, _38012_);
  or (_38293_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_38294_, _38293_, _38012_);
  nand (_38295_, _38101_, _36025_);
  and (_38296_, _38295_, _38294_);
  or (_38297_, _38296_, _38292_);
  and (_13672_, _38297_, _42355_);
  nor (_38298_, _38047_, _38043_);
  nor (_38299_, _38298_, _38048_);
  and (_38300_, _38299_, _29858_);
  and (_38301_, _23871_, _18853_);
  and (_38302_, _38076_, _19748_);
  nor (_38303_, _38076_, _19748_);
  or (_38304_, _38303_, _38302_);
  and (_38305_, _38304_, _30283_);
  or (_38306_, _29584_, _20081_);
  nor (_38307_, _38078_, _30566_);
  and (_38308_, _38307_, _38306_);
  nor (_38309_, _31758_, _22171_);
  nor (_38310_, _30980_, _19748_);
  and (_38311_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or (_38312_, _38311_, _38310_);
  or (_38313_, _38312_, _38309_);
  or (_38314_, _38313_, _38308_);
  or (_38315_, _38314_, _38305_);
  or (_38316_, _38315_, _38301_);
  or (_38317_, _38316_, _38300_);
  and (_38318_, _38317_, _38011_);
  or (_38319_, _38101_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_38320_, _38319_, _38012_);
  nand (_38321_, _38101_, _36752_);
  and (_38322_, _38321_, _38320_);
  or (_38323_, _38322_, _38318_);
  and (_13683_, _38323_, _42355_);
  nand (_38324_, _38110_, _32444_);
  or (_38325_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_38326_, _38325_, _42355_);
  and (_13694_, _38326_, _38324_);
  nand (_38327_, _38110_, _33119_);
  or (_38328_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_38329_, _38328_, _42355_);
  and (_13705_, _38329_, _38327_);
  nand (_38330_, _38110_, _33837_);
  or (_38331_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_38332_, _38331_, _42355_);
  and (_13716_, _38332_, _38330_);
  or (_38333_, _38109_, _34566_);
  or (_38334_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_38335_, _38334_, _42355_);
  and (_13727_, _38335_, _38333_);
  or (_38336_, _38109_, _35229_);
  or (_38337_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_38338_, _38337_, _42355_);
  and (_13738_, _38338_, _38336_);
  nand (_38339_, _38110_, _36025_);
  or (_38340_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_38341_, _38340_, _42355_);
  and (_13749_, _38341_, _38339_);
  nand (_38342_, _38110_, _36752_);
  or (_38343_, _38110_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_38344_, _38343_, _42355_);
  and (_13760_, _38344_, _38342_);
  not (_38345_, _27961_);
  nor (_38346_, _38345_, _27830_);
  and (_38347_, _38346_, _31965_);
  and (_38348_, _38347_, _28455_);
  not (_38349_, _31922_);
  nor (_38350_, _38349_, _31889_);
  not (_38351_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_38352_, _31922_, _38351_);
  or (_38353_, _38352_, _38350_);
  and (_38354_, _38353_, _38348_);
  nor (_38355_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_38356_, _38355_);
  nand (_38357_, _38356_, _31889_);
  and (_38358_, _38355_, _38351_);
  nor (_38359_, _38358_, _38348_);
  and (_38360_, _38359_, _38357_);
  nor (_38361_, _28433_, _38345_);
  nor (_38362_, _27830_, _28137_);
  and (_38363_, _37877_, _27633_);
  and (_38364_, _38363_, _38362_);
  and (_38365_, _38364_, _38361_);
  or (_38366_, _38365_, _38360_);
  or (_38367_, _38366_, _38354_);
  nand (_38368_, _38365_, _37963_);
  and (_38369_, _38368_, _42355_);
  and (_15163_, _38369_, _38367_);
  and (_38370_, _38361_, _38362_);
  and (_38371_, _38370_, _38363_);
  and (_38372_, _38348_, _33228_);
  nand (_38373_, _38372_, _31889_);
  or (_38374_, _38372_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_38375_, _38374_, _38373_);
  or (_38376_, _38375_, _38371_);
  nand (_38377_, _38365_, _37934_);
  and (_38378_, _38377_, _42355_);
  and (_17344_, _38378_, _38376_);
  and (_38379_, _31410_, _29771_);
  not (_38380_, _29771_);
  and (_38383_, _31430_, _38380_);
  or (_38385_, _38383_, _38379_);
  and (_38386_, _38385_, _28543_);
  not (_38387_, _28565_);
  nand (_38388_, _30217_, _38387_);
  or (_38389_, _30217_, _28575_);
  and (_38390_, _29858_, _38389_);
  and (_38391_, _38390_, _38388_);
  and (_38392_, _38071_, _25420_);
  and (_38393_, _38069_, _24210_);
  nand (_38394_, _38393_, _38392_);
  nand (_38396_, _38394_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_38405_, _38396_, _38391_);
  or (_38411_, _38405_, _38386_);
  or (_38417_, _23966_, _23935_);
  or (_38420_, _38417_, _23998_);
  or (_38421_, _38420_, _24040_);
  or (_38422_, _38421_, _24072_);
  or (_38423_, _38422_, _24115_);
  or (_38424_, _38423_, _24146_);
  and (_38425_, _38424_, _18853_);
  or (_38426_, _38425_, _38411_);
  or (_38427_, _38426_, _28510_);
  nor (_38428_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_38429_, _38428_, _38348_);
  and (_38430_, _38429_, _38427_);
  and (_38431_, _33990_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_38432_, _38431_, _34001_);
  and (_38433_, _38432_, _38348_);
  or (_38434_, _38433_, _38365_);
  or (_38435_, _38434_, _38430_);
  nand (_38436_, _38365_, _37927_);
  and (_38437_, _38436_, _42355_);
  and (_17355_, _38437_, _38435_);
  and (_38438_, _38348_, _34653_);
  nand (_38439_, _38438_, _31889_);
  not (_38440_, _38365_);
  or (_38441_, _38438_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_38442_, _38441_, _38440_);
  and (_38443_, _38442_, _38439_);
  nor (_38446_, _38440_, _37920_);
  or (_38447_, _38446_, _38443_);
  and (_17366_, _38447_, _42355_);
  not (_38448_, _38348_);
  or (_38449_, _38448_, _35338_);
  not (_38450_, _38371_);
  and (_38451_, _38450_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_38452_, _38450_, _37912_);
  nor (_38453_, _38452_, _38451_);
  nor (_38482_, _38453_, rst);
  and (_38454_, _38482_, _38449_);
  and (_38455_, _35328_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_38456_, _38455_, _35371_);
  and (_38457_, _38348_, _42355_);
  and (_38458_, _38457_, _38456_);
  or (_17377_, _38458_, _38454_);
  and (_38459_, _38348_, _36112_);
  nand (_38460_, _38459_, _31889_);
  or (_38461_, _38459_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_38462_, _38461_, _38440_);
  and (_38463_, _38462_, _38460_);
  nor (_38464_, _38440_, _37904_);
  or (_38465_, _38464_, _38463_);
  and (_17388_, _38465_, _42355_);
  not (_38466_, _36851_);
  nor (_38467_, _38466_, _31889_);
  or (_38468_, _36851_, _34315_);
  nand (_38469_, _38468_, _38348_);
  or (_38470_, _38469_, _38467_);
  and (_38471_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_38472_, _29858_, _30119_);
  and (_38473_, _29727_, _28543_);
  or (_38474_, _38473_, _38472_);
  and (_38475_, _38474_, _38471_);
  nand (_38476_, _38471_, _30980_);
  and (_38477_, _38476_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_38478_, _38477_, _38348_);
  or (_38479_, _38478_, _38475_);
  and (_38481_, _38479_, _38440_);
  nor (_38485_, _38440_, _37896_);
  or (_38491_, _38485_, _38481_);
  and (_38496_, _38491_, _42355_);
  and (_17399_, _38496_, _38470_);
  not (_38510_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38518_, _38010_, _38510_);
  and (_38519_, _38518_, _38098_);
  nor (_38520_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_38521_, _38520_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_38522_, _27633_, _28290_);
  and (_38523_, _28433_, _38345_);
  and (_38524_, _38523_, _38362_);
  and (_38525_, _38524_, _38522_);
  and (_38526_, _38525_, _31301_);
  nor (_38527_, _38526_, _38521_);
  nor (_38528_, _38527_, _31234_);
  and (_38529_, _28433_, _28290_);
  and (_38530_, _38529_, _27972_);
  not (_38531_, _31965_);
  nor (_38532_, _38531_, _28137_);
  and (_38533_, _38532_, _38530_);
  and (_38534_, _38533_, _31922_);
  and (_38535_, _38534_, _31889_);
  nor (_38536_, _38534_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_38537_, _38521_, _38518_);
  not (_38538_, _38537_);
  nor (_38539_, _38538_, _38526_);
  not (_38540_, _38539_);
  nor (_38541_, _38540_, _38536_);
  not (_38542_, _38541_);
  nor (_38543_, _38542_, _38535_);
  nor (_38544_, _38543_, _38518_);
  not (_38545_, _38544_);
  nor (_38546_, _38545_, _38528_);
  nor (_38547_, _38546_, _38519_);
  and (_17968_, _38547_, _42355_);
  not (_38548_, _38518_);
  nor (_38549_, _38548_, _38137_);
  not (_38550_, _38527_);
  and (_38551_, _38550_, _32444_);
  not (_38552_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_38553_, _38533_, _38552_);
  not (_38554_, _38553_);
  and (_38560_, _32531_, _27633_);
  nor (_38571_, _27633_, _38552_);
  nor (_38572_, _38571_, _38560_);
  nand (_38573_, _38539_, _38533_);
  or (_38574_, _38573_, _38572_);
  and (_38585_, _38574_, _38527_);
  and (_38591_, _38585_, _38554_);
  nor (_38592_, _38591_, _38518_);
  not (_38593_, _38592_);
  nor (_38594_, _38593_, _38551_);
  nor (_38595_, _38594_, _38549_);
  nor (_19759_, _38595_, rst);
  nor (_38596_, _38527_, _33119_);
  and (_38597_, _38533_, _33228_);
  and (_38598_, _38597_, _31889_);
  nor (_38599_, _38597_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_38600_, _38599_, _38540_);
  not (_38601_, _38600_);
  nor (_38602_, _38601_, _38598_);
  or (_38603_, _38602_, _38596_);
  and (_38604_, _38603_, _38548_);
  nor (_38605_, _38548_, _38168_);
  or (_38606_, _38605_, _38604_);
  and (_19771_, _38606_, _42355_);
  and (_38607_, _38518_, _38198_);
  nor (_38608_, _38527_, _33837_);
  and (_38609_, _38533_, _33979_);
  nor (_38610_, _38609_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_38611_, _38610_);
  and (_38612_, _38609_, _31889_);
  nor (_38613_, _38612_, _38540_);
  and (_38614_, _38613_, _38611_);
  nor (_38615_, _38614_, _38518_);
  not (_38616_, _38615_);
  nor (_38617_, _38616_, _38608_);
  nor (_38618_, _38617_, _38607_);
  and (_19783_, _38618_, _42355_);
  and (_38619_, _38518_, _38226_);
  or (_38620_, _38527_, _34566_);
  not (_38621_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_38622_, _38533_, _38621_);
  nor (_38623_, _34653_, _38621_);
  or (_38624_, _38623_, _34664_);
  and (_38625_, _38624_, _38533_);
  or (_38626_, _38625_, _38550_);
  or (_38627_, _38626_, _38622_);
  and (_38628_, _38627_, _38548_);
  and (_38629_, _38628_, _38620_);
  or (_38630_, _38629_, _38619_);
  and (_19795_, _38630_, _42355_);
  or (_38631_, _38548_, _38256_);
  and (_38632_, _38550_, _35229_);
  and (_38633_, _38533_, _35317_);
  or (_38634_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_38635_, _38633_, _31889_);
  and (_38636_, _38635_, _38539_);
  and (_38637_, _38636_, _38634_);
  or (_38638_, _38637_, _38518_);
  or (_38639_, _38638_, _38632_);
  and (_38640_, _38639_, _38631_);
  and (_19807_, _38640_, _42355_);
  and (_38641_, _38518_, _38291_);
  nor (_38642_, _38527_, _36025_);
  and (_38643_, _38533_, _36112_);
  and (_38644_, _38643_, _31889_);
  nor (_38645_, _38643_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_38646_, _38645_, _38540_);
  not (_38647_, _38646_);
  nor (_38648_, _38647_, _38644_);
  nor (_38649_, _38648_, _38518_);
  not (_38650_, _38649_);
  nor (_38651_, _38650_, _38642_);
  nor (_38652_, _38651_, _38641_);
  and (_19819_, _38652_, _42355_);
  and (_38653_, _38518_, _38317_);
  and (_38654_, _38550_, _36752_);
  not (_38655_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_38656_, _38533_, _38655_);
  nor (_38657_, _38656_, _38550_);
  not (_38658_, _38657_);
  not (_38659_, _38533_);
  nor (_38660_, _36851_, _38655_);
  nor (_38661_, _38660_, _38467_);
  nor (_38662_, _38661_, _38659_);
  nor (_38663_, _38662_, _38658_);
  nor (_38664_, _38663_, _38518_);
  not (_38665_, _38664_);
  nor (_38666_, _38665_, _38654_);
  nor (_38667_, _38666_, _38653_);
  nor (_19831_, _38667_, rst);
  and (_38668_, _27961_, _27830_);
  and (_38669_, _38529_, _28148_);
  and (_38670_, _38669_, _38668_);
  and (_38671_, _38670_, _31922_);
  nand (_38672_, _38671_, _31889_);
  or (_38673_, _38671_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38674_, _38673_, _31965_);
  and (_38675_, _38674_, _38672_);
  and (_38676_, _37882_, _38522_);
  nand (_38677_, _38676_, _37963_);
  or (_38678_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_38679_, _38678_, _31301_);
  and (_38680_, _38679_, _38677_);
  not (_38681_, _31300_);
  and (_38682_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_38683_, _38682_, rst);
  or (_38684_, _38683_, _38680_);
  or (_31035_, _38684_, _38675_);
  and (_38685_, _38668_, _28455_);
  and (_38686_, _38685_, _31922_);
  nand (_38687_, _38686_, _31889_);
  or (_38688_, _38686_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_38689_, _38688_, _31965_);
  and (_38690_, _38689_, _38687_);
  and (_38691_, _38361_, _37881_);
  and (_38692_, _38691_, _38522_);
  nand (_38693_, _38692_, _37963_);
  or (_38694_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_38695_, _38694_, _31301_);
  and (_38696_, _38695_, _38693_);
  and (_38697_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_38698_, _38697_, rst);
  or (_38699_, _38698_, _38696_);
  or (_31058_, _38699_, _38690_);
  and (_38700_, _38345_, _27830_);
  and (_38701_, _38700_, _38669_);
  and (_38702_, _38701_, _31922_);
  nand (_38703_, _38702_, _31889_);
  or (_38704_, _38702_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_38705_, _38704_, _31965_);
  and (_38706_, _38705_, _38703_);
  and (_38707_, _38523_, _37881_);
  and (_38708_, _38707_, _38522_);
  not (_38709_, _38708_);
  nor (_38710_, _38709_, _37963_);
  and (_38711_, _38709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_38712_, _38711_, _38710_);
  and (_38713_, _38712_, _31301_);
  and (_38714_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_38715_, _38714_, rst);
  or (_38716_, _38715_, _38713_);
  or (_31081_, _38716_, _38706_);
  and (_38717_, _38700_, _28455_);
  and (_38718_, _38717_, _31922_);
  nand (_38719_, _38718_, _31889_);
  or (_38720_, _38718_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_38721_, _38720_, _31965_);
  and (_38722_, _38721_, _38719_);
  nor (_38723_, _28433_, _27961_);
  and (_38724_, _37881_, _38723_);
  and (_38725_, _38724_, _38522_);
  not (_38726_, _38725_);
  nor (_38727_, _38726_, _37963_);
  and (_38728_, _38726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_38729_, _38728_, _38727_);
  and (_38730_, _38729_, _31301_);
  and (_38731_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_38732_, _38731_, rst);
  or (_38733_, _38732_, _38730_);
  or (_31103_, _38733_, _38722_);
  or (_38734_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_38735_, _38734_, _31965_);
  and (_38736_, _38670_, _27633_);
  nand (_38737_, _38736_, _31889_);
  and (_38738_, _38737_, _38735_);
  nand (_38739_, _38676_, _37941_);
  and (_38740_, _38739_, _31301_);
  and (_38741_, _38740_, _38734_);
  not (_38742_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_38743_, _31300_, _38742_);
  or (_38744_, _38743_, rst);
  or (_38745_, _38744_, _38741_);
  or (_40047_, _38745_, _38738_);
  and (_38746_, _33228_, _28290_);
  and (_38747_, _38746_, _37882_);
  nand (_38748_, _38747_, _31889_);
  or (_38749_, _38747_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_38750_, _38749_, _31965_);
  and (_38751_, _38750_, _38748_);
  nand (_38752_, _38676_, _37934_);
  or (_38753_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_38754_, _38753_, _31301_);
  and (_38755_, _38754_, _38752_);
  and (_38756_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_38757_, _38756_, rst);
  or (_38758_, _38757_, _38755_);
  or (_40048_, _38758_, _38751_);
  not (_38759_, _34675_);
  nand (_38760_, _38670_, _38759_);
  and (_38761_, _38760_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_38762_, _34012_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_38763_, _38762_, _34001_);
  and (_38764_, _38763_, _38670_);
  or (_38765_, _38764_, _38761_);
  and (_38774_, _38765_, _31965_);
  nand (_38785_, _38676_, _37927_);
  or (_38796_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_38805_, _38796_, _31301_);
  and (_38811_, _38805_, _38785_);
  and (_38822_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_38833_, _38822_, rst);
  or (_38844_, _38833_, _38811_);
  or (_40050_, _38844_, _38774_);
  nand (_38865_, _38670_, _27369_);
  and (_38876_, _38865_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_38887_, _38759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_38898_, _38887_, _34664_);
  and (_38909_, _38898_, _38670_);
  or (_38920_, _38909_, _38876_);
  and (_38931_, _38920_, _31965_);
  nand (_38942_, _38676_, _37920_);
  or (_38953_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_38964_, _38953_, _31301_);
  and (_38975_, _38964_, _38942_);
  and (_38979_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_38980_, _38979_, rst);
  or (_38981_, _38980_, _38975_);
  or (_40052_, _38981_, _38931_);
  not (_38982_, _38670_);
  or (_38983_, _38982_, _35338_);
  and (_38984_, _38983_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_38985_, _35328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_38986_, _38985_, _35371_);
  and (_38987_, _38986_, _38670_);
  or (_38988_, _38987_, _38984_);
  and (_38989_, _38988_, _31965_);
  nand (_38990_, _38676_, _37912_);
  or (_38991_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_38992_, _38991_, _31301_);
  and (_38993_, _38992_, _38990_);
  and (_38994_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_38995_, _38994_, rst);
  or (_38996_, _38995_, _38993_);
  or (_40054_, _38996_, _38989_);
  and (_38997_, _38670_, _36112_);
  nand (_38998_, _38997_, _31889_);
  or (_38999_, _38997_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39000_, _38999_, _31965_);
  and (_39001_, _39000_, _38998_);
  nand (_39002_, _38676_, _37904_);
  or (_39003_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_39004_, _39003_, _31301_);
  and (_39005_, _39004_, _39002_);
  and (_39006_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_39007_, _39006_, rst);
  or (_39008_, _39007_, _39005_);
  or (_40056_, _39008_, _39001_);
  and (_39009_, _38670_, _36851_);
  nand (_39010_, _39009_, _31889_);
  or (_39011_, _39009_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39012_, _39011_, _31965_);
  and (_39013_, _39012_, _39010_);
  nand (_39014_, _38676_, _37896_);
  or (_39015_, _38676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_39016_, _39015_, _31301_);
  and (_39017_, _39016_, _39014_);
  and (_39018_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_39019_, _39018_, rst);
  or (_39020_, _39019_, _39017_);
  or (_40058_, _39020_, _39013_);
  and (_39021_, _38685_, _27633_);
  nand (_39022_, _39021_, _31889_);
  or (_39023_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_39024_, _39023_, _31965_);
  and (_39025_, _39024_, _39022_);
  nand (_39026_, _38692_, _37941_);
  and (_39027_, _39026_, _31301_);
  and (_39028_, _39027_, _39023_);
  not (_39029_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_39030_, _31300_, _39029_);
  or (_39031_, _39030_, rst);
  or (_39032_, _39031_, _39028_);
  or (_40060_, _39032_, _39025_);
  and (_39033_, _38685_, _33228_);
  nand (_39034_, _39033_, _31889_);
  or (_39035_, _39033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39036_, _39035_, _31965_);
  and (_39037_, _39036_, _39034_);
  nand (_39038_, _38692_, _37934_);
  or (_39039_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39040_, _39039_, _31301_);
  and (_39041_, _39040_, _39038_);
  and (_39042_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_39043_, _39042_, rst);
  or (_39044_, _39043_, _39041_);
  or (_40062_, _39044_, _39037_);
  and (_39045_, _38685_, _33979_);
  nand (_39046_, _39045_, _31889_);
  or (_39047_, _39045_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39048_, _39047_, _31965_);
  and (_39049_, _39048_, _39046_);
  nand (_39050_, _38692_, _37927_);
  or (_39051_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_39052_, _39051_, _31301_);
  and (_39053_, _39052_, _39050_);
  and (_39054_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_39055_, _39054_, rst);
  or (_39056_, _39055_, _39053_);
  or (_40064_, _39056_, _39049_);
  and (_39057_, _38685_, _34653_);
  nand (_39058_, _39057_, _31889_);
  or (_39059_, _39057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39060_, _39059_, _31965_);
  and (_39061_, _39060_, _39058_);
  nand (_39062_, _38692_, _37920_);
  or (_39063_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39064_, _39063_, _31301_);
  and (_39065_, _39064_, _39062_);
  and (_39066_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_39067_, _39066_, rst);
  or (_39068_, _39067_, _39065_);
  or (_40066_, _39068_, _39061_);
  and (_39069_, _38685_, _35317_);
  nand (_39070_, _39069_, _31889_);
  or (_39071_, _39069_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39072_, _39071_, _31965_);
  and (_39073_, _39072_, _39070_);
  nand (_39074_, _38692_, _37912_);
  or (_39075_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_39076_, _39075_, _31301_);
  and (_39077_, _39076_, _39074_);
  and (_39078_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_39079_, _39078_, rst);
  or (_39080_, _39079_, _39077_);
  or (_40068_, _39080_, _39073_);
  and (_39081_, _38685_, _36112_);
  nand (_39082_, _39081_, _31889_);
  or (_39083_, _39081_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39084_, _39083_, _31965_);
  and (_39085_, _39084_, _39082_);
  nand (_39086_, _38692_, _37904_);
  or (_39087_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_39088_, _39087_, _31301_);
  and (_39089_, _39088_, _39086_);
  and (_39090_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_39091_, _39090_, rst);
  or (_39092_, _39091_, _39089_);
  or (_40070_, _39092_, _39085_);
  and (_39093_, _38685_, _36851_);
  nand (_39094_, _39093_, _31889_);
  or (_39095_, _39093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39096_, _39095_, _31965_);
  and (_39097_, _39096_, _39094_);
  nand (_39098_, _38692_, _37896_);
  or (_39099_, _38692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_39100_, _39099_, _31301_);
  and (_39101_, _39100_, _39098_);
  and (_39102_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_39103_, _39102_, rst);
  or (_39104_, _39103_, _39101_);
  or (_40072_, _39104_, _39097_);
  nand (_39105_, _38708_, _31889_);
  or (_39106_, _38708_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_39107_, _39106_, _31965_);
  and (_39108_, _39107_, _39105_);
  nor (_39109_, _38709_, _37941_);
  not (_39110_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_39111_, _38708_, _39110_);
  or (_39112_, _39111_, _39109_);
  and (_39113_, _39112_, _31301_);
  nor (_39114_, _31300_, _39110_);
  or (_39115_, _39114_, rst);
  or (_39116_, _39115_, _39113_);
  or (_40074_, _39116_, _39108_);
  and (_39117_, _38701_, _33228_);
  nand (_39118_, _39117_, _31889_);
  or (_39119_, _39117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_39120_, _39119_, _31965_);
  and (_39121_, _39120_, _39118_);
  nor (_39122_, _38709_, _37934_);
  and (_39123_, _38709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39124_, _39123_, _39122_);
  and (_39125_, _39124_, _31301_);
  and (_39126_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_39127_, _39126_, rst);
  or (_39128_, _39127_, _39125_);
  or (_40076_, _39128_, _39121_);
  and (_39129_, _38701_, _33979_);
  nand (_39130_, _39129_, _31889_);
  or (_39131_, _39129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_39132_, _39131_, _31965_);
  and (_39133_, _39132_, _39130_);
  nor (_39134_, _38709_, _37927_);
  and (_39135_, _38709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39136_, _39135_, _39134_);
  and (_39137_, _39136_, _31301_);
  and (_39138_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_39139_, _39138_, rst);
  or (_39140_, _39139_, _39137_);
  or (_40078_, _39140_, _39133_);
  and (_39141_, _38701_, _34653_);
  nand (_39142_, _39141_, _31889_);
  or (_39143_, _39141_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_39144_, _39143_, _31965_);
  and (_39145_, _39144_, _39142_);
  nor (_39146_, _38709_, _37920_);
  and (_39147_, _38709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39148_, _39147_, _39146_);
  and (_39149_, _39148_, _31301_);
  and (_39150_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_39151_, _39150_, rst);
  or (_39152_, _39151_, _39149_);
  or (_40079_, _39152_, _39145_);
  and (_39153_, _38701_, _35317_);
  nand (_39154_, _39153_, _31889_);
  or (_39155_, _39153_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_39156_, _39155_, _31965_);
  and (_39157_, _39156_, _39154_);
  nor (_39158_, _38709_, _37912_);
  and (_39159_, _38709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39160_, _39159_, _39158_);
  and (_39161_, _39160_, _31301_);
  and (_39162_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_39163_, _39162_, rst);
  or (_39164_, _39163_, _39161_);
  or (_40081_, _39164_, _39157_);
  and (_39165_, _38701_, _36112_);
  nand (_39166_, _39165_, _31889_);
  or (_39167_, _39165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_39168_, _39167_, _31965_);
  and (_39169_, _39168_, _39166_);
  nor (_39170_, _38709_, _37904_);
  and (_39171_, _38709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39172_, _39171_, _39170_);
  and (_39173_, _39172_, _31301_);
  and (_39174_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_39175_, _39174_, rst);
  or (_39176_, _39175_, _39173_);
  or (_40083_, _39176_, _39169_);
  and (_39177_, _38701_, _36851_);
  nand (_39178_, _39177_, _31889_);
  or (_39179_, _39177_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_39180_, _39179_, _31965_);
  and (_39181_, _39180_, _39178_);
  nor (_39182_, _38709_, _37896_);
  and (_39183_, _38709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39184_, _39183_, _39182_);
  and (_39185_, _39184_, _31301_);
  and (_39186_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_39187_, _39186_, rst);
  or (_39188_, _39187_, _39185_);
  or (_40085_, _39188_, _39181_);
  and (_39189_, _38717_, _27633_);
  nand (_39190_, _39189_, _31889_);
  or (_39191_, _39189_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_39192_, _39191_, _31965_);
  and (_39193_, _39192_, _39190_);
  nor (_39194_, _38726_, _37941_);
  not (_39195_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_39200_, _38725_, _39195_);
  or (_39206_, _39200_, _39194_);
  and (_39207_, _39206_, _31301_);
  nor (_39208_, _31300_, _39195_);
  or (_39209_, _39208_, rst);
  or (_39210_, _39209_, _39207_);
  or (_40087_, _39210_, _39193_);
  and (_39211_, _38717_, _33228_);
  nand (_39212_, _39211_, _31889_);
  or (_39213_, _39211_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_39214_, _39213_, _31965_);
  and (_39215_, _39214_, _39212_);
  nor (_39216_, _38726_, _37934_);
  and (_39217_, _38726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39218_, _39217_, _39216_);
  and (_39219_, _39218_, _31301_);
  and (_39220_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_39221_, _39220_, rst);
  or (_39222_, _39221_, _39219_);
  or (_40089_, _39222_, _39215_);
  and (_39223_, _38717_, _33979_);
  nand (_39224_, _39223_, _31889_);
  or (_39225_, _39223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_39226_, _39225_, _31965_);
  and (_39227_, _39226_, _39224_);
  nor (_39228_, _38726_, _37927_);
  and (_39229_, _38726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39230_, _39229_, _39228_);
  and (_39231_, _39230_, _31301_);
  and (_39232_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_39233_, _39232_, rst);
  or (_39234_, _39233_, _39231_);
  or (_40091_, _39234_, _39227_);
  and (_39235_, _38717_, _34653_);
  nand (_39236_, _39235_, _31889_);
  or (_39237_, _39235_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_39238_, _39237_, _31965_);
  and (_39239_, _39238_, _39236_);
  nor (_39240_, _38726_, _37920_);
  and (_39241_, _38726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39242_, _39241_, _39240_);
  and (_39243_, _39242_, _31301_);
  and (_39244_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_39245_, _39244_, rst);
  or (_39246_, _39245_, _39243_);
  or (_40093_, _39246_, _39239_);
  and (_39247_, _38717_, _35317_);
  nand (_39248_, _39247_, _31889_);
  or (_39249_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_39250_, _39249_, _31965_);
  and (_39251_, _39250_, _39248_);
  nor (_39252_, _38726_, _37912_);
  and (_39253_, _38726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39254_, _39253_, _39252_);
  and (_39255_, _39254_, _31301_);
  and (_39256_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_39257_, _39256_, rst);
  or (_39258_, _39257_, _39255_);
  or (_40095_, _39258_, _39251_);
  and (_39259_, _38717_, _36112_);
  nand (_39260_, _39259_, _31889_);
  or (_39261_, _39259_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_39262_, _39261_, _31965_);
  and (_39263_, _39262_, _39260_);
  nor (_39264_, _38726_, _37904_);
  and (_39265_, _38726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39266_, _39265_, _39264_);
  and (_39267_, _39266_, _31301_);
  and (_39268_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_39269_, _39268_, rst);
  or (_39270_, _39269_, _39267_);
  or (_40097_, _39270_, _39263_);
  and (_39271_, _38717_, _36851_);
  nand (_39272_, _39271_, _31889_);
  or (_39273_, _39271_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_39274_, _39273_, _31965_);
  and (_39275_, _39274_, _39272_);
  nor (_39276_, _38726_, _37896_);
  and (_39277_, _38726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39278_, _39277_, _39276_);
  and (_39279_, _39278_, _31301_);
  and (_39280_, _38681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_39281_, _39280_, rst);
  or (_39282_, _39281_, _39279_);
  or (_40099_, _39282_, _39275_);
  and (_40549_, t0_i, _42355_);
  and (_40552_, t1_i, _42355_);
  not (_39283_, _31301_);
  nor (_39284_, _39283_, _28290_);
  and (_39285_, _39284_, _34653_);
  and (_39286_, _39285_, _37882_);
  nand (_39287_, _39286_, _37963_);
  nor (_39288_, _27369_, _28290_);
  and (_39289_, _39288_, _33217_);
  and (_39290_, _39289_, _37882_);
  and (_39291_, _39290_, _31301_);
  not (_39292_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_39293_, _39292_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39304_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_39315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39304_);
  nor (_39326_, _39315_, _39293_);
  nor (_39337_, _39326_, _39291_);
  not (_39348_, _39337_);
  and (_39355_, _39348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_39357_, t1_i);
  and (_39358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39357_);
  nor (_39359_, _39358_, _39356_);
  not (_39360_, _39359_);
  not (_39361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_39362_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39361_);
  nor (_39363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_39364_, _39363_);
  and (_39365_, _39364_, _39362_);
  and (_39366_, _39365_, _39360_);
  not (_39367_, _39366_);
  nand (_39368_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_39369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_39370_, _39369_, _39368_);
  nor (_39371_, _39370_, _39367_);
  and (_39372_, _39371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_39373_, _39372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_39374_, _39373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_39375_, _39374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_39376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_39377_, _39370_, _39376_);
  and (_39378_, _39377_, _39366_);
  and (_39379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_39380_, _39379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_39381_, _39380_, _39378_);
  nor (_39382_, _39381_, _39326_);
  and (_39383_, _39382_, _39375_);
  and (_39384_, _39381_, _39293_);
  and (_39385_, _39384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39386_, _39385_, _39383_);
  nor (_39387_, _39386_, _39291_);
  or (_39388_, _39387_, _39355_);
  or (_39389_, _39286_, _39388_);
  and (_39390_, _39389_, _42355_);
  and (_40555_, _39390_, _39287_);
  nand (_39391_, _39291_, _37963_);
  not (_39392_, _39286_);
  and (_39393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39394_, _39393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39395_, _39394_, _39378_);
  and (_39396_, _39395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_39397_, _39396_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39398_, _39397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_39399_, _39398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_39400_, _39399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_39401_, _39399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_39402_, _39401_, _39380_);
  not (_39403_, _39315_);
  nor (_39404_, _39380_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_39405_, _39404_, _39403_);
  nor (_39406_, _39405_, _39402_);
  and (_39407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_39408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39409_, _39408_);
  nor (_39410_, _39401_, _39409_);
  or (_39411_, _39410_, _39407_);
  or (_39412_, _39411_, _39406_);
  and (_39413_, _39412_, _39400_);
  or (_39414_, _39413_, _39291_);
  and (_39415_, _39414_, _39392_);
  and (_39416_, _39415_, _39391_);
  and (_39417_, _39284_, _38100_);
  and (_39419_, _39417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_39425_, _39419_, _39416_);
  and (_40558_, _39425_, _42355_);
  and (_39426_, _39367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_39427_, _39426_, _39402_);
  and (_39428_, _39427_, _39315_);
  or (_39429_, _39426_, _39401_);
  and (_39430_, _39429_, _39408_);
  nand (_39431_, _39366_, _39292_);
  and (_39432_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_39433_, _39432_, _39431_);
  or (_39434_, _39433_, _39384_);
  or (_39435_, _39434_, _39430_);
  or (_39436_, _39435_, _39428_);
  nor (_39437_, _39291_, rst);
  and (_39438_, _39437_, _39392_);
  and (_40561_, _39438_, _39436_);
  and (_39439_, _39284_, _35317_);
  and (_39440_, _39439_, _37882_);
  nor (_39441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_39442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_39443_, t0_i);
  and (_39444_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39443_);
  nor (_39445_, _39444_, _39442_);
  not (_39446_, _39445_);
  not (_39447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_39448_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_39449_, _39448_, _39447_);
  and (_39450_, _39449_, _39446_);
  and (_39451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_39452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39453_, _39452_, _39451_);
  and (_39454_, _39453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_39455_, _39454_, _39450_);
  and (_39456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_39457_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_39458_, _39457_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39459_, _39458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_39460_, _39459_, _39456_);
  and (_39461_, _39460_, _39455_);
  and (_39462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_39463_, _39462_, _39461_);
  and (_39464_, _39463_, _39441_);
  not (_39465_, _39450_);
  and (_39466_, _39465_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_39467_, _39462_, _39460_);
  or (_39468_, _39467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_39469_, _39441_);
  and (_39470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_39471_, _39470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_39472_, _39471_, _39455_);
  and (_39473_, _39472_, _39469_);
  and (_39474_, _39473_, _39468_);
  or (_39475_, _39474_, _39466_);
  or (_39476_, _39475_, _39464_);
  nand (_39477_, _39476_, _42355_);
  nor (_39478_, _39477_, _39440_);
  and (_39479_, _39284_, _33979_);
  and (_39480_, _39479_, _37882_);
  not (_39481_, _39480_);
  and (_40564_, _39481_, _39478_);
  nand (_39482_, _39480_, _37963_);
  not (_39483_, _39440_);
  or (_39484_, _39483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_39485_, _39441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_39486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_39487_, _39486_, _39455_);
  or (_39488_, _39487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_39489_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_39490_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _39489_);
  nand (_39491_, _39490_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_39492_, _39491_, _39472_);
  and (_39493_, _39492_, _39469_);
  or (_39494_, _39493_, _39440_);
  and (_39495_, _39494_, _39488_);
  or (_39496_, _39495_, _39485_);
  and (_39497_, _39496_, _39484_);
  or (_39498_, _39497_, _39480_);
  and (_39499_, _39498_, _42355_);
  and (_40567_, _39499_, _39482_);
  nand (_39500_, _39440_, _37963_);
  and (_39501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _39489_);
  or (_39505_, _39490_, _39501_);
  not (_39513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_39514_, _39471_, _39454_);
  and (_39515_, _39450_, _39489_);
  and (_39516_, _39515_, _39514_);
  and (_39517_, _39516_, _39460_);
  and (_39518_, _39517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_39519_, _39518_, _39513_);
  and (_39520_, _39518_, _39513_);
  or (_39521_, _39520_, _39519_);
  and (_39522_, _39521_, _39505_);
  and (_39523_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39524_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_39525_, _39524_, _39459_);
  and (_39526_, _39525_, _39456_);
  and (_39527_, _39526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_39528_, _39527_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_39529_, _39524_, _39467_);
  and (_39530_, _39529_, _39528_);
  and (_39531_, _39530_, _39523_);
  and (_39532_, _39461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_39533_, _39532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_39534_, _39463_, _39469_);
  and (_39535_, _39534_, _39533_);
  or (_39536_, _39535_, _39531_);
  or (_39537_, _39536_, _39522_);
  or (_39538_, _39537_, _39440_);
  and (_39539_, _39538_, _39481_);
  and (_39540_, _39539_, _39500_);
  and (_39541_, _39480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_39542_, _39541_, _39540_);
  and (_40570_, _39542_, _42355_);
  not (_39543_, _39524_);
  or (_39544_, _39543_, _39467_);
  or (_39545_, _39524_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_39546_, _39523_, _42355_);
  and (_39547_, _39546_, _39545_);
  nand (_39548_, _39547_, _39544_);
  nor (_39549_, _39548_, _39440_);
  and (_40573_, _39549_, _39481_);
  nor (_39550_, _31900_, _28290_);
  and (_39551_, _39550_, _37883_);
  and (_39552_, _39551_, _31301_);
  or (_39553_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_39554_, _39553_, _42355_);
  nand (_39555_, _39552_, _37963_);
  and (_40576_, _39555_, _39554_);
  not (_39556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_39557_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_39558_, _39557_, _39291_);
  and (_39559_, _39558_, _39366_);
  nor (_39560_, _39559_, _39556_);
  and (_39561_, _39559_, _39556_);
  or (_39562_, _39561_, _39560_);
  and (_39563_, _39380_, _39377_);
  and (_39564_, _39563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_39565_, _39564_, _39293_);
  nor (_39566_, _39565_, _39291_);
  or (_39567_, _39566_, _39286_);
  or (_39568_, _39567_, _39562_);
  nand (_39569_, _39286_, _37941_);
  and (_39570_, _39569_, _42355_);
  and (_41062_, _39570_, _39568_);
  and (_39571_, _39366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_39572_, _39571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_39573_, _39571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_39574_, _39573_, _39572_);
  nand (_39575_, _39574_, _39558_);
  or (_39576_, _39558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_39577_, _39576_, _39575_);
  nand (_39578_, _39384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_39579_, _39578_, _39291_);
  or (_39580_, _39579_, _39417_);
  or (_39581_, _39580_, _39577_);
  nand (_39586_, _39417_, _37934_);
  and (_39587_, _39586_, _42355_);
  and (_41064_, _39587_, _39581_);
  not (_39588_, _39417_);
  nor (_39589_, _39572_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_39590_, _39572_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_39591_, _39590_, _39589_);
  and (_39592_, _39591_, _39558_);
  not (_39593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_39594_, _39558_, _39593_);
  nand (_39595_, _39384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_39596_, _39595_, _39291_);
  or (_39597_, _39596_, _39594_);
  or (_39598_, _39597_, _39592_);
  and (_39599_, _39598_, _39588_);
  nor (_39600_, _39588_, _37927_);
  or (_39601_, _39600_, _39599_);
  and (_41066_, _39601_, _42355_);
  not (_39611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_39612_, _39558_, _39611_);
  or (_39613_, _39590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_39614_, _39557_, _39371_);
  and (_39615_, _39614_, _39613_);
  and (_39616_, _39384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_39617_, _39616_, _39615_);
  nor (_39618_, _39617_, _39291_);
  or (_39619_, _39618_, _39612_);
  and (_39620_, _39619_, _39588_);
  nor (_39621_, _39588_, _37920_);
  or (_39622_, _39621_, _39620_);
  and (_41067_, _39622_, _42355_);
  nor (_39623_, _39371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_39624_, _39623_, _39378_);
  and (_39625_, _39624_, _39558_);
  nor (_39626_, _39558_, _39376_);
  nand (_39627_, _39384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_39628_, _39627_, _39291_);
  or (_39629_, _39628_, _39626_);
  or (_39630_, _39629_, _39625_);
  and (_39631_, _39630_, _39588_);
  nor (_39632_, _39588_, _37912_);
  or (_39633_, _39632_, _39631_);
  and (_41069_, _39633_, _42355_);
  nand (_39634_, _39286_, _37904_);
  and (_39635_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_39636_, _39378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_39637_, _39636_, _39635_);
  and (_39638_, _39637_, _39337_);
  and (_39639_, _39348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand (_39640_, _39384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_39641_, _39640_, _39291_);
  or (_39642_, _39641_, _39639_);
  or (_39643_, _39642_, _39638_);
  or (_39644_, _39643_, _39286_);
  and (_39645_, _39644_, _42355_);
  and (_41071_, _39645_, _39634_);
  nand (_39646_, _39286_, _37896_);
  and (_39647_, _39348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_39648_, _39293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_39649_, _39648_, _39366_);
  and (_39650_, _39649_, _39563_);
  nor (_39651_, _39635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_39652_, _39651_, _39326_);
  nor (_39653_, _39652_, _39374_);
  nor (_39654_, _39653_, _39650_);
  nor (_39655_, _39654_, _39291_);
  or (_39656_, _39655_, _39647_);
  or (_39657_, _39656_, _39286_);
  and (_39658_, _39657_, _42355_);
  and (_41073_, _39658_, _39646_);
  nand (_39659_, _39291_, _37941_);
  not (_39660_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_39661_, _39378_, _39304_);
  nor (_39662_, _39380_, _39292_);
  not (_39663_, _39662_);
  and (_39664_, _39663_, _39661_);
  nor (_39665_, _39664_, _39660_);
  and (_39666_, _39664_, _39660_);
  or (_39667_, _39666_, _39665_);
  or (_39668_, _39667_, _39291_);
  and (_39669_, _39668_, _39659_);
  or (_39670_, _39669_, _39417_);
  nand (_39671_, _39417_, _39660_);
  and (_39672_, _39671_, _42355_);
  and (_41075_, _39672_, _39670_);
  nand (_39673_, _39291_, _37934_);
  nor (_39674_, _39381_, _39403_);
  not (_39675_, _39674_);
  nor (_39676_, _39661_, _39315_);
  nor (_39677_, _39676_, _39660_);
  and (_39678_, _39677_, _39675_);
  or (_39679_, _39678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_39680_, _39678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_39681_, _39680_, _39679_);
  or (_39682_, _39681_, _39291_);
  and (_39683_, _39682_, _39392_);
  and (_39684_, _39683_, _39673_);
  and (_39685_, _39286_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_39686_, _39685_, _39684_);
  and (_41077_, _39686_, _42355_);
  nand (_39687_, _39291_, _37927_);
  nand (_39688_, _39395_, _39304_);
  or (_39689_, _39688_, _39662_);
  and (_39690_, _39689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_39691_, _39662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_39692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39693_, _39393_, _39692_);
  nand (_39694_, _39693_, _39378_);
  nor (_39695_, _39694_, _39691_);
  or (_39696_, _39695_, _39690_);
  or (_39697_, _39696_, _39291_);
  and (_39698_, _39697_, _39392_);
  and (_39699_, _39698_, _39687_);
  and (_39700_, _39286_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_39701_, _39700_, _39699_);
  and (_41079_, _39701_, _42355_);
  nand (_39702_, _39291_, _37920_);
  and (_39703_, _39395_, _39380_);
  nor (_39704_, _39703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_39705_, _39396_, _39380_);
  nor (_39706_, _39705_, _39704_);
  or (_39707_, _39706_, _39403_);
  nor (_39708_, _39688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_39709_, _39688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39710_, _39709_, _39315_);
  or (_39711_, _39710_, _39708_);
  and (_39712_, _39711_, _39707_);
  or (_39713_, _39712_, _39291_);
  and (_39714_, _39713_, _39392_);
  and (_39715_, _39714_, _39702_);
  and (_39716_, _39286_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39717_, _39716_, _39715_);
  and (_41081_, _39717_, _42355_);
  nand (_39718_, _39291_, _37912_);
  or (_39719_, _39705_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39720_, _39705_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_39721_, _39720_, _39403_);
  and (_39722_, _39721_, _39719_);
  and (_39723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39724_, _39393_, _39377_);
  and (_39725_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_39726_, _39725_, _39366_);
  and (_39727_, _39726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_39728_, _39727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_39729_, _39727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_39730_, _39729_, _39728_);
  and (_39731_, _39730_, _39408_);
  or (_39732_, _39731_, _39723_);
  or (_39733_, _39732_, _39722_);
  or (_39734_, _39733_, _39291_);
  and (_39735_, _39734_, _39392_);
  and (_39736_, _39735_, _39718_);
  and (_39737_, _39417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_39738_, _39737_, _39736_);
  and (_41083_, _39738_, _42355_);
  nand (_39739_, _39291_, _37904_);
  and (_39740_, _39397_, _39408_);
  and (_39741_, _39720_, _39315_);
  nor (_39742_, _39741_, _39740_);
  nor (_39743_, _39742_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_39744_, _39742_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_39745_, _39744_, _39743_);
  or (_39746_, _39745_, _39291_);
  and (_39747_, _39746_, _39392_);
  and (_39748_, _39747_, _39739_);
  and (_39749_, _39286_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_39750_, _39749_, _39748_);
  and (_41084_, _39750_, _42355_);
  nand (_39751_, _39291_, _37896_);
  not (_39752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  not (_39753_, _39691_);
  nand (_39754_, _39753_, _39398_);
  nand (_39755_, _39754_, _39752_);
  or (_39756_, _39754_, _39752_);
  and (_39757_, _39756_, _39755_);
  or (_39758_, _39757_, _39291_);
  and (_39759_, _39758_, _39392_);
  and (_39760_, _39759_, _39751_);
  and (_39761_, _39417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_39762_, _39761_, _39760_);
  and (_41086_, _39762_, _42355_);
  nor (_39763_, _39465_, _39440_);
  or (_39764_, _39763_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39765_, _39450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_39766_, _39490_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_39767_, _39766_, _39514_);
  nand (_39768_, _39767_, _39765_);
  or (_39769_, _39768_, _39440_);
  and (_39770_, _39769_, _39764_);
  or (_39771_, _39770_, _39480_);
  nand (_39772_, _39480_, _37941_);
  and (_39773_, _39772_, _42355_);
  and (_41088_, _39773_, _39771_);
  nor (_39774_, _39765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_39775_, _39765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_39776_, _39775_, _39774_);
  and (_39777_, _39490_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_39778_, _39777_, _39472_);
  nor (_39779_, _39778_, _39776_);
  nor (_39780_, _39779_, _39440_);
  and (_39781_, _39440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_39782_, _39781_, _39780_);
  and (_39783_, _39782_, _39481_);
  nor (_39784_, _39481_, _37934_);
  or (_39785_, _39784_, _39783_);
  and (_41090_, _39785_, _42355_);
  nor (_39786_, _39775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_39787_, _39765_, _39451_);
  nor (_39788_, _39787_, _39786_);
  and (_39789_, _39490_, _39472_);
  and (_39790_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_39791_, _39790_, _39788_);
  nor (_39792_, _39791_, _39440_);
  and (_39793_, _39440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_39794_, _39793_, _39792_);
  and (_39795_, _39794_, _39481_);
  nor (_39796_, _39481_, _37927_);
  or (_39797_, _39796_, _39795_);
  and (_41092_, _39797_, _42355_);
  and (_39798_, _39453_, _39450_);
  nor (_39799_, _39787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_39800_, _39799_, _39798_);
  and (_39801_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_39802_, _39801_, _39800_);
  nor (_39803_, _39802_, _39440_);
  and (_39804_, _39440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_39805_, _39804_, _39803_);
  and (_39806_, _39805_, _39481_);
  nor (_39807_, _39481_, _37920_);
  or (_39808_, _39807_, _39806_);
  and (_41094_, _39808_, _42355_);
  nor (_39809_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_39810_, _39809_, _39455_);
  and (_39811_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_39812_, _39811_, _39810_);
  or (_39813_, _39812_, _39440_);
  or (_39814_, _39483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_39815_, _39814_, _39481_);
  and (_39816_, _39815_, _39813_);
  nor (_39817_, _39481_, _37912_);
  or (_39818_, _39817_, _39816_);
  and (_41096_, _39818_, _42355_);
  and (_39819_, _39284_, _38107_);
  nand (_39820_, _39819_, _37904_);
  not (_39821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_39822_, _39455_, _39469_);
  and (_39823_, _39822_, _39821_);
  and (_39824_, _39789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_39825_, _39824_, _39823_);
  nor (_39826_, _39825_, _39440_);
  and (_39827_, _39822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_39828_, _39827_);
  or (_39829_, _39828_, _39440_);
  and (_39830_, _39829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_39831_, _39830_, _39826_);
  or (_39832_, _39831_, _39819_);
  and (_39833_, _39832_, _42355_);
  and (_41098_, _39833_, _39820_);
  and (_39834_, _39490_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_39835_, _39834_, _39450_);
  and (_39836_, _39835_, _39514_);
  nor (_39837_, _39828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_39838_, _39837_, _39836_);
  nor (_39839_, _39838_, _39440_);
  and (_39840_, _39829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_39841_, _39840_, _39839_);
  and (_39842_, _39841_, _39481_);
  nor (_39843_, _39481_, _37896_);
  or (_39844_, _39843_, _39842_);
  and (_41100_, _39844_, _42355_);
  nor (_39845_, _39516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_39846_, _39516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_39847_, _39846_, _39845_);
  and (_39848_, _39847_, _39505_);
  and (_39849_, _39524_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_39850_, _39524_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_39851_, _39850_, _39523_);
  nor (_39852_, _39851_, _39849_);
  and (_39853_, _39455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_39854_, _39455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_39855_, _39854_, _39441_);
  nor (_39856_, _39855_, _39853_);
  or (_39857_, _39856_, _39852_);
  or (_39858_, _39857_, _39848_);
  or (_39859_, _39858_, _39440_);
  nand (_39860_, _39440_, _37941_);
  and (_39861_, _39860_, _39859_);
  or (_39862_, _39861_, _39480_);
  or (_39863_, _39481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_39864_, _39863_, _42355_);
  and (_41101_, _39864_, _39862_);
  nand (_39865_, _39440_, _37934_);
  or (_39866_, _39846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_39867_, _39514_, _39450_);
  and (_39868_, _39867_, _39457_);
  not (_39869_, _39868_);
  or (_39870_, _39869_, _39490_);
  and (_39871_, _39870_, _39505_);
  and (_39872_, _39871_, _39866_);
  and (_39873_, _39524_, _39457_);
  or (_39874_, _39849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_39875_, _39874_, _39523_);
  nor (_39876_, _39875_, _39873_);
  and (_39877_, _39853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_39878_, _39853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_39879_, _39878_, _39441_);
  nor (_39880_, _39879_, _39877_);
  or (_39881_, _39880_, _39876_);
  or (_39882_, _39881_, _39872_);
  or (_39883_, _39882_, _39440_);
  and (_39884_, _39883_, _39865_);
  or (_39885_, _39884_, _39480_);
  or (_39886_, _39481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_39887_, _39886_, _42355_);
  and (_41103_, _39887_, _39885_);
  nand (_39888_, _39440_, _37927_);
  or (_39889_, _39868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39890_, _39867_, _39458_);
  not (_39891_, _39890_);
  and (_39892_, _39891_, _39501_);
  and (_39893_, _39892_, _39889_);
  or (_39894_, _39877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39895_, _39458_, _39455_);
  nor (_39896_, _39895_, _39469_);
  and (_39897_, _39896_, _39894_);
  and (_39898_, _39873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_39899_, _39898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39900_, _39524_, _39458_);
  nand (_39901_, _39900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_39902_, _39901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39903_, _39902_, _39899_);
  or (_39904_, _39903_, _39897_);
  or (_39905_, _39904_, _39893_);
  nor (_39906_, _39905_, _39440_);
  nor (_39907_, _39906_, _39819_);
  and (_39908_, _39907_, _39888_);
  and (_39909_, _39480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_39910_, _39909_, _39908_);
  and (_41105_, _39910_, _42355_);
  nand (_39911_, _39440_, _37920_);
  not (_39912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_39913_, _39890_, _39489_);
  nor (_39914_, _39913_, _39912_);
  and (_39915_, _39913_, _39912_);
  or (_39916_, _39915_, _39914_);
  and (_39917_, _39916_, _39505_);
  or (_39918_, _39900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_39919_, _39525_);
  and (_39920_, _39919_, _39523_);
  and (_39921_, _39920_, _39918_);
  or (_39922_, _39895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_39923_, _39459_, _39455_);
  nor (_39924_, _39923_, _39469_);
  and (_39925_, _39924_, _39922_);
  or (_39926_, _39925_, _39921_);
  or (_39927_, _39926_, _39917_);
  nor (_39928_, _39927_, _39440_);
  nor (_39929_, _39928_, _39819_);
  and (_39930_, _39929_, _39911_);
  and (_39931_, _39480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_39932_, _39931_, _39930_);
  and (_41107_, _39932_, _42355_);
  nand (_39933_, _39440_, _37912_);
  or (_39934_, _39923_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_39935_, _39877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_39936_, _39935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_39937_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_39938_, _39937_, _39469_);
  and (_39939_, _39938_, _39934_);
  and (_39940_, _39867_, _39459_);
  or (_39941_, _39940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_39942_, _39940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_39943_, _39942_, _39501_);
  and (_39944_, _39943_, _39941_);
  and (_39945_, _39525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_39946_, _39945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_39947_, _39946_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_39948_, _39525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_39949_, _39948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_39950_, _39949_, _39947_);
  or (_39951_, _39950_, _39944_);
  or (_39952_, _39951_, _39939_);
  or (_39953_, _39952_, _39440_);
  and (_39954_, _39953_, _39481_);
  and (_39955_, _39954_, _39933_);
  and (_39956_, _39480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_39957_, _39956_, _39955_);
  and (_41109_, _39957_, _42355_);
  not (_39958_, _39937_);
  nor (_39959_, _39958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_39960_, _39958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_39961_, _39960_, _39959_);
  and (_39962_, _39961_, _39441_);
  nor (_39963_, _39942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_39964_, _39963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_39965_, _39963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_39966_, _39965_, _39505_);
  and (_39967_, _39966_, _39964_);
  not (_39968_, _39526_);
  and (_39969_, _39968_, _39523_);
  or (_39970_, _39948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_39971_, _39970_, _39969_);
  or (_39972_, _39971_, _39967_);
  or (_39973_, _39972_, _39962_);
  or (_39974_, _39973_, _39440_);
  nand (_39975_, _39440_, _37904_);
  and (_39976_, _39975_, _39974_);
  or (_39977_, _39976_, _39480_);
  or (_39978_, _39481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_39979_, _39978_, _42355_);
  and (_41111_, _39979_, _39977_);
  nand (_39980_, _39440_, _37896_);
  or (_39981_, _39517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_39982_, _39981_, _39505_);
  nor (_39983_, _39982_, _39518_);
  or (_39984_, _39526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_39985_, _39527_);
  and (_39986_, _39985_, _39523_);
  and (_39987_, _39986_, _39984_);
  or (_39988_, _39461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_39989_, _39532_, _39469_);
  and (_39990_, _39989_, _39988_);
  or (_39991_, _39990_, _39987_);
  or (_39992_, _39991_, _39983_);
  nor (_39993_, _39992_, _39440_);
  nor (_39994_, _39993_, _39819_);
  and (_39995_, _39994_, _39980_);
  and (_39996_, _39480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_39997_, _39996_, _39995_);
  and (_41113_, _39997_, _42355_);
  nand (_39998_, _39552_, _37941_);
  or (_39999_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_40000_, _39999_, _42355_);
  and (_41115_, _40000_, _39998_);
  or (_40001_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_40002_, _40001_, _42355_);
  nand (_40003_, _39552_, _37934_);
  and (_41117_, _40003_, _40002_);
  or (_40004_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_40005_, _40004_, _42355_);
  nand (_40006_, _39552_, _37927_);
  and (_41118_, _40006_, _40005_);
  or (_40007_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_40008_, _40007_, _42355_);
  nand (_40009_, _39552_, _37920_);
  and (_41120_, _40009_, _40008_);
  or (_40010_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_40011_, _40010_, _42355_);
  nand (_40012_, _39552_, _37912_);
  and (_41122_, _40012_, _40011_);
  or (_40013_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_40014_, _40013_, _42355_);
  nand (_40015_, _39552_, _37904_);
  and (_41124_, _40015_, _40014_);
  or (_40016_, _39552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_40017_, _40016_, _42355_);
  nand (_40018_, _39552_, _37896_);
  and (_41126_, _40018_, _40017_);
  nor (_40019_, _28433_, _28290_);
  and (_40020_, _40019_, _38532_);
  and (_40021_, _40020_, _38700_);
  and (_40022_, _40021_, _31922_);
  nand (_40023_, _40022_, _31889_);
  and (_40024_, _37877_, _31922_);
  and (_40025_, _40024_, _38724_);
  not (_40026_, _40025_);
  or (_40027_, _40022_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_40028_, _40027_, _40026_);
  and (_40029_, _40028_, _40023_);
  not (_40030_, _37963_);
  and (_40031_, _38718_, _31301_);
  and (_40032_, _40031_, _40030_);
  or (_40033_, _40032_, _40029_);
  and (_42293_, _40033_, _42355_);
  and (_40034_, _39284_, _27633_);
  and (_40035_, _40034_, _38707_);
  not (_40036_, _40035_);
  and (_40037_, _28433_, _28301_);
  and (_40038_, _40037_, _38532_);
  and (_40039_, _40038_, _38700_);
  and (_40040_, _40039_, _31922_);
  or (_40041_, _40040_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40042_, _40041_, _40036_);
  nand (_40043_, _40040_, _31889_);
  and (_40044_, _40043_, _40042_);
  nor (_40045_, _40036_, _37963_);
  or (_40046_, _40045_, _40044_);
  and (_42296_, _40046_, _42355_);
  and (_40049_, _40034_, _37882_);
  nor (_40051_, _38531_, _28290_);
  and (_40053_, _40051_, _28433_);
  and (_40055_, _40053_, _28148_);
  and (_40057_, _40055_, _38668_);
  nand (_40059_, _40057_, _27611_);
  and (_40061_, _40059_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40063_, _40061_, _40049_);
  or (_40065_, _27622_, _33968_);
  and (_40067_, _40065_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_40069_, _40067_, _38467_);
  and (_40071_, _40069_, _40057_);
  or (_40073_, _40071_, _40063_);
  nand (_40075_, _40049_, _37896_);
  and (_40077_, _40075_, _42355_);
  and (_42298_, _40077_, _40073_);
  not (_40080_, _40049_);
  nor (_40082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_40084_, _40082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_40086_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_40088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_40090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40090_);
  and (_40094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40096_, _40094_, _40092_);
  nor (_40098_, _40096_, _40088_);
  or (_40100_, _40098_, _40086_);
  and (_40101_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_40102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_40103_, _40102_, _40101_);
  nor (_40104_, _40103_, _40088_);
  and (_40105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40090_);
  and (_40106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40107_, _40106_, _40105_);
  nand (_40108_, _40107_, _40104_);
  or (_40109_, _40108_, _40100_);
  and (_40110_, _40109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_40111_, _40110_, _40084_);
  and (_40112_, _37882_, _31922_);
  and (_40113_, _40112_, _40051_);
  or (_40114_, _40113_, _40111_);
  and (_40115_, _40114_, _40080_);
  nand (_40116_, _40113_, _31889_);
  and (_40117_, _40116_, _40115_);
  nor (_40118_, _40080_, _37963_);
  or (_40119_, _40118_, _40117_);
  and (_42300_, _40119_, _42355_);
  and (_40120_, _39290_, _31965_);
  nand (_40121_, _40120_, _31889_);
  not (_40122_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_40123_, _40122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_40124_, _40107_, _40088_);
  not (_40125_, _40124_);
  or (_40126_, _40125_, _40104_);
  or (_40127_, _40126_, _40100_);
  and (_40128_, _40127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_40129_, _40128_, _40123_);
  or (_40130_, _40129_, _40120_);
  and (_40131_, _40130_, _40121_);
  or (_40132_, _40131_, _40049_);
  nand (_40133_, _40049_, _37904_);
  and (_40134_, _40133_, _42355_);
  and (_42302_, _40134_, _40132_);
  not (_40135_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_40136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40135_);
  nand (_40137_, _40098_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_40138_, _40124_, _40104_);
  or (_40139_, _40138_, _40137_);
  and (_40140_, _40139_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_40141_, _40140_, _40136_);
  and (_40142_, _39551_, _31965_);
  or (_40143_, _40142_, _40141_);
  and (_40144_, _40143_, _40080_);
  nand (_40145_, _40142_, _31889_);
  and (_40146_, _40145_, _40144_);
  nor (_40147_, _40080_, _37934_);
  or (_40148_, _40147_, _40146_);
  and (_42304_, _40148_, _42355_);
  and (_40149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_40150_, _40137_, _40126_);
  and (_40151_, _40150_, _40149_);
  and (_40152_, _40051_, _38100_);
  or (_40153_, _40152_, _40151_);
  and (_40154_, _40153_, _40080_);
  nand (_40155_, _40152_, _31889_);
  and (_40156_, _40155_, _40154_);
  nor (_40157_, _40080_, _37920_);
  or (_40158_, _40157_, _40156_);
  and (_42306_, _40158_, _42355_);
  nand (_40159_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_40160_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40090_);
  and (_40161_, _40160_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_40162_, _40161_, _40159_);
  or (_40163_, _40162_, _40088_);
  and (_40164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40165_, _40164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_40166_, _40165_);
  and (_40167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40168_, _40167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_40169_, _40168_);
  and (_40170_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40171_, _40170_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40173_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_40174_, _40173_, _40171_);
  and (_40175_, _40174_, _40169_);
  and (_40176_, _40175_, _40166_);
  not (_40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_40178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_40179_, _40178_, _40177_);
  nand (_40180_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_40181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_40182_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_40183_, _40182_, _40181_);
  and (_40184_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_40185_, _40184_);
  and (_40186_, _40185_, _40180_);
  nand (_40187_, _40186_, _40176_);
  and (_40188_, _40187_, _40163_);
  and (_40189_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_40190_, _40189_, _40090_);
  and (_40191_, _40190_, _40188_);
  not (_40192_, _40191_);
  not (_40193_, _40190_);
  and (_40194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40088_);
  not (_40195_, _40194_);
  not (_40196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40197_, _40167_, _40196_);
  not (_40198_, _40197_);
  not (_40199_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40200_, _40170_, _40199_);
  not (_40201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40202_, _40172_, _40201_);
  nor (_40203_, _40202_, _40200_);
  and (_40204_, _40203_, _40198_);
  nor (_40205_, _40204_, _40195_);
  not (_40206_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40207_, _40179_, _40206_);
  not (_40208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40209_, _40183_, _40208_);
  nor (_40210_, _40209_, _40207_);
  not (_40211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40212_, _40164_, _40211_);
  not (_40213_, _40212_);
  and (_40214_, _40213_, _40210_);
  nor (_40215_, _40214_, _40195_);
  nor (_40216_, _40215_, _40205_);
  or (_40217_, _40216_, _40193_);
  and (_40218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42355_);
  and (_40219_, _40218_, _40217_);
  and (_42342_, _40219_, _40192_);
  nor (_40220_, _40189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_40221_, _40220_);
  not (_40222_, _40188_);
  and (_40223_, _40216_, _40222_);
  nor (_40224_, _40223_, _40221_);
  nand (_40225_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42355_);
  nor (_42344_, _40225_, _40224_);
  and (_40226_, _40186_, _40166_);
  nand (_40227_, _40226_, _40188_);
  or (_40228_, _40215_, _40188_);
  and (_40229_, _40228_, _40190_);
  and (_40230_, _40229_, _40227_);
  or (_40231_, _40230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_40232_, _40192_, _40175_);
  nor (_40233_, _40193_, _40188_);
  nand (_40234_, _40233_, _40205_);
  and (_40235_, _40234_, _42355_);
  and (_40236_, _40235_, _40232_);
  and (_42345_, _40236_, _40231_);
  and (_40237_, _40227_, _40220_);
  or (_40238_, _40237_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_40239_, _40220_, _40188_);
  not (_40240_, _40239_);
  or (_40241_, _40240_, _40175_);
  or (_40242_, _40215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_40243_, _40220_, _40205_);
  and (_40244_, _40243_, _40242_);
  or (_40245_, _40244_, _40188_);
  and (_40246_, _40245_, _42355_);
  and (_40247_, _40246_, _40241_);
  and (_42347_, _40247_, _40238_);
  nand (_40248_, _40223_, _40088_);
  nor (_40249_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_40250_, _40249_, _40189_);
  and (_40251_, _40250_, _42355_);
  and (_42349_, _40251_, _40248_);
  and (_40252_, _40223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_40253_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_40254_, _40253_, _40249_);
  nor (_40255_, _40254_, _40222_);
  or (_40256_, _40255_, _40189_);
  or (_40257_, _40256_, _40252_);
  not (_40258_, _40189_);
  or (_40259_, _40254_, _40258_);
  and (_40260_, _40259_, _42355_);
  and (_42351_, _40260_, _40257_);
  and (_40261_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42355_);
  and (_42353_, _40261_, _40189_);
  nor (_42358_, _40082_, rst);
  and (_42360_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _42355_);
  nor (_40262_, _40223_, _40189_);
  and (_40263_, _40189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_40264_, _40263_, _40262_);
  and (_00131_, _40264_, _42355_);
  and (_40265_, _40189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_40266_, _40265_, _40262_);
  and (_00133_, _40266_, _42355_);
  and (_40267_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42355_);
  and (_00134_, _40267_, _40189_);
  not (_40268_, _40202_);
  nor (_40269_, _40209_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_40270_, _40269_, _40207_);
  or (_40271_, _40270_, _40212_);
  and (_40272_, _40271_, _40268_);
  or (_40273_, _40272_, _40200_);
  nor (_40274_, _40216_, _40188_);
  and (_40275_, _40274_, _40198_);
  and (_40276_, _40275_, _40273_);
  not (_40277_, _40173_);
  or (_40278_, _40184_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40279_, _40278_, _40180_);
  or (_40280_, _40279_, _40165_);
  and (_40281_, _40280_, _40277_);
  or (_40282_, _40281_, _40171_);
  and (_40283_, _40188_, _40169_);
  and (_40284_, _40283_, _40282_);
  or (_40285_, _40284_, _40189_);
  or (_40286_, _40285_, _40276_);
  or (_40287_, _40258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_40288_, _40287_, _42355_);
  and (_00136_, _40288_, _40286_);
  nor (_40289_, _40200_, _40197_);
  or (_40290_, _40212_, _40202_);
  and (_40291_, _40210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40292_, _40291_, _40290_);
  and (_40293_, _40292_, _40289_);
  and (_40294_, _40293_, _40274_);
  not (_40295_, _40171_);
  or (_40296_, _40173_, _40165_);
  and (_40297_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_40298_, _40297_, _40296_);
  and (_40299_, _40298_, _40295_);
  and (_40300_, _40299_, _40283_);
  or (_40301_, _40300_, _40189_);
  or (_40302_, _40301_, _40294_);
  or (_40303_, _40258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_40304_, _40303_, _42355_);
  and (_00138_, _40304_, _40302_);
  and (_40305_, _40213_, _40194_);
  nand (_40306_, _40305_, _40204_);
  or (_40307_, _40306_, _40210_);
  nor (_40308_, _40307_, _40188_);
  not (_40309_, _40186_);
  and (_40316_, _40309_, _40176_);
  and (_40317_, _40316_, _40163_);
  or (_40323_, _40317_, _40189_);
  or (_40329_, _40323_, _40308_);
  or (_40335_, _40258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_40338_, _40335_, _42355_);
  and (_00140_, _40338_, _40329_);
  and (_40339_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42355_);
  and (_00142_, _40339_, _40189_);
  and (_40340_, _40189_, _40090_);
  or (_40341_, _40340_, _40224_);
  or (_40342_, _40341_, _40233_);
  and (_00144_, _40342_, _42355_);
  not (_40343_, _40262_);
  and (_40344_, _40343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_40345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_40346_, _40184_, _40090_);
  or (_40347_, _40346_, _40345_);
  nor (_40348_, _40180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40349_, _40348_, _40165_);
  nand (_40355_, _40349_, _40347_);
  or (_40356_, _40166_, _40094_);
  and (_40360_, _40356_, _40355_);
  or (_40361_, _40360_, _40173_);
  or (_40363_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40090_);
  or (_40364_, _40363_, _40277_);
  and (_40370_, _40364_, _40295_);
  and (_40373_, _40370_, _40361_);
  and (_40374_, _40171_, _40094_);
  or (_40375_, _40374_, _40168_);
  or (_40378_, _40375_, _40373_);
  or (_40384_, _40363_, _40169_);
  and (_40386_, _40384_, _40188_);
  and (_40387_, _40386_, _40378_);
  and (_40389_, _40209_, _40090_);
  or (_40395_, _40389_, _40345_);
  and (_40398_, _40207_, _40090_);
  nor (_40399_, _40398_, _40212_);
  nand (_40400_, _40399_, _40395_);
  or (_40403_, _40213_, _40094_);
  and (_40409_, _40403_, _40400_);
  or (_40411_, _40409_, _40202_);
  not (_40414_, _40200_);
  or (_40415_, _40363_, _40268_);
  and (_40421_, _40415_, _40414_);
  and (_40423_, _40421_, _40411_);
  and (_40425_, _40200_, _40094_);
  or (_40426_, _40425_, _40197_);
  or (_40432_, _40426_, _40423_);
  and (_40435_, _40363_, _40274_);
  or (_40436_, _40435_, _40275_);
  and (_40438_, _40436_, _40432_);
  or (_40444_, _40438_, _40387_);
  and (_40447_, _40444_, _40258_);
  or (_40448_, _40447_, _40344_);
  and (_00145_, _40448_, _42355_);
  or (_40451_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40090_);
  and (_40457_, _40451_, _40169_);
  or (_40459_, _40457_, _40175_);
  or (_40460_, _40346_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40463_, _40460_, _40349_);
  nand (_40469_, _40165_, _40106_);
  nand (_40471_, _40469_, _40174_);
  or (_40472_, _40471_, _40463_);
  and (_40474_, _40472_, _40459_);
  nand (_40480_, _40168_, _40106_);
  nand (_40483_, _40480_, _40188_);
  or (_40484_, _40483_, _40474_);
  or (_40486_, _40389_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40492_, _40486_, _40399_);
  and (_40495_, _40212_, _40106_);
  or (_40496_, _40495_, _40492_);
  and (_40497_, _40496_, _40203_);
  not (_40502_, _40203_);
  and (_40507_, _40451_, _40502_);
  or (_40508_, _40507_, _40197_);
  or (_40509_, _40508_, _40497_);
  or (_40514_, _40198_, _40106_);
  nand (_40519_, _40514_, _40509_);
  nand (_40520_, _40519_, _40274_);
  and (_40521_, _40520_, _40484_);
  or (_40525_, _40521_, _40189_);
  or (_40531_, _40262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_40532_, _40531_, _42355_);
  and (_00147_, _40532_, _40525_);
  and (_40536_, _40343_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_40541_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40542_, _40541_, _40169_);
  and (_40543_, _40542_, _40188_);
  not (_40544_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_40545_, _40184_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40546_, _40545_, _40544_);
  nor (_40547_, _40180_, _40090_);
  nor (_40548_, _40547_, _40165_);
  nand (_40550_, _40548_, _40546_);
  or (_40551_, _40166_, _40092_);
  and (_40553_, _40551_, _40550_);
  or (_40554_, _40553_, _40173_);
  or (_40556_, _40541_, _40277_);
  and (_40557_, _40556_, _40295_);
  and (_40559_, _40557_, _40554_);
  and (_40560_, _40171_, _40092_);
  or (_40562_, _40560_, _40168_);
  or (_40563_, _40562_, _40559_);
  and (_40565_, _40563_, _40543_);
  or (_40566_, _40541_, _40198_);
  and (_40568_, _40209_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_40569_, _40568_, _40544_);
  and (_40571_, _40207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_40572_, _40571_, _40212_);
  nand (_40574_, _40572_, _40569_);
  or (_40575_, _40213_, _40092_);
  and (_40577_, _40575_, _40574_);
  or (_40578_, _40577_, _40202_);
  or (_40579_, _40541_, _40268_);
  and (_40580_, _40579_, _40414_);
  and (_40581_, _40580_, _40578_);
  and (_40582_, _40200_, _40092_);
  or (_40583_, _40582_, _40197_);
  or (_40584_, _40583_, _40581_);
  and (_40585_, _40584_, _40274_);
  and (_40586_, _40585_, _40566_);
  or (_40587_, _40586_, _40565_);
  and (_40588_, _40587_, _40258_);
  or (_40589_, _40588_, _40536_);
  and (_00149_, _40589_, _42355_);
  or (_40590_, _40545_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40591_, _40590_, _40548_);
  and (_40592_, _40165_, _40105_);
  or (_40593_, _40592_, _40591_);
  and (_40594_, _40593_, _40174_);
  not (_40595_, _40174_);
  or (_40596_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_40597_, _40596_, _40595_);
  or (_40598_, _40597_, _40168_);
  or (_40599_, _40598_, _40594_);
  or (_40600_, _40169_, _40105_);
  and (_40601_, _40600_, _40188_);
  and (_40602_, _40601_, _40599_);
  and (_40603_, _40223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_40604_, _40603_, _40602_);
  or (_40605_, _40568_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40606_, _40605_, _40572_);
  and (_40607_, _40212_, _40105_);
  or (_40608_, _40607_, _40606_);
  and (_40609_, _40608_, _40203_);
  and (_40610_, _40596_, _40502_);
  or (_40611_, _40610_, _40197_);
  or (_40612_, _40611_, _40609_);
  or (_40613_, _40198_, _40105_);
  and (_40614_, _40613_, _40274_);
  and (_40615_, _40614_, _40612_);
  or (_40616_, _40615_, _40189_);
  or (_40617_, _40616_, _40604_);
  or (_40618_, _40258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_40619_, _40618_, _42355_);
  and (_00151_, _40619_, _40617_);
  or (_40620_, _40221_, _40216_);
  and (_40621_, _40620_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_40622_, _40621_, _40239_);
  and (_00153_, _40622_, _42355_);
  and (_40623_, _40217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_40624_, _40623_, _40191_);
  and (_00155_, _40624_, _42355_);
  and (_40625_, _40057_, _27633_);
  or (_40626_, _40625_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40627_, _40626_, _40080_);
  nand (_40628_, _40625_, _31889_);
  and (_40629_, _40628_, _40627_);
  nor (_40630_, _40080_, _37941_);
  or (_40631_, _40630_, _40629_);
  and (_00156_, _40631_, _42355_);
  and (_40632_, _40057_, _33979_);
  or (_40633_, _40632_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_40634_, _40633_, _40080_);
  nand (_40635_, _40632_, _31889_);
  and (_40636_, _40635_, _40634_);
  nor (_40637_, _40080_, _37927_);
  or (_40638_, _40637_, _40636_);
  and (_00158_, _40638_, _42355_);
  and (_40639_, _40057_, _35317_);
  or (_40640_, _40639_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_40641_, _40640_, _40080_);
  nand (_40642_, _40639_, _31889_);
  and (_40643_, _40642_, _40641_);
  nor (_40644_, _40080_, _37912_);
  or (_40645_, _40644_, _40643_);
  and (_00160_, _40645_, _42355_);
  and (_40646_, _40039_, _27633_);
  or (_40647_, _40646_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_40648_, _40647_, _40036_);
  nand (_40649_, _40646_, _31889_);
  and (_40650_, _40649_, _40648_);
  nor (_40651_, _40036_, _37941_);
  or (_40652_, _40651_, _40650_);
  and (_00162_, _40652_, _42355_);
  and (_40653_, _40039_, _33228_);
  or (_40654_, _40653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_40655_, _40654_, _40036_);
  nand (_40656_, _40653_, _31889_);
  and (_40657_, _40656_, _40655_);
  nor (_40658_, _40036_, _37934_);
  or (_40659_, _40658_, _40657_);
  and (_00164_, _40659_, _42355_);
  nand (_40660_, _40039_, _38759_);
  and (_40661_, _40660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40662_, _40661_, _40035_);
  and (_40663_, _34012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40664_, _40663_, _34001_);
  and (_40665_, _40664_, _40039_);
  or (_40666_, _40665_, _40662_);
  nand (_40667_, _40035_, _37927_);
  and (_40668_, _40667_, _42355_);
  and (_00166_, _40668_, _40666_);
  and (_40669_, _40039_, _34653_);
  or (_40670_, _40669_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_40671_, _40670_, _40036_);
  nand (_40672_, _40669_, _31889_);
  and (_40673_, _40672_, _40671_);
  nor (_40674_, _40036_, _37920_);
  or (_40675_, _40674_, _40673_);
  and (_00167_, _40675_, _42355_);
  and (_40676_, _40039_, _35317_);
  or (_40677_, _40676_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_40678_, _40677_, _40036_);
  nand (_40679_, _40676_, _31889_);
  and (_40680_, _40679_, _40678_);
  nor (_40681_, _40036_, _37912_);
  or (_40682_, _40681_, _40680_);
  and (_00169_, _40682_, _42355_);
  and (_40683_, _40039_, _36112_);
  or (_40684_, _40683_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_40685_, _40684_, _40036_);
  nand (_40686_, _40683_, _31889_);
  and (_40687_, _40686_, _40685_);
  nor (_40688_, _40036_, _37904_);
  or (_40689_, _40688_, _40687_);
  and (_00171_, _40689_, _42355_);
  and (_40690_, _40039_, _36851_);
  or (_40691_, _40690_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_40692_, _40691_, _40036_);
  nand (_40693_, _40690_, _31889_);
  and (_40694_, _40693_, _40692_);
  nor (_40695_, _40036_, _37896_);
  or (_40696_, _40695_, _40694_);
  and (_00173_, _40696_, _42355_);
  and (_40697_, _40021_, _27633_);
  nand (_40698_, _40697_, _31889_);
  or (_40699_, _40697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40700_, _40699_, _40026_);
  and (_40701_, _40700_, _40698_);
  and (_40702_, _40031_, _37942_);
  or (_40703_, _40702_, _40701_);
  and (_00175_, _40703_, _42355_);
  and (_40704_, _40021_, _33228_);
  nand (_40705_, _40704_, _31889_);
  or (_40706_, _40704_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40707_, _40706_, _40026_);
  and (_40708_, _40707_, _40705_);
  not (_40709_, _37934_);
  and (_40710_, _40031_, _40709_);
  or (_40711_, _40710_, _40708_);
  and (_00177_, _40711_, _42355_);
  and (_40712_, _34012_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40713_, _40712_, _34001_);
  and (_40714_, _40713_, _40021_);
  nand (_40715_, _40021_, _38759_);
  and (_40716_, _40715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_40717_, _40716_, _40025_);
  or (_40718_, _40717_, _40714_);
  nand (_40719_, _40025_, _37927_);
  and (_40720_, _40719_, _42355_);
  and (_00178_, _40720_, _40718_);
  and (_40721_, _40021_, _34653_);
  nand (_40722_, _40721_, _31889_);
  or (_40723_, _40721_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_40724_, _40723_, _40026_);
  and (_40725_, _40724_, _40722_);
  not (_40726_, _37920_);
  and (_40727_, _40031_, _40726_);
  or (_40728_, _40727_, _40725_);
  and (_00180_, _40728_, _42355_);
  and (_40729_, _40021_, _35317_);
  nand (_40730_, _40729_, _31889_);
  or (_40731_, _40729_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40732_, _40731_, _40026_);
  and (_40733_, _40732_, _40730_);
  not (_40734_, _37912_);
  and (_40735_, _40031_, _40734_);
  or (_40736_, _40735_, _40733_);
  and (_00182_, _40736_, _42355_);
  and (_40737_, _40021_, _36112_);
  nand (_40738_, _40737_, _31889_);
  or (_40739_, _40737_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40740_, _40739_, _40026_);
  and (_40741_, _40740_, _40738_);
  not (_40742_, _37904_);
  and (_40743_, _40031_, _40742_);
  or (_40744_, _40743_, _40741_);
  and (_00184_, _40744_, _42355_);
  and (_40745_, _40021_, _36851_);
  and (_40746_, _40745_, _31889_);
  nor (_40747_, _40745_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_40748_, _40747_, _40746_);
  nand (_40749_, _40748_, _40026_);
  nand (_40750_, _40025_, _37896_);
  and (_40751_, _40750_, _42355_);
  and (_00186_, _40751_, _40749_);
  and (_40752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_40753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_40754_, _40082_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_40755_, _40754_, _40753_);
  not (_40756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_40757_, _40756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_40758_, _40757_, _40755_);
  nor (_40759_, _40758_, _40752_);
  or (_40760_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_40761_, _40760_, _42355_);
  nor (_00546_, _40761_, _40759_);
  nor (_40762_, _40759_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_40763_, _40762_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_40764_, _40762_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_40765_, _40764_, _42355_);
  and (_00549_, _40765_, _40763_);
  not (_40766_, rxd_i);
  and (_40767_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _40766_);
  nor (_40768_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_40769_, _40768_);
  and (_40770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_40771_, _40770_, _40769_);
  and (_40772_, _40771_, _40767_);
  not (_40773_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_40774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _40773_);
  and (_40775_, _40774_, _40768_);
  or (_40776_, _40775_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_40777_, _40776_, _40772_);
  and (_40778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _42355_);
  and (_00551_, _40778_, _40777_);
  and (_40779_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_40780_, _40779_, _40769_);
  not (_40781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_40782_, _40768_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_40783_, _40782_, _40781_);
  nor (_40784_, _40783_, _40780_);
  not (_40785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_40786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _40785_);
  not (_40787_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_40788_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _40787_);
  and (_40789_, _40788_, _40786_);
  not (_40790_, _40789_);
  or (_40791_, _40790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_40792_, _40789_, _40780_);
  and (_40793_, _40780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_40794_, _40793_, _40792_);
  and (_40795_, _40794_, _40791_);
  or (_40796_, _40795_, _40784_);
  and (_40797_, _40768_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_40798_, _40797_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not (_40799_, _40798_);
  or (_40800_, _40799_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_40801_, _40800_, _40796_);
  nand (_00554_, _40801_, _40778_);
  not (_40802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_40803_, _40780_);
  nor (_40804_, _40781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_40805_, _40804_);
  not (_40806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_40807_, _40768_, _40806_);
  and (_40808_, _40807_, _40805_);
  and (_40809_, _40808_, _40803_);
  nor (_40810_, _40809_, _40802_);
  and (_40811_, _40809_, rxd_i);
  or (_40812_, _40811_, rst);
  or (_00557_, _40812_, _40810_);
  nor (_40813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_40814_, _40813_, _40786_);
  and (_40815_, _40814_, _40793_);
  nand (_40816_, _40815_, _40766_);
  or (_40817_, _40815_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_40818_, _40817_, _42355_);
  and (_00559_, _40818_, _40816_);
  and (_40819_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_40820_, _40819_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_40821_, _40820_, _40785_);
  and (_40822_, _40821_, _40793_);
  and (_40823_, _40771_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_40824_, _40823_, _40793_);
  nor (_40825_, _40820_, _40803_);
  or (_40826_, _40825_, _40824_);
  and (_40827_, _40826_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_40828_, _40827_, _40822_);
  and (_00562_, _40828_, _42355_);
  and (_40829_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _42355_);
  nand (_40830_, _40829_, _40806_);
  nand (_40831_, _40778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_00565_, _40831_, _40830_);
  and (_40832_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _40806_);
  not (_40833_, _40771_);
  not (_40834_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_40835_, _40775_, _40834_);
  and (_40836_, _40835_, _40833_);
  and (_40837_, _40836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_40838_, _40837_, _40780_);
  or (_40839_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_40840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_40841_, _40840_, _40792_);
  and (_40842_, _40841_, _40839_);
  and (_40843_, _40842_, _40838_);
  or (_40844_, _40843_, _40798_);
  nand (_40845_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_40846_, _40845_, _40780_);
  or (_40847_, _40846_, _40790_);
  and (_40848_, _40847_, _40799_);
  or (_40849_, _40848_, rxd_i);
  and (_40850_, _40849_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_40851_, _40850_, _40844_);
  or (_40852_, _40851_, _40832_);
  and (_00567_, _40852_, _42355_);
  and (_40853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_40854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_40855_, _40754_, _40854_);
  or (_40856_, _40855_, _40757_);
  nor (_40857_, _40856_, _40853_);
  or (_40858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_40859_, _40858_, _42355_);
  nor (_00570_, _40859_, _40857_);
  nor (_40860_, _40857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_40861_, _40860_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_40862_, _40860_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_40863_, _40862_, _42355_);
  and (_00573_, _40863_, _40861_);
  and (_40864_, _40797_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_40865_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_40866_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_40867_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_40868_, _40867_, _40866_);
  and (_40869_, _40868_, _40865_);
  not (_40870_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_40871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_40872_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_40873_, _40872_, _40871_);
  and (_40874_, _40873_, _40870_);
  and (_40875_, _40874_, _40869_);
  or (_40876_, _40875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_40877_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_40878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_40879_, _40878_, _40877_);
  and (_40880_, _40769_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_40881_, _40880_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_40882_, _40881_, _40879_);
  not (_40883_, _40882_);
  or (_40884_, _40883_, _40876_);
  and (_40885_, _40879_, _40880_);
  not (_40886_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or (_40887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _40886_);
  or (_40888_, _40887_, _40885_);
  and (_40889_, _40888_, _40884_);
  or (_40890_, _40889_, _40864_);
  not (_40891_, _40864_);
  not (_40892_, _40875_);
  or (_40893_, _40892_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_40894_, _40893_, _40876_);
  or (_40895_, _40894_, _40891_);
  nand (_40896_, _40895_, _40890_);
  and (_40897_, _39550_, _33217_);
  and (_40898_, _40897_, _31301_);
  and (_40899_, _40898_, _38691_);
  nor (_40900_, _40899_, rst);
  nand (_40901_, _40900_, _40896_);
  not (_40902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_40903_, _40899_, _42355_);
  nand (_40904_, _40903_, _40902_);
  and (_00575_, _40904_, _40901_);
  nor (_40905_, _40892_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_40906_, _40885_, _40905_);
  and (_40907_, _40875_, _40864_);
  or (_40908_, _40886_, rst);
  nor (_40909_, _40908_, _40907_);
  and (_40910_, _40909_, _40906_);
  or (_00578_, _40910_, _40903_);
  or (_40911_, _40883_, _40905_);
  or (_40912_, _40885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_40913_, _40797_, _40886_);
  and (_40914_, _40913_, _40912_);
  and (_40915_, _40914_, _40911_);
  or (_40916_, _40915_, _40907_);
  and (_00581_, _40916_, _40900_);
  and (_40917_, _40881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_40918_, _40917_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_40919_, _40918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_40920_, _40919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_40921_, _40919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_40922_, _40921_, _40920_);
  and (_00583_, _40922_, _40900_);
  and (_40923_, _40903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_40924_, _40882_, _40864_);
  and (_40925_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_40926_, _40925_, _40900_);
  or (_00586_, _40926_, _40923_);
  and (_40927_, _40024_, _37882_);
  or (_40928_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_40929_, _40928_, _42355_);
  nand (_40930_, _40927_, _37963_);
  and (_00589_, _40930_, _40929_);
  and (_40931_, _40020_, _38668_);
  and (_40932_, _40931_, _31922_);
  nand (_40933_, _40932_, _31889_);
  and (_40934_, _40034_, _38691_);
  not (_40935_, _40934_);
  or (_40936_, _40932_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_40937_, _40936_, _40935_);
  and (_40938_, _40937_, _40933_);
  nor (_40939_, _40935_, _37963_);
  or (_40940_, _40939_, _40938_);
  and (_00591_, _40940_, _42355_);
  nor (_40941_, _40798_, _40792_);
  not (_40942_, _40941_);
  nor (_40943_, _40836_, _40780_);
  nor (_40944_, _40943_, _40942_);
  nor (_40945_, _40944_, _40806_);
  or (_40946_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_40947_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _40806_);
  or (_40948_, _40947_, _40941_);
  and (_40949_, _40948_, _42355_);
  and (_01209_, _40949_, _40946_);
  or (_40950_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_40951_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _40806_);
  or (_40952_, _40951_, _40941_);
  and (_40953_, _40952_, _42355_);
  and (_01211_, _40953_, _40950_);
  or (_40954_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_40955_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _40806_);
  or (_40956_, _40955_, _40941_);
  and (_40957_, _40956_, _42355_);
  and (_01213_, _40957_, _40954_);
  or (_40958_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_40959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _40806_);
  or (_40960_, _40959_, _40941_);
  and (_40961_, _40960_, _42355_);
  and (_01215_, _40961_, _40958_);
  or (_40962_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_40963_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _40806_);
  or (_40964_, _40963_, _40941_);
  and (_40965_, _40964_, _42355_);
  and (_01217_, _40965_, _40962_);
  or (_40966_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_40967_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _40806_);
  or (_40968_, _40967_, _40941_);
  and (_40969_, _40968_, _42355_);
  and (_01219_, _40969_, _40966_);
  or (_40970_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_40971_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _40806_);
  or (_40972_, _40971_, _40941_);
  and (_40973_, _40972_, _42355_);
  and (_01221_, _40973_, _40970_);
  or (_40974_, _40945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_40975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _40806_);
  or (_40976_, _40975_, _40941_);
  and (_40977_, _40976_, _42355_);
  and (_01223_, _40977_, _40974_);
  nor (_40978_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_40979_, _40978_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_40980_, _40790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_40981_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_40982_, _40981_, _40780_);
  and (_40983_, _40982_, _40980_);
  or (_40984_, _40771_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_40985_, _40984_, _40835_);
  and (_40986_, _40985_, _40803_);
  or (_40987_, _40986_, _40983_);
  or (_40988_, _40987_, _40798_);
  or (_40989_, _40799_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_40990_, _40989_, _40778_);
  and (_40991_, _40990_, _40988_);
  or (_01225_, _40991_, _40979_);
  and (_40992_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_40993_, _40992_, _40836_);
  or (_40994_, _40993_, _40944_);
  and (_40995_, _40994_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_40996_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _40806_);
  nand (_40997_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_40998_, _40997_, _40941_);
  or (_40999_, _40998_, _40996_);
  or (_41000_, _40999_, _40995_);
  and (_01227_, _41000_, _42355_);
  not (_41001_, _40945_);
  and (_41002_, _41001_, _40829_);
  or (_41003_, _40993_, _40942_);
  and (_41004_, _40778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_41005_, _41004_, _41003_);
  or (_01229_, _41005_, _41002_);
  or (_41006_, _40822_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_41007_, _40822_, _40766_);
  and (_41008_, _41007_, _42355_);
  and (_01231_, _41008_, _41006_);
  or (_41009_, _40824_, _40787_);
  or (_41010_, _40793_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_41011_, _41010_, _42355_);
  and (_01232_, _41011_, _41009_);
  and (_41012_, _40824_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_41013_, _40813_, _40819_);
  and (_41014_, _41013_, _40793_);
  or (_41015_, _41014_, _41012_);
  and (_01234_, _41015_, _42355_);
  and (_41016_, _40826_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_41017_, _40819_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41018_, _41017_, _40825_);
  or (_41019_, _41018_, _41016_);
  and (_01236_, _41019_, _42355_);
  and (_41020_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _40806_);
  and (_41021_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41022_, _41021_, _41020_);
  and (_01238_, _41022_, _42355_);
  and (_41023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _40806_);
  and (_41024_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41025_, _41024_, _41023_);
  and (_01240_, _41025_, _42355_);
  and (_41026_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _40806_);
  and (_41027_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41028_, _41027_, _41026_);
  and (_01242_, _41028_, _42355_);
  and (_41029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _40806_);
  and (_41030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41031_, _41030_, _41029_);
  and (_01244_, _41031_, _42355_);
  and (_41032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _40806_);
  and (_41033_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41034_, _41033_, _41032_);
  and (_01246_, _41034_, _42355_);
  and (_41035_, _40778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01248_, _41035_, _40979_);
  and (_41036_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_41037_, _41036_, _40996_);
  and (_01250_, _41037_, _42355_);
  nor (_41038_, _40881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_41039_, _41038_, _40917_);
  and (_01252_, _41039_, _40900_);
  nor (_41040_, _40917_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_41041_, _41040_, _40918_);
  and (_01254_, _41041_, _40900_);
  nor (_41042_, _40918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_41043_, _41042_, _40919_);
  and (_01256_, _41043_, _40900_);
  or (_41044_, _40882_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41045_, _40883_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41046_, _41045_, _41044_);
  and (_41047_, _41046_, _40891_);
  and (_41048_, _40875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_41049_, _41048_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_41050_, _41049_, _40864_);
  or (_41051_, _41050_, _41047_);
  and (_41052_, _41051_, _40900_);
  nor (_41053_, _40769_, _37941_);
  and (_41054_, _41053_, _40903_);
  or (_01258_, _41054_, _41052_);
  not (_41055_, _40924_);
  and (_41056_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_41057_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_41058_, _41057_, _41056_);
  and (_41059_, _41058_, _40900_);
  nand (_41060_, _40768_, _37934_);
  nand (_41061_, _40769_, _37941_);
  and (_41063_, _41061_, _40903_);
  and (_41065_, _41063_, _41060_);
  or (_01260_, _41065_, _41059_);
  nor (_41068_, _40924_, _40870_);
  and (_41070_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_41072_, _41070_, _41068_);
  and (_41074_, _41072_, _40900_);
  nand (_41076_, _40768_, _37927_);
  nand (_41078_, _40769_, _37934_);
  and (_41080_, _41078_, _40903_);
  and (_41082_, _41080_, _41076_);
  or (_01262_, _41082_, _41074_);
  nor (_41085_, _40924_, _40866_);
  and (_41087_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_41089_, _41087_, _41085_);
  and (_41091_, _41089_, _40900_);
  nand (_41093_, _40769_, _37927_);
  nand (_41095_, _40768_, _37920_);
  and (_41097_, _41095_, _40903_);
  and (_41099_, _41097_, _41093_);
  or (_01264_, _41099_, _41091_);
  and (_41102_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_41104_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or (_41106_, _41104_, _41102_);
  and (_41108_, _41106_, _40900_);
  nand (_41110_, _40768_, _37912_);
  nand (_41112_, _40769_, _37920_);
  and (_41114_, _41112_, _40903_);
  and (_41116_, _41114_, _41110_);
  or (_01266_, _41116_, _41108_);
  and (_41119_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_41121_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_41123_, _41121_, _41119_);
  and (_41125_, _41123_, _40900_);
  nand (_41127_, _40769_, _37912_);
  nand (_41128_, _40768_, _37904_);
  and (_41129_, _41128_, _40903_);
  and (_41130_, _41129_, _41127_);
  or (_01267_, _41130_, _41125_);
  and (_41131_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_41132_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_41133_, _41132_, _41131_);
  and (_41134_, _41133_, _40900_);
  nand (_41135_, _40768_, _37896_);
  nand (_41136_, _40769_, _37904_);
  and (_41137_, _41136_, _40903_);
  and (_41138_, _41137_, _41135_);
  or (_01269_, _41138_, _41134_);
  and (_41139_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41140_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_41141_, _41140_, _41139_);
  and (_41142_, _41141_, _40900_);
  nand (_41143_, _40768_, _37963_);
  nand (_41144_, _40769_, _37896_);
  and (_41145_, _41144_, _40903_);
  and (_41146_, _41145_, _41143_);
  or (_01271_, _41146_, _41142_);
  and (_41147_, _40899_, _40769_);
  nand (_41148_, _41147_, _37963_);
  and (_41149_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_41150_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41151_, _41150_, _41149_);
  or (_41152_, _41151_, _40899_);
  and (_41153_, _41152_, _42355_);
  and (_01273_, _41153_, _41148_);
  and (_41154_, _41055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_41155_, _40924_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_41156_, _41155_, _41154_);
  and (_41157_, _41156_, _40900_);
  or (_41158_, _40756_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41159_, _41158_, _40769_);
  and (_41160_, _41159_, _40903_);
  or (_01275_, _41160_, _41157_);
  nand (_41161_, _40927_, _37941_);
  or (_41162_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_41163_, _41162_, _42355_);
  and (_01277_, _41163_, _41161_);
  or (_41164_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_41165_, _41164_, _42355_);
  nand (_41166_, _40927_, _37934_);
  and (_01279_, _41166_, _41165_);
  or (_41167_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_41168_, _41167_, _42355_);
  nand (_41169_, _40927_, _37927_);
  and (_01281_, _41169_, _41168_);
  or (_41170_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_41171_, _41170_, _42355_);
  nand (_41172_, _40927_, _37920_);
  and (_01283_, _41172_, _41171_);
  or (_41173_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_41174_, _41173_, _42355_);
  nand (_41175_, _40927_, _37912_);
  and (_01285_, _41175_, _41174_);
  or (_41176_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_41177_, _41176_, _42355_);
  nand (_41178_, _40927_, _37904_);
  and (_01287_, _41178_, _41177_);
  or (_41179_, _40927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_41180_, _41179_, _42355_);
  nand (_41181_, _40927_, _37896_);
  and (_01289_, _41181_, _41180_);
  not (_41182_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_41183_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41182_);
  or (_41184_, _41183_, _40768_);
  nor (_41185_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_41186_, _41185_, _41184_);
  or (_41187_, _41186_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_41188_, _41187_, _40931_);
  or (_41189_, _27633_, _40773_);
  nand (_41190_, _41189_, _40931_);
  or (_41191_, _41190_, _38560_);
  and (_41192_, _41191_, _41188_);
  or (_41193_, _41192_, _40934_);
  nand (_41194_, _40934_, _37941_);
  and (_41195_, _41194_, _42355_);
  and (_01291_, _41195_, _41193_);
  or (_41196_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_41197_, _41196_, _40931_);
  not (_41198_, _33228_);
  nor (_41199_, _41198_, _31889_);
  nand (_41200_, _41198_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_41201_, _41200_, _40931_);
  or (_41202_, _41201_, _41199_);
  and (_41203_, _41202_, _41197_);
  or (_41204_, _41203_, _40934_);
  nand (_41205_, _40934_, _37934_);
  and (_41206_, _41205_, _42355_);
  and (_01293_, _41206_, _41204_);
  not (_41207_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not (_41208_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_41209_, _40782_, _41208_);
  nor (_41210_, _41209_, _41207_);
  and (_41211_, _41209_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_41212_, _41211_, _41210_);
  or (_41213_, _41212_, _40931_);
  or (_41214_, _33979_, _41207_);
  nand (_41215_, _41214_, _40931_);
  or (_41216_, _41215_, _34001_);
  and (_41217_, _41216_, _41213_);
  or (_41218_, _41217_, _40934_);
  nand (_41219_, _40934_, _37927_);
  and (_41220_, _41219_, _42355_);
  and (_01295_, _41220_, _41218_);
  and (_41221_, _40931_, _34653_);
  nand (_41222_, _41221_, _31889_);
  or (_41223_, _41221_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_41224_, _41223_, _40935_);
  and (_41225_, _41224_, _41222_);
  nor (_41226_, _40935_, _37920_);
  or (_41227_, _41226_, _41225_);
  and (_01297_, _41227_, _42355_);
  and (_41228_, _40931_, _35317_);
  nand (_41229_, _41228_, _31889_);
  or (_41230_, _41228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_41231_, _41230_, _40935_);
  and (_41232_, _41231_, _41229_);
  nor (_41233_, _40935_, _37912_);
  or (_41234_, _41233_, _41232_);
  and (_01299_, _41234_, _42355_);
  and (_41235_, _40931_, _36112_);
  nand (_41236_, _41235_, _31889_);
  or (_41237_, _41235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_41238_, _41237_, _40935_);
  and (_41239_, _41238_, _41236_);
  nor (_41240_, _40935_, _37904_);
  or (_41241_, _41240_, _41239_);
  and (_01301_, _41241_, _42355_);
  and (_41242_, _40931_, _36851_);
  nand (_41243_, _41242_, _31889_);
  or (_41244_, _41242_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_41245_, _41244_, _40935_);
  and (_41246_, _41245_, _41243_);
  nor (_41247_, _40935_, _37896_);
  or (_41248_, _41247_, _41246_);
  and (_01302_, _41248_, _42355_);
  and (_01629_, t2_i, _42355_);
  nor (_41249_, t2_i, rst);
  and (_01632_, _41249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_41250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _42355_);
  nor (_01635_, _41250_, t2ex_i);
  and (_01638_, t2ex_i, _42355_);
  and (_41251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_41252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_41253_, _41252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41254_, _41253_, _41251_);
  not (_41255_, _41254_);
  and (_41256_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41257_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_41258_, _41257_, _41256_);
  and (_41259_, _37879_, _38362_);
  and (_41260_, _41259_, _39479_);
  nor (_41261_, _41260_, _41258_);
  and (_41262_, _27611_, _33957_);
  and (_41263_, _39550_, _41262_);
  and (_41264_, _41259_, _41263_);
  and (_41265_, _41264_, _31301_);
  not (_41266_, _41265_);
  nor (_41267_, _41266_, _37963_);
  or (_41268_, _41267_, _41261_);
  and (_41269_, _41259_, _39285_);
  not (_41270_, _41269_);
  and (_41271_, _41270_, _41268_);
  and (_41272_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_41273_, _41272_, _41271_);
  and (_01641_, _41273_, _42355_);
  nand (_41274_, _41269_, _37963_);
  nor (_41275_, _41260_, _41255_);
  or (_41276_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_41277_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_41278_, _41275_, _41277_);
  and (_41279_, _41278_, _41276_);
  or (_41280_, _41279_, _41269_);
  and (_41281_, _41280_, _42355_);
  and (_01644_, _41281_, _41274_);
  not (_41282_, _41252_);
  or (_41283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_41284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_41285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _41284_);
  and (_41286_, _41285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_41287_, _41286_, _41283_);
  and (_41288_, _41287_, _41282_);
  and (_41289_, _41259_, _39439_);
  and (_41290_, _39284_, _36112_);
  and (_41291_, _41290_, _41259_);
  nor (_41292_, _41291_, _41289_);
  and (_41293_, _41292_, _41288_);
  or (_41294_, _41293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_41295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41296_, _41295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_41297_, _41296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_41298_, _41297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_41299_, _41298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_41300_, _41299_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_41301_, _41300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41302_, _41301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41303_, _41302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_41304_, _41303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_41305_, _41304_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_41306_, _41305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_41307_, _41306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_41308_, _41307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_41309_, _41308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_41310_, _41309_);
  nand (_41311_, _41310_, _41293_);
  and (_41312_, _41311_, _42355_);
  and (_01647_, _41312_, _41294_);
  nand (_41313_, _41289_, _37963_);
  and (_41314_, _41259_, _36112_);
  and (_41315_, _41314_, _39284_);
  not (_41316_, _41315_);
  not (_41317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41318_, _41251_, _41317_);
  and (_41319_, _41318_, _41252_);
  and (_41320_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not (_41321_, _41319_);
  and (_41322_, _41300_, _41287_);
  or (_41323_, _41322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_41324_, _41322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_41325_, _41324_, _41323_);
  not (_41326_, _41253_);
  and (_41327_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_41328_, _41309_, _41287_);
  and (_41329_, _41328_, _41327_);
  or (_41330_, _41329_, _41325_);
  and (_41331_, _41330_, _41321_);
  or (_41332_, _41331_, _41320_);
  or (_41333_, _41332_, _41289_);
  and (_41334_, _41333_, _41316_);
  and (_41335_, _41334_, _41313_);
  and (_41336_, _41315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_41337_, _41336_, _41335_);
  and (_01650_, _41337_, _42355_);
  nand (_41338_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_41339_, _41338_, _41287_);
  nand (_41340_, _41339_, _41309_);
  and (_41341_, _41308_, _41287_);
  or (_41342_, _41341_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_41343_, _41342_, _41321_);
  and (_41344_, _41343_, _41340_);
  nand (_41345_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_41346_, _41345_, _41292_);
  or (_41347_, _41346_, _41344_);
  nand (_41348_, _41289_, _41277_);
  and (_41349_, _41348_, _42355_);
  and (_41350_, _41349_, _41347_);
  nand (_41351_, _41315_, _37963_);
  and (_01653_, _41351_, _41350_);
  and (_41352_, _41287_, _41252_);
  and (_41353_, _41352_, _41321_);
  nand (_41354_, _41353_, _41309_);
  nand (_41355_, _41354_, _41292_);
  or (_41356_, _41292_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41357_, _41356_, _42355_);
  and (_01656_, _41357_, _41355_);
  or (_41358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41359_, _40038_, _38346_);
  or (_41360_, _41359_, _41358_);
  nand (_41361_, _38349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_41362_, _41361_, _41359_);
  or (_41363_, _41362_, _38350_);
  and (_41364_, _41363_, _41360_);
  and (_41365_, _41259_, _40034_);
  or (_41366_, _41365_, _41364_);
  nand (_41367_, _41365_, _37963_);
  and (_41368_, _41367_, _42355_);
  and (_01659_, _41368_, _41366_);
  not (_41369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_41370_, _41254_, _41369_);
  and (_41371_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_41372_, _41371_, _41370_);
  or (_41373_, _41372_, _41260_);
  nand (_41374_, _41260_, _37941_);
  and (_41375_, _41374_, _41373_);
  or (_41376_, _41375_, _41269_);
  nand (_41377_, _41269_, _41369_);
  and (_41378_, _41377_, _42355_);
  and (_02110_, _41378_, _41376_);
  nand (_41379_, _41260_, _37934_);
  and (_41380_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41381_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_41382_, _41381_, _41380_);
  or (_41383_, _41382_, _41260_);
  and (_41384_, _41383_, _41379_);
  or (_41385_, _41384_, _41269_);
  or (_41386_, _41270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41387_, _41386_, _42355_);
  and (_02112_, _41387_, _41385_);
  and (_41388_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41389_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_41390_, _41389_, _41388_);
  nor (_41391_, _41390_, _41260_);
  nor (_41392_, _41266_, _37927_);
  or (_41393_, _41392_, _41391_);
  and (_41394_, _41393_, _41270_);
  and (_41395_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_41396_, _41395_, _41394_);
  and (_02113_, _41396_, _42355_);
  and (_41397_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41398_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_41399_, _41398_, _41397_);
  nor (_41400_, _41399_, _41260_);
  nor (_41401_, _41266_, _37920_);
  or (_41402_, _41401_, _41400_);
  and (_41403_, _41402_, _41270_);
  and (_41404_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_41405_, _41404_, _41403_);
  and (_02115_, _41405_, _42355_);
  and (_41406_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_41407_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_41408_, _41407_, _41406_);
  nor (_41409_, _41408_, _41260_);
  nor (_41410_, _41266_, _37912_);
  or (_41411_, _41410_, _41409_);
  and (_41412_, _41411_, _41270_);
  and (_41413_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_41414_, _41413_, _41412_);
  and (_02117_, _41414_, _42355_);
  and (_41415_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41416_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_41417_, _41416_, _41415_);
  nor (_41418_, _41417_, _41260_);
  nor (_41419_, _41266_, _37904_);
  or (_41420_, _41419_, _41418_);
  and (_41421_, _41420_, _41270_);
  and (_41422_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_41423_, _41422_, _41421_);
  and (_02119_, _41423_, _42355_);
  and (_41424_, _41255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41425_, _41254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_41426_, _41425_, _41424_);
  nor (_41427_, _41426_, _41260_);
  nor (_41428_, _41266_, _37896_);
  or (_41429_, _41428_, _41427_);
  and (_41430_, _41429_, _41270_);
  and (_41431_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_41432_, _41431_, _41430_);
  and (_02120_, _41432_, _42355_);
  or (_41433_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_41434_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_41435_, _41275_, _41434_);
  and (_41436_, _41435_, _41433_);
  or (_41437_, _41436_, _41269_);
  nand (_41438_, _41269_, _37941_);
  and (_41439_, _41438_, _42355_);
  and (_02122_, _41439_, _41437_);
  and (_41440_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  not (_41441_, _41275_);
  and (_41442_, _41441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_41443_, _41442_, _41440_);
  and (_41444_, _41443_, _41270_);
  nor (_41445_, _41270_, _37934_);
  or (_41446_, _41445_, _41444_);
  and (_02124_, _41446_, _42355_);
  nand (_41447_, _41269_, _37927_);
  and (_41448_, _41441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41449_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_41450_, _41449_, _41448_);
  or (_41451_, _41450_, _41269_);
  and (_41452_, _41451_, _42355_);
  and (_02126_, _41452_, _41447_);
  nand (_41453_, _41269_, _37920_);
  and (_41454_, _41441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41455_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41456_, _41455_, _41454_);
  or (_41457_, _41456_, _41269_);
  and (_41458_, _41457_, _42355_);
  and (_02127_, _41458_, _41453_);
  nand (_41459_, _41269_, _37912_);
  and (_41460_, _41441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_41461_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41462_, _41461_, _41460_);
  or (_41463_, _41462_, _41269_);
  and (_41464_, _41463_, _42355_);
  and (_02129_, _41464_, _41459_);
  nand (_41465_, _41269_, _37904_);
  and (_41466_, _41441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41467_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41468_, _41467_, _41466_);
  or (_41469_, _41468_, _41269_);
  and (_41470_, _41469_, _42355_);
  and (_02131_, _41470_, _41465_);
  nand (_41471_, _41269_, _37896_);
  and (_41472_, _41441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41473_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_41474_, _41473_, _41472_);
  or (_41475_, _41474_, _41269_);
  and (_41476_, _41475_, _42355_);
  and (_02133_, _41476_, _41471_);
  and (_41477_, _41287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_41478_, _41253_, _41369_);
  nand (_41479_, _41478_, _41309_);
  nand (_41480_, _41479_, _41477_);
  or (_41481_, _41287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_41482_, _41481_, _41321_);
  and (_41483_, _41482_, _41480_);
  and (_41484_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_41485_, _41484_, _41289_);
  or (_41486_, _41485_, _41483_);
  and (_41487_, _41289_, _37941_);
  nor (_41488_, _41487_, _41315_);
  and (_41489_, _41488_, _41486_);
  and (_41490_, _41315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_41491_, _41490_, _41489_);
  and (_02134_, _41491_, _42355_);
  and (_41492_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_41493_, _41492_, _41287_);
  and (_41494_, _41493_, _41309_);
  or (_41495_, _41477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_41496_, _41295_, _41287_);
  and (_41497_, _41496_, _41495_);
  or (_41498_, _41497_, _41494_);
  and (_41499_, _41498_, _41321_);
  and (_41500_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_41501_, _41500_, _41289_);
  or (_41502_, _41501_, _41499_);
  nand (_41503_, _41289_, _37934_);
  and (_41504_, _41503_, _41316_);
  and (_41505_, _41504_, _41502_);
  and (_41506_, _41315_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_41507_, _41506_, _41505_);
  and (_02136_, _41507_, _42355_);
  not (_41508_, _41289_);
  nor (_41509_, _41508_, _37927_);
  and (_41510_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41511_, _41510_, _41328_);
  and (_41512_, _41496_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_41513_, _41496_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_41514_, _41513_, _41319_);
  or (_41515_, _41514_, _41512_);
  or (_41516_, _41515_, _41511_);
  or (_41517_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_41518_, _41517_, _41292_);
  and (_41519_, _41518_, _41516_);
  and (_41520_, _41291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_41521_, _41520_, _41519_);
  or (_41522_, _41521_, _41509_);
  and (_02138_, _41522_, _42355_);
  nor (_41523_, _41508_, _37920_);
  and (_41524_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41525_, _41524_, _41328_);
  nand (_41526_, _41296_, _41287_);
  and (_41527_, _41526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_41528_, _41526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_41529_, _41528_, _41319_);
  or (_41530_, _41529_, _41527_);
  or (_41531_, _41530_, _41525_);
  or (_41532_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_41533_, _41532_, _41292_);
  and (_41534_, _41533_, _41531_);
  and (_41535_, _41291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_41536_, _41535_, _41534_);
  or (_41537_, _41536_, _41523_);
  and (_02140_, _41537_, _42355_);
  nor (_41538_, _41508_, _37912_);
  and (_41539_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_41540_, _41539_, _41328_);
  nand (_41541_, _41297_, _41287_);
  and (_41542_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_41543_, _41541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_41544_, _41543_, _41319_);
  or (_41545_, _41544_, _41542_);
  or (_41546_, _41545_, _41540_);
  or (_41547_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_41548_, _41547_, _41292_);
  and (_41549_, _41548_, _41546_);
  and (_41550_, _41291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_41551_, _41550_, _41549_);
  or (_41552_, _41551_, _41538_);
  and (_02141_, _41552_, _42355_);
  nor (_41553_, _41508_, _37904_);
  and (_41554_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41555_, _41554_, _41328_);
  nand (_41556_, _41298_, _41287_);
  and (_41557_, _41556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_41558_, _41556_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_41559_, _41558_, _41319_);
  or (_41560_, _41559_, _41557_);
  or (_41561_, _41560_, _41555_);
  or (_41562_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_41563_, _41562_, _41292_);
  and (_41564_, _41563_, _41561_);
  and (_41565_, _41291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_41566_, _41565_, _41564_);
  or (_41567_, _41566_, _41553_);
  and (_02143_, _41567_, _42355_);
  nor (_41568_, _41508_, _37896_);
  and (_41569_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41570_, _41569_, _41328_);
  and (_41571_, _41299_, _41287_);
  nor (_41572_, _41571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_41573_, _41572_, _41322_);
  or (_41574_, _41573_, _41319_);
  or (_41575_, _41574_, _41570_);
  or (_41576_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_41577_, _41576_, _41292_);
  and (_41578_, _41577_, _41575_);
  and (_41579_, _41291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_41580_, _41579_, _41578_);
  or (_41581_, _41580_, _41568_);
  and (_02145_, _41581_, _42355_);
  not (_41582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_41583_, _41253_, _41582_);
  and (_41584_, _41583_, _41328_);
  and (_41585_, _41301_, _41287_);
  or (_41586_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_41587_, _41585_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41588_, _41587_, _41586_);
  or (_41589_, _41588_, _41319_);
  or (_41590_, _41589_, _41584_);
  nand (_41591_, _41319_, _41582_);
  and (_41592_, _41591_, _41292_);
  and (_41593_, _41592_, _41590_);
  and (_41594_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_41595_, _41315_, _37942_);
  or (_41596_, _41595_, _41594_);
  or (_41597_, _41596_, _41593_);
  and (_02147_, _41597_, _42355_);
  and (_41598_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_41599_, _41598_, _41328_);
  and (_41600_, _41302_, _41287_);
  or (_41601_, _41600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_41602_, _41600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_41603_, _41602_, _41601_);
  or (_41604_, _41603_, _41319_);
  or (_41605_, _41604_, _41599_);
  or (_41606_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_41607_, _41606_, _41292_);
  and (_41608_, _41607_, _41605_);
  and (_41609_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_41610_, _41316_, _37934_);
  or (_41611_, _41610_, _41609_);
  or (_41612_, _41611_, _41608_);
  and (_02148_, _41612_, _42355_);
  and (_41613_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41614_, _41613_, _41328_);
  and (_41615_, _41303_, _41287_);
  or (_41616_, _41615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand (_41617_, _41615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_41618_, _41617_, _41616_);
  or (_41619_, _41618_, _41319_);
  or (_41620_, _41619_, _41614_);
  or (_41621_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_41622_, _41621_, _41292_);
  and (_41623_, _41622_, _41620_);
  and (_41624_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_41625_, _41316_, _37927_);
  or (_41626_, _41625_, _41624_);
  or (_41627_, _41626_, _41623_);
  and (_02150_, _41627_, _42355_);
  and (_41628_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41629_, _41628_, _41328_);
  nand (_41630_, _41304_, _41287_);
  nor (_41631_, _41630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_41632_, _41630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41633_, _41632_, _41319_);
  or (_41634_, _41633_, _41631_);
  or (_41635_, _41634_, _41629_);
  or (_41636_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_41637_, _41636_, _41292_);
  and (_41638_, _41637_, _41635_);
  and (_41639_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_41640_, _41639_, _41638_);
  and (_41641_, _41259_, _39289_);
  and (_41642_, _41641_, _31301_);
  and (_41643_, _41642_, _40726_);
  or (_41644_, _41643_, _41640_);
  and (_02152_, _41644_, _42355_);
  and (_41645_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_41646_, _41645_, _41328_);
  nand (_41647_, _41305_, _41287_);
  nor (_41648_, _41647_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_41649_, _41647_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41650_, _41649_, _41319_);
  or (_41651_, _41650_, _41648_);
  or (_41652_, _41651_, _41646_);
  or (_41653_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_41654_, _41653_, _41292_);
  and (_41655_, _41654_, _41652_);
  and (_41656_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_41657_, _41656_, _41655_);
  and (_41658_, _41642_, _40734_);
  or (_41659_, _41658_, _41657_);
  and (_02154_, _41659_, _42355_);
  and (_41660_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41661_, _41660_, _41328_);
  nand (_41662_, _41306_, _41287_);
  and (_41663_, _41662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_41664_, _41662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_41665_, _41664_, _41319_);
  or (_41666_, _41665_, _41663_);
  or (_41667_, _41666_, _41661_);
  or (_41668_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_41669_, _41668_, _41292_);
  and (_41670_, _41669_, _41667_);
  and (_41671_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_41672_, _41316_, _37904_);
  or (_41673_, _41672_, _41671_);
  or (_41674_, _41673_, _41670_);
  and (_02155_, _41674_, _42355_);
  and (_41675_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_41676_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41677_, _41676_, _41328_);
  and (_41678_, _41307_, _41287_);
  nor (_41679_, _41678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_41680_, _41679_, _41341_);
  or (_41681_, _41680_, _41319_);
  or (_41682_, _41681_, _41677_);
  or (_41683_, _41321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_41684_, _41683_, _41292_);
  and (_41685_, _41684_, _41682_);
  or (_41686_, _41685_, _41675_);
  not (_41687_, _37896_);
  and (_41688_, _41642_, _41687_);
  or (_41689_, _41688_, _41686_);
  and (_02156_, _41689_, _42355_);
  not (_41690_, _41365_);
  and (_41691_, _41359_, _27633_);
  or (_41692_, _41691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_41693_, _41692_, _41690_);
  nand (_41694_, _41691_, _31889_);
  and (_41695_, _41694_, _41693_);
  nor (_41696_, _41690_, _37941_);
  or (_41697_, _41696_, _41695_);
  and (_02157_, _41697_, _42355_);
  and (_41698_, _41359_, _33228_);
  or (_41699_, _41698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_41700_, _41699_, _41690_);
  nand (_41701_, _41698_, _31889_);
  and (_41702_, _41701_, _41700_);
  nor (_41703_, _41690_, _37934_);
  or (_41704_, _41703_, _41702_);
  and (_02158_, _41704_, _42355_);
  nand (_41705_, _41359_, _38759_);
  and (_41706_, _41705_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_41707_, _41706_, _41365_);
  and (_41708_, _34012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_41709_, _41708_, _34001_);
  and (_41710_, _41709_, _41359_);
  or (_41711_, _41710_, _41707_);
  nand (_41712_, _41365_, _37927_);
  and (_41713_, _41712_, _42355_);
  and (_02159_, _41713_, _41711_);
  and (_41714_, _41359_, _34653_);
  or (_41715_, _41714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_41716_, _41715_, _41690_);
  nand (_41717_, _41714_, _31889_);
  and (_41718_, _41717_, _41716_);
  nor (_41719_, _41690_, _37920_);
  or (_41720_, _41719_, _41718_);
  and (_02160_, _41720_, _42355_);
  and (_41721_, _41359_, _35317_);
  or (_41722_, _41721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_41723_, _41722_, _41690_);
  nand (_41724_, _41721_, _31889_);
  and (_41725_, _41724_, _41723_);
  nor (_41726_, _41690_, _37912_);
  or (_41727_, _41726_, _41725_);
  and (_02161_, _41727_, _42355_);
  and (_41728_, _41359_, _36112_);
  or (_41729_, _41728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_41730_, _41729_, _41690_);
  nand (_41731_, _41728_, _31889_);
  and (_41732_, _41731_, _41730_);
  nor (_41733_, _41690_, _37904_);
  or (_41734_, _41733_, _41732_);
  and (_02162_, _41734_, _42355_);
  not (_41735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_41736_, _41251_, _41735_);
  or (_41737_, _41736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_41738_, _41737_, _41359_);
  nand (_41739_, _38466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_41740_, _41739_, _41359_);
  or (_41741_, _41740_, _38467_);
  and (_41742_, _41741_, _41738_);
  or (_41743_, _41742_, _41365_);
  nand (_41744_, _41365_, _37896_);
  and (_41745_, _41744_, _42355_);
  and (_02163_, _41745_, _41743_);
  and (_41746_, _31278_, _28115_);
  and (_41747_, _37965_, _37875_);
  not (_41748_, _41747_);
  not (_41749_, _37874_);
  nor (_41750_, _41749_, _37839_);
  not (_41751_, _37025_);
  and (_41752_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_41753_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_41754_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_41755_, _41754_, _41753_);
  and (_41756_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_41757_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_41758_, _41757_, _41756_);
  and (_41759_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_41760_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_41761_, _41760_, _41759_);
  and (_41762_, _41761_, _41758_);
  and (_41763_, _41762_, _41755_);
  nor (_41764_, _37156_, _41751_);
  not (_41765_, _41764_);
  nor (_41766_, _41765_, _41763_);
  nor (_41767_, _41766_, _41752_);
  not (_41768_, _41767_);
  and (_41769_, _41768_, _41750_);
  not (_41770_, _41769_);
  not (_41771_, _37740_);
  and (_41772_, _41749_, _37839_);
  and (_41773_, _38450_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_41774_, _41773_, _38446_);
  nor (_41775_, _41774_, _37750_);
  and (_41776_, _41775_, _38453_);
  and (_41777_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_41778_, _41774_, _37633_);
  and (_41779_, _41778_, _38453_);
  and (_41780_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_41781_, _41780_, _41777_);
  not (_41782_, _38453_);
  and (_41783_, _41775_, _41782_);
  and (_41784_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_41785_, _41774_, _37750_);
  and (_41786_, _41785_, _41782_);
  and (_41787_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_41788_, _41787_, _41784_);
  and (_41789_, _41788_, _41781_);
  not (_41790_, _28433_);
  nor (_41791_, _38453_, _41790_);
  and (_41792_, _38453_, _41790_);
  nor (_41793_, _41792_, _41791_);
  and (_41794_, _37633_, _27611_);
  nor (_41795_, _37633_, _27611_);
  nor (_41796_, _41795_, _41794_);
  and (_41797_, _27830_, _28137_);
  not (_41798_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_41799_, _31278_, _41798_);
  and (_41800_, _41799_, _34012_);
  and (_41801_, _41800_, _41797_);
  and (_41802_, _41801_, _41796_);
  and (_41803_, _41802_, _27961_);
  and (_41804_, _41774_, _28301_);
  nor (_41805_, _41774_, _28301_);
  nor (_41806_, _41805_, _41804_);
  and (_41807_, _41806_, _41803_);
  and (_41808_, _41807_, _41793_);
  not (_41809_, _41808_);
  and (_41810_, _41778_, _41782_);
  and (_41811_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_41812_, _41774_, _37633_);
  and (_41813_, _41812_, _38453_);
  and (_41814_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_41815_, _41814_, _41811_);
  and (_41816_, _41812_, _41782_);
  and (_41817_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_41818_, _41785_, _38453_);
  and (_41819_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_41820_, _41819_, _41817_);
  and (_41821_, _41820_, _41815_);
  and (_41822_, _41821_, _41809_);
  and (_41823_, _41822_, _41789_);
  and (_41824_, _41808_, _37963_);
  nor (_41825_, _41824_, _41823_);
  and (_41826_, _41825_, _41772_);
  nor (_41827_, _41826_, _41771_);
  and (_41828_, _41827_, _41770_);
  and (_41829_, _41828_, _41748_);
  not (_41830_, _37778_);
  and (_41831_, _41830_, _37758_);
  and (_41832_, _37610_, _37724_);
  nor (_41833_, _41832_, _37768_);
  and (_41834_, _37724_, _37752_);
  nor (_41835_, _41834_, _37774_);
  and (_41836_, _41835_, _41833_);
  and (_41837_, _37826_, _37790_);
  and (_41838_, _41837_, _41836_);
  and (_41839_, _41838_, _41831_);
  nor (_41840_, _41839_, _36982_);
  nor (_41841_, _37788_, _37784_);
  not (_41842_, _37722_);
  nor (_41843_, _41842_, _41841_);
  nor (_41844_, _41843_, _41840_);
  not (_41845_, _41844_);
  and (_41846_, _41845_, _41829_);
  and (_41847_, _37740_, _37874_);
  and (_41848_, _41847_, _37839_);
  and (_41849_, _41848_, _41782_);
  and (_41850_, _41750_, _37740_);
  and (_41851_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_41852_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_41853_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_41854_, _41853_, _41852_);
  and (_41855_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_41856_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_41857_, _41856_, _41855_);
  and (_41858_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_41859_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_41860_, _41859_, _41858_);
  and (_41861_, _41860_, _41857_);
  and (_41862_, _41861_, _41854_);
  nor (_41863_, _41862_, _41765_);
  nor (_41864_, _41863_, _41851_);
  not (_41865_, _41864_);
  and (_41866_, _41865_, _41850_);
  nor (_41867_, _41866_, _41849_);
  and (_41868_, _41772_, _37740_);
  and (_41869_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_41870_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_41871_, _41870_, _41869_);
  and (_41872_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_41873_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_41874_, _41873_, _41872_);
  and (_41875_, _41874_, _41871_);
  and (_41876_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_41877_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_41878_, _41877_, _41876_);
  and (_41879_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_41880_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_41881_, _41880_, _41879_);
  and (_41882_, _41881_, _41878_);
  and (_41883_, _41882_, _41809_);
  and (_41884_, _41883_, _41875_);
  and (_41885_, _41808_, _37912_);
  nor (_41886_, _41885_, _41884_);
  and (_41887_, _41886_, _41868_);
  not (_41888_, _41887_);
  not (_41889_, _37997_);
  and (_41890_, _41889_, _37876_);
  and (_41891_, _41771_, _37874_);
  nor (_41892_, _41891_, _41890_);
  and (_41893_, _41892_, _41888_);
  and (_41894_, _41893_, _41867_);
  not (_41895_, _41894_);
  and (_41896_, _41895_, _41846_);
  and (_41897_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_41898_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_41899_, _41898_, _41897_);
  and (_41900_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_41901_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_41902_, _41901_, _41900_);
  and (_41903_, _41902_, _41899_);
  and (_41904_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_41905_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_41906_, _41905_, _41904_);
  and (_41907_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_41908_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_41909_, _41908_, _41907_);
  and (_41910_, _41909_, _41906_);
  and (_41911_, _41910_, _41809_);
  and (_41912_, _41911_, _41903_);
  and (_41913_, _41808_, _37934_);
  nor (_41914_, _41913_, _41912_);
  and (_41915_, _41914_, _41868_);
  and (_41916_, _41772_, _41771_);
  not (_41917_, _37979_);
  and (_41918_, _41917_, _37876_);
  or (_41919_, _41918_, _41916_);
  and (_41920_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_41921_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_41922_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_41923_, _41922_, _41921_);
  and (_41924_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_41925_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_41926_, _41925_, _41924_);
  and (_41927_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_41928_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_41929_, _41928_, _41927_);
  and (_41930_, _41929_, _41926_);
  and (_41931_, _41930_, _41923_);
  nor (_41932_, _41931_, _41765_);
  nor (_41933_, _41932_, _41920_);
  not (_41934_, _41933_);
  and (_41935_, _41934_, _41850_);
  and (_41936_, _41848_, _37657_);
  or (_41937_, _41936_, _41935_);
  or (_41938_, _41937_, _41919_);
  nor (_41939_, _41938_, _41915_);
  nor (_41940_, _41939_, _41845_);
  nor (_41941_, _41940_, _41896_);
  and (_41942_, _28137_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_41943_, _41942_, _41790_);
  nor (_41944_, _27490_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_41945_, _41944_, _41943_);
  nand (_41946_, _41945_, _41941_);
  or (_41947_, _41945_, _41941_);
  and (_41948_, _41947_, _41946_);
  and (_41949_, _41942_, _28301_);
  nor (_41950_, _27611_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_41951_, _41950_, _41949_);
  not (_41952_, _41951_);
  not (_41953_, _41774_);
  and (_41954_, _41848_, _41953_);
  and (_41955_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_41956_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_41957_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_41958_, _41957_, _41956_);
  and (_41959_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_41960_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_41961_, _41960_, _41959_);
  and (_41962_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_41963_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_41964_, _41963_, _41962_);
  and (_41965_, _41964_, _41961_);
  and (_41966_, _41965_, _41958_);
  nor (_41967_, _41966_, _41765_);
  nor (_41968_, _41967_, _41955_);
  not (_41969_, _41968_);
  and (_41970_, _41969_, _41850_);
  nor (_41971_, _41970_, _41954_);
  not (_41972_, _37991_);
  and (_41973_, _41972_, _37876_);
  and (_41974_, _41808_, _37920_);
  and (_41975_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_41976_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_41977_, _41976_, _41975_);
  and (_41978_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_41979_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_41980_, _41979_, _41978_);
  and (_41981_, _41980_, _41977_);
  and (_41982_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_41983_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_41984_, _41983_, _41982_);
  and (_41985_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_41986_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_41987_, _41986_, _41985_);
  and (_41988_, _41987_, _41984_);
  and (_41989_, _41988_, _41809_);
  and (_41990_, _41989_, _41981_);
  nor (_41991_, _41990_, _41974_);
  and (_41992_, _41991_, _41868_);
  nor (_41993_, _41992_, _41973_);
  and (_41994_, _41993_, _41971_);
  not (_41995_, _41994_);
  and (_41996_, _41995_, _41846_);
  and (_41997_, _41848_, _37633_);
  and (_41998_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_41999_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_42000_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_42001_, _42000_, _41999_);
  and (_42002_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42003_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_42004_, _42003_, _42002_);
  and (_42005_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_42006_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_42007_, _42006_, _42005_);
  and (_42008_, _42007_, _42004_);
  and (_42009_, _42008_, _42001_);
  nor (_42010_, _42009_, _41765_);
  nor (_42011_, _42010_, _41998_);
  not (_42012_, _42011_);
  and (_42013_, _42012_, _41850_);
  nor (_42014_, _42013_, _41997_);
  not (_42015_, _37973_);
  and (_42016_, _42015_, _37876_);
  and (_42017_, _41808_, _37941_);
  and (_42018_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_42019_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_42020_, _42019_, _42018_);
  and (_42021_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_42022_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_42023_, _42022_, _42021_);
  and (_42024_, _42023_, _42020_);
  and (_42025_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_42026_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_42027_, _42026_, _42025_);
  and (_42028_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_42029_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_42030_, _42029_, _42028_);
  and (_42031_, _42030_, _42027_);
  and (_42032_, _42031_, _41809_);
  and (_42033_, _42032_, _42024_);
  nor (_42034_, _42033_, _42017_);
  and (_42035_, _42034_, _41868_);
  nor (_42036_, _42035_, _42016_);
  and (_42037_, _42036_, _42014_);
  nor (_42038_, _42037_, _41845_);
  nor (_42039_, _42038_, _41996_);
  and (_42040_, _42039_, _41952_);
  nor (_42041_, _42039_, _41952_);
  nor (_42042_, _42041_, _42040_);
  not (_42043_, _42042_);
  nor (_42044_, _42043_, _41948_);
  and (_42045_, _41942_, _37880_);
  nor (_42046_, _41942_, _28290_);
  nor (_42047_, _42046_, _42045_);
  nor (_42048_, _41772_, _37740_);
  and (_42049_, _41808_, _37896_);
  and (_42050_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_42051_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_42052_, _42051_, _42050_);
  and (_42053_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_42054_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_42055_, _42054_, _42053_);
  and (_42056_, _42055_, _42052_);
  and (_42057_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_42058_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_42059_, _42058_, _42057_);
  and (_42060_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_42061_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_42062_, _42061_, _42060_);
  and (_42063_, _42062_, _42059_);
  and (_42064_, _42063_, _41809_);
  and (_42065_, _42064_, _42056_);
  nor (_42066_, _42065_, _42049_);
  and (_42067_, _42066_, _41868_);
  nor (_42068_, _42067_, _42048_);
  not (_42069_, _38009_);
  and (_42070_, _42069_, _37876_);
  and (_42071_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_42072_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42073_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_42074_, _42073_, _42072_);
  and (_42075_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_42076_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_42077_, _42076_, _42075_);
  and (_42078_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_42079_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_42080_, _42079_, _42078_);
  and (_42081_, _42080_, _42077_);
  and (_42082_, _42081_, _42074_);
  nor (_42083_, _42082_, _41765_);
  nor (_42084_, _42083_, _42071_);
  not (_42085_, _42084_);
  and (_42086_, _42085_, _41850_);
  nor (_42087_, _42086_, _42070_);
  and (_42088_, _42087_, _42068_);
  and (_42089_, _42088_, _41846_);
  nor (_42090_, _41995_, _41846_);
  nor (_42091_, _42090_, _42089_);
  nor (_42092_, _42091_, _42047_);
  and (_42093_, _42091_, _42047_);
  nor (_42094_, _42093_, _42092_);
  not (_42095_, _41846_);
  and (_42096_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_42097_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor (_42098_, _42097_, _42096_);
  and (_42099_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_42100_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_42101_, _42100_, _42099_);
  and (_42102_, _42101_, _42098_);
  and (_42103_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_42104_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_42105_, _42104_, _42103_);
  and (_42106_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_42107_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_42108_, _42107_, _42106_);
  and (_42109_, _42108_, _42105_);
  and (_42110_, _42109_, _41809_);
  and (_42111_, _42110_, _42102_);
  and (_42112_, _41808_, _37904_);
  nor (_42113_, _42112_, _42111_);
  and (_42114_, _42113_, _41868_);
  and (_42115_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_42116_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_42117_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_42118_, _42117_, _42116_);
  and (_42119_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42120_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_42121_, _42120_, _42119_);
  and (_42122_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_42123_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_42124_, _42123_, _42122_);
  and (_42125_, _42124_, _42121_);
  and (_42126_, _42125_, _42118_);
  nor (_42127_, _42126_, _41765_);
  nor (_42128_, _42127_, _42115_);
  not (_42129_, _42128_);
  and (_42130_, _42129_, _41850_);
  nor (_42131_, _42130_, _42114_);
  nor (_42132_, _38003_, _37874_);
  nor (_42133_, _42132_, _41771_);
  not (_42134_, _42133_);
  nor (_42135_, _41750_, _41772_);
  and (_42136_, _42135_, _42134_);
  not (_42137_, _42136_);
  and (_42138_, _42137_, _42131_);
  nor (_42139_, _42138_, _42095_);
  and (_42140_, _41848_, _37679_);
  and (_42141_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_42142_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42143_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_42144_, _42143_, _42142_);
  and (_42145_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_42146_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_42147_, _42146_, _42145_);
  and (_42148_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_42149_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_42150_, _42149_, _42148_);
  and (_42151_, _42150_, _42147_);
  and (_42152_, _42151_, _42144_);
  nor (_42153_, _42152_, _41765_);
  nor (_42154_, _42153_, _42141_);
  not (_42155_, _42154_);
  and (_42156_, _42155_, _41850_);
  nor (_42157_, _42156_, _42140_);
  not (_42158_, _37985_);
  and (_42159_, _42158_, _37876_);
  and (_42160_, _41808_, _37927_);
  and (_42161_, _41783_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_42162_, _41810_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_42163_, _42162_, _42161_);
  and (_42164_, _41786_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_42165_, _41813_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_42166_, _42165_, _42164_);
  and (_42167_, _42166_, _42163_);
  and (_42168_, _41776_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_42169_, _41779_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_42170_, _42169_, _42168_);
  and (_42171_, _41816_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_42172_, _41818_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_42173_, _42172_, _42171_);
  and (_42174_, _42173_, _42170_);
  and (_42175_, _42174_, _41809_);
  and (_42176_, _42175_, _42167_);
  nor (_42177_, _42176_, _42160_);
  and (_42178_, _42177_, _41868_);
  nor (_42179_, _42178_, _42159_);
  and (_42180_, _42179_, _42157_);
  nor (_42181_, _42180_, _41845_);
  nor (_42182_, _42181_, _42139_);
  and (_42183_, _41942_, _38345_);
  nor (_42184_, _27369_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_42185_, _42184_, _42183_);
  not (_42186_, _42185_);
  nor (_42187_, _42186_, _42182_);
  and (_42188_, _42186_, _42182_);
  nor (_42189_, _42188_, _42187_);
  and (_42190_, _42189_, _42094_);
  and (_42191_, _42190_, _42044_);
  and (_42192_, _42191_, _41746_);
  nor (_42193_, _42088_, _41846_);
  nor (_42194_, _41942_, _27830_);
  not (_42195_, _42194_);
  nor (_42196_, _42195_, _42193_);
  and (_42197_, _42195_, _42193_);
  nor (_42198_, _42197_, _42196_);
  nor (_42199_, _41894_, _41846_);
  nor (_42200_, _41942_, _28433_);
  not (_42201_, _42200_);
  nor (_42202_, _42201_, _42199_);
  and (_42203_, _42201_, _42199_);
  nor (_42204_, _42203_, _42202_);
  and (_42205_, _42138_, _42095_);
  nor (_42206_, _41942_, _38345_);
  not (_42207_, _42206_);
  nor (_42208_, _42207_, _42205_);
  and (_42209_, _42207_, _42205_);
  nor (_42210_, _41829_, _28137_);
  and (_42211_, _41829_, _28137_);
  nor (_42212_, _42211_, _42210_);
  or (_42213_, _42212_, _42209_);
  nor (_42214_, _42213_, _42208_);
  and (_42215_, _42214_, _42204_);
  and (_42216_, _42215_, _42198_);
  and (_42217_, _42216_, _42192_);
  not (_42218_, _42182_);
  not (_42219_, _42039_);
  and (_42220_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_42221_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_42222_, _42221_, _41941_);
  or (_42223_, _42222_, _42220_);
  and (_42224_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_42225_, _41941_);
  and (_42226_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_42227_, _42226_, _42225_);
  or (_42228_, _42227_, _42224_);
  and (_42229_, _42228_, _42223_);
  or (_42230_, _42229_, _42218_);
  not (_42231_, _42091_);
  and (_42232_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_42233_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_42234_, _42233_, _41941_);
  or (_42235_, _42234_, _42232_);
  and (_42236_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_42237_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_42238_, _42237_, _42225_);
  or (_42239_, _42238_, _42236_);
  and (_42240_, _42239_, _42235_);
  or (_42241_, _42240_, _42182_);
  and (_42242_, _42241_, _42231_);
  and (_42243_, _42242_, _42230_);
  or (_42244_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_42245_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_42246_, _42245_, _42244_);
  or (_42247_, _42246_, _42225_);
  or (_42248_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_42249_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_42250_, _42249_, _42248_);
  or (_42251_, _42250_, _41941_);
  and (_42252_, _42251_, _42247_);
  or (_42253_, _42252_, _42218_);
  or (_42254_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_42255_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_42256_, _42255_, _42254_);
  or (_42257_, _42256_, _42225_);
  or (_42258_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_42259_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_42260_, _42259_, _42258_);
  or (_42261_, _42260_, _41941_);
  and (_42262_, _42261_, _42257_);
  or (_42263_, _42262_, _42182_);
  and (_42264_, _42263_, _42091_);
  and (_42265_, _42264_, _42253_);
  or (_42266_, _42265_, _42243_);
  or (_42267_, _42266_, _42217_);
  not (_42268_, _42217_);
  or (_42269_, _42268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_42270_, _42192_);
  nor (_42271_, _42217_, _42270_);
  nor (_42272_, _42271_, rst);
  and (_42273_, _42272_, _42269_);
  and (_42274_, _42273_, _42267_);
  and (_42275_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_42276_, _42275_, _29233_);
  nor (_42277_, _42276_, _31889_);
  nand (_42278_, _29233_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42279_, _20625_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42280_, _42279_, _42278_);
  nor (_42281_, _37963_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42282_, _42281_, _42280_);
  or (_42283_, _42282_, _42277_);
  and (_39583_, _42283_, _42355_);
  and (_42284_, _39583_, _42271_);
  or (_02567_, _42284_, _42274_);
  not (_42285_, _41746_);
  nor (_42286_, _41951_, _42285_);
  nor (_42287_, _42285_, _41945_);
  and (_42288_, _42287_, _42286_);
  nor (_42289_, _42047_, _42285_);
  nor (_42290_, _42285_, _42185_);
  and (_42291_, _42290_, _42289_);
  and (_42292_, _42291_, _42288_);
  and (_42294_, _42283_, _41746_);
  and (_42295_, _42294_, _42292_);
  not (_42297_, _42292_);
  and (_42299_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_02577_, _42299_, _42295_);
  nor (_42301_, _42290_, _42289_);
  nor (_42303_, _42287_, _42286_);
  and (_42305_, _42303_, _41746_);
  and (_42307_, _42305_, _42301_);
  and (_42308_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _29222_);
  and (_42309_, _42308_, _29266_);
  not (_42310_, _42309_);
  nor (_42311_, _42310_, _31889_);
  not (_42312_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42313_, _37941_, _42312_);
  or (_42314_, _19466_, _42312_);
  and (_42315_, _42314_, _42310_);
  and (_42316_, _42315_, _42313_);
  or (_42317_, _42316_, _42311_);
  and (_42318_, _42317_, _42307_);
  not (_42319_, _42307_);
  and (_42320_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_02801_, _42320_, _42318_);
  nand (_42321_, _42308_, _29310_);
  nor (_42322_, _42321_, _31889_);
  nor (_42323_, _37934_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42324_, _42308_, _29332_);
  and (_42325_, _42308_, _29233_);
  or (_42326_, _42325_, _42275_);
  or (_42327_, _42326_, _42324_);
  and (_42328_, _42327_, _20451_);
  or (_42329_, _42328_, _42323_);
  or (_42330_, _42329_, _42322_);
  and (_42331_, _42330_, _42307_);
  and (_42332_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_02806_, _42332_, _42331_);
  and (_42333_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_42334_, _42308_, _29343_);
  nor (_42335_, _42334_, _31889_);
  nor (_42336_, _37927_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42337_, _42308_, _29299_);
  or (_42338_, _42337_, _42326_);
  and (_42339_, _42338_, _19104_);
  or (_42340_, _42339_, _42336_);
  or (_42341_, _42340_, _42335_);
  and (_42343_, _42341_, _42307_);
  or (_02811_, _42343_, _42333_);
  and (_42346_, _42325_, _32531_);
  nor (_42348_, _37920_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_42350_, _42324_, _42275_);
  or (_42352_, _42350_, _42337_);
  and (_42354_, _42352_, _20136_);
  or (_42356_, _42354_, _42348_);
  or (_42357_, _42356_, _42346_);
  and (_42359_, _42357_, _42307_);
  and (_42361_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_02816_, _42361_, _42359_);
  and (_42362_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_42363_, _42275_, _29266_);
  nor (_42364_, _42363_, _31889_);
  nor (_42365_, _37912_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42366_, _29266_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42367_, _19302_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42368_, _42367_, _42366_);
  or (_42369_, _42368_, _42365_);
  or (_42370_, _42369_, _42364_);
  and (_42371_, _42370_, _42307_);
  or (_02821_, _42371_, _42362_);
  nand (_42372_, _42275_, _29310_);
  nor (_42373_, _42372_, _31889_);
  nor (_42374_, _37904_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42375_, _29310_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42376_, _20288_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42377_, _42376_, _42375_);
  or (_42378_, _42377_, _42374_);
  or (_42379_, _42378_, _42373_);
  and (_42380_, _42379_, _42307_);
  and (_42381_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_02826_, _42381_, _42380_);
  and (_42382_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand (_42383_, _42275_, _29343_);
  nor (_42384_, _42383_, _31889_);
  nor (_42385_, _37896_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_42386_, _29343_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_42387_, _19640_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_42388_, _42387_, _42386_);
  or (_42389_, _42388_, _42385_);
  or (_42390_, _42389_, _42384_);
  and (_42391_, _42390_, _42307_);
  or (_02831_, _42391_, _42382_);
  and (_42392_, _42319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_42393_, _42307_, _42283_);
  or (_02834_, _42393_, _42392_);
  and (_42394_, _42317_, _41746_);
  and (_42395_, _42286_, _41945_);
  and (_42396_, _42395_, _42301_);
  and (_42397_, _42396_, _42394_);
  not (_42398_, _42396_);
  and (_42399_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_02842_, _42399_, _42397_);
  and (_42400_, _42330_, _41746_);
  and (_42401_, _42396_, _42400_);
  and (_42402_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_02845_, _42402_, _42401_);
  and (_42403_, _42341_, _41746_);
  and (_42404_, _42396_, _42403_);
  and (_42405_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_02848_, _42405_, _42404_);
  and (_42406_, _42357_, _41746_);
  and (_42407_, _42396_, _42406_);
  and (_42408_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_02852_, _42408_, _42407_);
  and (_42409_, _42370_, _41746_);
  and (_42410_, _42396_, _42409_);
  and (_42411_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_02856_, _42411_, _42410_);
  and (_42412_, _42379_, _41746_);
  and (_42413_, _42396_, _42412_);
  and (_42414_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_02859_, _42414_, _42413_);
  and (_42415_, _42390_, _41746_);
  and (_42416_, _42396_, _42415_);
  and (_42417_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_02862_, _42417_, _42416_);
  and (_42418_, _42396_, _42294_);
  and (_42419_, _42398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_02865_, _42419_, _42418_);
  and (_42420_, _42287_, _41951_);
  and (_42421_, _42420_, _42301_);
  and (_42422_, _42421_, _42394_);
  not (_42423_, _42421_);
  and (_42424_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_02871_, _42424_, _42422_);
  and (_42425_, _42421_, _42400_);
  and (_42426_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_02875_, _42426_, _42425_);
  and (_42427_, _42421_, _42403_);
  and (_42428_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_02879_, _42428_, _42427_);
  and (_42429_, _42421_, _42406_);
  and (_42430_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_02882_, _42430_, _42429_);
  and (_42431_, _42421_, _42409_);
  and (_42432_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_02886_, _42432_, _42431_);
  and (_42433_, _42421_, _42412_);
  and (_42434_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_02889_, _42434_, _42433_);
  and (_42435_, _42421_, _42415_);
  and (_42436_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_02893_, _42436_, _42435_);
  and (_42437_, _42421_, _42294_);
  and (_42438_, _42423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_02895_, _42438_, _42437_);
  and (_42439_, _42301_, _42288_);
  and (_42440_, _42439_, _42394_);
  not (_42441_, _42439_);
  and (_42442_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_02901_, _42442_, _42440_);
  and (_42443_, _42439_, _42400_);
  and (_42444_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_02904_, _42444_, _42443_);
  and (_42445_, _42439_, _42403_);
  and (_42446_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_02907_, _42446_, _42445_);
  and (_42447_, _42439_, _42406_);
  and (_42448_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_02911_, _42448_, _42447_);
  and (_42449_, _42439_, _42409_);
  and (_42450_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_02913_, _42450_, _42449_);
  and (_42451_, _42439_, _42412_);
  and (_42452_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_02917_, _42452_, _42451_);
  and (_42453_, _42439_, _42415_);
  and (_42454_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_02921_, _42454_, _42453_);
  and (_42455_, _42439_, _42294_);
  and (_42456_, _42441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_02924_, _42456_, _42455_);
  and (_42457_, _42290_, _42047_);
  and (_42458_, _42457_, _42303_);
  and (_42459_, _42458_, _42394_);
  not (_42460_, _42458_);
  and (_42461_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_02933_, _42461_, _42459_);
  and (_42462_, _42458_, _42400_);
  and (_42463_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_02936_, _42463_, _42462_);
  and (_42464_, _42458_, _42403_);
  and (_42465_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_02940_, _42465_, _42464_);
  and (_42466_, _42458_, _42406_);
  and (_42467_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_02944_, _42467_, _42466_);
  and (_42468_, _42458_, _42409_);
  and (_42469_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_02948_, _42469_, _42468_);
  and (_42470_, _42458_, _42412_);
  and (_42471_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_02951_, _42471_, _42470_);
  and (_42472_, _42458_, _42415_);
  and (_42473_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_02955_, _42473_, _42472_);
  and (_42474_, _42458_, _42294_);
  and (_42475_, _42460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_02959_, _42475_, _42474_);
  and (_42476_, _42457_, _42395_);
  and (_42477_, _42476_, _42394_);
  not (_42478_, _42476_);
  and (_42479_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_02964_, _42479_, _42477_);
  and (_42480_, _42476_, _42400_);
  and (_42481_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_02968_, _42481_, _42480_);
  and (_42482_, _42476_, _42403_);
  and (_42483_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_02973_, _42483_, _42482_);
  and (_42484_, _42476_, _42406_);
  and (_42485_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_02976_, _42485_, _42484_);
  and (_42486_, _42476_, _42409_);
  and (_42487_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_02980_, _42487_, _42486_);
  and (_42488_, _42476_, _42412_);
  and (_42489_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_02985_, _42489_, _42488_);
  and (_42490_, _42476_, _42415_);
  and (_42491_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_02989_, _42491_, _42490_);
  and (_42492_, _42476_, _42294_);
  and (_42493_, _42478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_02992_, _42493_, _42492_);
  and (_42494_, _42457_, _42420_);
  and (_42495_, _42494_, _42394_);
  not (_42496_, _42494_);
  and (_42497_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_02996_, _42497_, _42495_);
  and (_42498_, _42494_, _42400_);
  and (_42499_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_03001_, _42499_, _42498_);
  and (_42500_, _42494_, _42403_);
  and (_42501_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_03004_, _42501_, _42500_);
  and (_42502_, _42494_, _42406_);
  and (_42503_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_03008_, _42503_, _42502_);
  and (_42504_, _42494_, _42409_);
  and (_42505_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_03013_, _42505_, _42504_);
  and (_42506_, _42494_, _42412_);
  and (_42507_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_03016_, _42507_, _42506_);
  and (_42508_, _42494_, _42415_);
  and (_42509_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_03019_, _42509_, _42508_);
  and (_42510_, _42494_, _42294_);
  and (_42511_, _42496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_03022_, _42511_, _42510_);
  and (_42512_, _42457_, _42288_);
  and (_42513_, _42512_, _42394_);
  not (_42514_, _42512_);
  and (_42515_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_03027_, _42515_, _42513_);
  and (_42516_, _42512_, _42400_);
  and (_42517_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_03030_, _42517_, _42516_);
  and (_42518_, _42512_, _42403_);
  and (_42519_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_03033_, _42519_, _42518_);
  and (_42520_, _42512_, _42406_);
  and (_42521_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_03036_, _42521_, _42520_);
  and (_42522_, _42512_, _42409_);
  and (_42523_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_03040_, _42523_, _42522_);
  and (_42524_, _42512_, _42412_);
  and (_42525_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_03043_, _42525_, _42524_);
  and (_42526_, _42512_, _42415_);
  and (_42527_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_03046_, _42527_, _42526_);
  and (_42528_, _42512_, _42294_);
  and (_42529_, _42514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_03049_, _42529_, _42528_);
  and (_42530_, _42289_, _42185_);
  and (_42531_, _42530_, _42303_);
  and (_42532_, _42531_, _42394_);
  not (_42533_, _42531_);
  and (_42534_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_03056_, _42534_, _42532_);
  and (_42535_, _42531_, _42400_);
  and (_42536_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_03060_, _42536_, _42535_);
  and (_42537_, _42531_, _42403_);
  and (_42538_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_03063_, _42538_, _42537_);
  and (_42539_, _42531_, _42406_);
  and (_42540_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_03067_, _42540_, _42539_);
  and (_42541_, _42531_, _42409_);
  and (_42542_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_03070_, _42542_, _42541_);
  and (_42543_, _42531_, _42412_);
  and (_42544_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_03074_, _42544_, _42543_);
  and (_42545_, _42531_, _42415_);
  and (_42546_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_03077_, _42546_, _42545_);
  and (_42547_, _42531_, _42294_);
  and (_42548_, _42533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_03080_, _42548_, _42547_);
  and (_42549_, _42530_, _42395_);
  and (_42550_, _42549_, _42394_);
  not (_42551_, _42549_);
  and (_42552_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_03085_, _42552_, _42550_);
  and (_42553_, _42549_, _42400_);
  and (_42554_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_03088_, _42554_, _42553_);
  and (_42555_, _42549_, _42403_);
  and (_42556_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_03092_, _42556_, _42555_);
  and (_42557_, _42549_, _42406_);
  and (_42558_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_03095_, _42558_, _42557_);
  and (_42559_, _42549_, _42409_);
  and (_42560_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_03099_, _42560_, _42559_);
  and (_42561_, _42549_, _42412_);
  and (_42562_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_03102_, _42562_, _42561_);
  and (_42563_, _42549_, _42415_);
  and (_42564_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_03106_, _42564_, _42563_);
  and (_42565_, _42549_, _42294_);
  and (_42566_, _42551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_03108_, _42566_, _42565_);
  and (_42567_, _42530_, _42420_);
  and (_42568_, _42567_, _42394_);
  not (_42569_, _42567_);
  and (_42570_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_03113_, _42570_, _42568_);
  and (_42571_, _42567_, _42400_);
  and (_42572_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_03116_, _42572_, _42571_);
  and (_42573_, _42567_, _42403_);
  and (_42574_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_03119_, _42574_, _42573_);
  and (_42575_, _42567_, _42406_);
  and (_42576_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_03123_, _42576_, _42575_);
  and (_42577_, _42567_, _42409_);
  and (_42578_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_03127_, _42578_, _42577_);
  and (_42579_, _42567_, _42412_);
  and (_42580_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_03130_, _42580_, _42579_);
  and (_42581_, _42567_, _42415_);
  and (_42582_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_03133_, _42582_, _42581_);
  and (_42583_, _42567_, _42294_);
  and (_42584_, _42569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_03136_, _42584_, _42583_);
  and (_42585_, _42530_, _42288_);
  and (_42586_, _42585_, _42394_);
  not (_42587_, _42585_);
  and (_42588_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_03140_, _42588_, _42586_);
  and (_42589_, _42585_, _42400_);
  and (_42590_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_03143_, _42590_, _42589_);
  and (_42591_, _42585_, _42403_);
  and (_42592_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_03146_, _42592_, _42591_);
  and (_42593_, _42585_, _42406_);
  and (_42594_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_03150_, _42594_, _42593_);
  and (_42595_, _42585_, _42409_);
  and (_42596_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_03153_, _42596_, _42595_);
  and (_42597_, _42585_, _42412_);
  and (_42598_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_03156_, _42598_, _42597_);
  and (_42599_, _42585_, _42415_);
  and (_42600_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_03159_, _42600_, _42599_);
  and (_42601_, _42585_, _42294_);
  and (_42602_, _42587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_03162_, _42602_, _42601_);
  and (_42603_, _42303_, _42291_);
  and (_42604_, _42603_, _42394_);
  not (_42605_, _42603_);
  and (_42606_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_03167_, _42606_, _42604_);
  and (_42607_, _42603_, _42400_);
  and (_42608_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_03170_, _42608_, _42607_);
  and (_42609_, _42603_, _42403_);
  and (_42610_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_03173_, _42610_, _42609_);
  and (_42611_, _42603_, _42406_);
  and (_42612_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_03176_, _42612_, _42611_);
  and (_42613_, _42603_, _42409_);
  and (_42614_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_03180_, _42614_, _42613_);
  and (_42615_, _42603_, _42412_);
  and (_42616_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_03183_, _42616_, _42615_);
  and (_42617_, _42603_, _42415_);
  and (_42618_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_03186_, _42618_, _42617_);
  and (_42619_, _42603_, _42294_);
  and (_42620_, _42605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_03189_, _42620_, _42619_);
  and (_42621_, _42395_, _42291_);
  and (_42622_, _42621_, _42394_);
  not (_42623_, _42621_);
  and (_42624_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_03193_, _42624_, _42622_);
  and (_42625_, _42621_, _42400_);
  and (_42626_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_03196_, _42626_, _42625_);
  and (_42627_, _42621_, _42403_);
  and (_42628_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_03199_, _42628_, _42627_);
  and (_42629_, _42621_, _42406_);
  and (_42630_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_03203_, _42630_, _42629_);
  and (_42631_, _42621_, _42409_);
  and (_42632_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_03206_, _42632_, _42631_);
  and (_42633_, _42621_, _42412_);
  and (_42634_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_03209_, _42634_, _42633_);
  and (_42635_, _42621_, _42415_);
  and (_42636_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_03213_, _42636_, _42635_);
  and (_42637_, _42621_, _42294_);
  and (_42638_, _42623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_03215_, _42638_, _42637_);
  and (_42639_, _42420_, _42291_);
  and (_42640_, _42639_, _42394_);
  not (_42641_, _42639_);
  and (_42642_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_03219_, _42642_, _42640_);
  and (_42643_, _42639_, _42400_);
  and (_42644_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_03222_, _42644_, _42643_);
  and (_42645_, _42639_, _42403_);
  and (_42646_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_03226_, _42646_, _42645_);
  and (_42647_, _42639_, _42406_);
  and (_42648_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_03229_, _42648_, _42647_);
  and (_42649_, _42639_, _42409_);
  and (_42650_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_03232_, _42650_, _42649_);
  and (_42651_, _42639_, _42412_);
  and (_42652_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_03236_, _42652_, _42651_);
  and (_42653_, _42639_, _42415_);
  and (_42654_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_03240_, _42654_, _42653_);
  and (_42655_, _42639_, _42294_);
  and (_42656_, _42641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_03243_, _42656_, _42655_);
  and (_42657_, _42394_, _42292_);
  and (_42658_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_03247_, _42658_, _42657_);
  and (_42659_, _42400_, _42292_);
  and (_42660_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_03251_, _42660_, _42659_);
  and (_42661_, _42403_, _42292_);
  and (_42662_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_03254_, _42662_, _42661_);
  and (_42663_, _42406_, _42292_);
  and (_42664_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_03257_, _42664_, _42663_);
  and (_42665_, _42409_, _42292_);
  and (_42666_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_03261_, _42666_, _42665_);
  and (_42667_, _42412_, _42292_);
  and (_42668_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_03264_, _42668_, _42667_);
  and (_42669_, _42415_, _42292_);
  and (_42670_, _42297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_03267_, _42670_, _42669_);
  and (_42671_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_42672_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_42673_, _42672_, _41941_);
  or (_42674_, _42673_, _42671_);
  and (_42675_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_42676_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_42677_, _42676_, _42225_);
  or (_42678_, _42677_, _42675_);
  and (_42679_, _42678_, _42674_);
  or (_42680_, _42679_, _42218_);
  and (_42681_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_42682_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_42683_, _42682_, _41941_);
  or (_42684_, _42683_, _42681_);
  and (_42685_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_42686_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_42687_, _42686_, _42225_);
  or (_42688_, _42687_, _42685_);
  and (_42689_, _42688_, _42684_);
  or (_42690_, _42689_, _42182_);
  and (_42691_, _42690_, _42231_);
  and (_42692_, _42691_, _42680_);
  or (_42693_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_42694_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_42695_, _42694_, _42693_);
  or (_42696_, _42695_, _42225_);
  or (_42697_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_42698_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_42699_, _42698_, _42697_);
  or (_42700_, _42699_, _41941_);
  and (_42701_, _42700_, _42696_);
  or (_42702_, _42701_, _42218_);
  or (_42703_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_42704_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_42705_, _42704_, _42703_);
  or (_42706_, _42705_, _42225_);
  or (_42707_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_42708_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_42709_, _42708_, _42707_);
  or (_42710_, _42709_, _41941_);
  and (_42711_, _42710_, _42706_);
  or (_42712_, _42711_, _42182_);
  and (_42713_, _42712_, _42091_);
  and (_42714_, _42713_, _42702_);
  or (_42715_, _42714_, _42692_);
  or (_42716_, _42715_, _42217_);
  or (_42717_, _42268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_42718_, _42717_, _42272_);
  and (_42719_, _42718_, _42716_);
  and (_39602_, _42317_, _42355_);
  and (_42720_, _39602_, _42271_);
  or (_05058_, _42720_, _42719_);
  and (_42721_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_42722_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_42723_, _42722_, _41941_);
  or (_42724_, _42723_, _42721_);
  and (_42725_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_42726_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_42727_, _42726_, _42225_);
  or (_42728_, _42727_, _42725_);
  and (_42729_, _42728_, _42724_);
  or (_42730_, _42729_, _42218_);
  and (_42731_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_42732_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_42733_, _42732_, _41941_);
  or (_42734_, _42733_, _42731_);
  and (_42735_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_42736_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_42737_, _42736_, _42225_);
  or (_42738_, _42737_, _42735_);
  and (_42739_, _42738_, _42734_);
  or (_42740_, _42739_, _42182_);
  and (_42741_, _42740_, _42231_);
  and (_42742_, _42741_, _42730_);
  or (_42743_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_42744_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_42745_, _42744_, _42743_);
  or (_42746_, _42745_, _42225_);
  or (_42747_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_42748_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_42749_, _42748_, _42747_);
  or (_42750_, _42749_, _41941_);
  and (_42751_, _42750_, _42746_);
  or (_42752_, _42751_, _42218_);
  or (_42753_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_42754_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_42755_, _42754_, _42753_);
  or (_42756_, _42755_, _42225_);
  or (_42757_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_42758_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_42759_, _42758_, _42757_);
  or (_42760_, _42759_, _41941_);
  and (_42761_, _42760_, _42756_);
  or (_42762_, _42761_, _42182_);
  and (_42763_, _42762_, _42091_);
  and (_42764_, _42763_, _42752_);
  or (_42765_, _42764_, _42742_);
  or (_42766_, _42765_, _42217_);
  or (_42767_, _42268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_42768_, _42767_, _42272_);
  and (_42769_, _42768_, _42766_);
  and (_39603_, _42330_, _42355_);
  and (_42770_, _39603_, _42271_);
  or (_05060_, _42770_, _42769_);
  and (_42771_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_42772_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_42773_, _42772_, _41941_);
  or (_42774_, _42773_, _42771_);
  and (_42775_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_42776_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_42777_, _42776_, _42225_);
  or (_42778_, _42777_, _42775_);
  and (_42779_, _42778_, _42774_);
  or (_42780_, _42779_, _42218_);
  and (_42781_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_42782_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_42783_, _42782_, _41941_);
  or (_42784_, _42783_, _42781_);
  and (_42785_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_42786_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_42787_, _42786_, _42225_);
  or (_42788_, _42787_, _42785_);
  and (_42789_, _42788_, _42784_);
  or (_42790_, _42789_, _42182_);
  and (_42791_, _42790_, _42231_);
  and (_42792_, _42791_, _42780_);
  or (_42793_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_42794_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_42795_, _42794_, _42793_);
  or (_42796_, _42795_, _42225_);
  or (_42797_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_42798_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_42799_, _42798_, _42797_);
  or (_42800_, _42799_, _41941_);
  and (_42801_, _42800_, _42796_);
  or (_42802_, _42801_, _42218_);
  or (_42803_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_42804_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_42805_, _42804_, _42803_);
  or (_42806_, _42805_, _42225_);
  or (_42807_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_42808_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_42809_, _42808_, _42807_);
  or (_42810_, _42809_, _41941_);
  and (_42811_, _42810_, _42806_);
  or (_42812_, _42811_, _42182_);
  and (_42813_, _42812_, _42091_);
  and (_42814_, _42813_, _42802_);
  or (_42815_, _42814_, _42792_);
  or (_42816_, _42815_, _42217_);
  or (_42817_, _42268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_42818_, _42817_, _42272_);
  and (_42819_, _42818_, _42816_);
  and (_39604_, _42341_, _42355_);
  and (_42820_, _39604_, _42271_);
  or (_05062_, _42820_, _42819_);
  or (_42821_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_42822_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_42823_, _42822_, _42821_);
  or (_42824_, _42823_, _41941_);
  or (_42825_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_42826_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_42827_, _42826_, _42825_);
  or (_42828_, _42827_, _42225_);
  and (_42829_, _42828_, _42091_);
  and (_42830_, _42829_, _42824_);
  and (_42831_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_42832_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_42833_, _42832_, _42225_);
  or (_42834_, _42833_, _42831_);
  and (_42835_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_42836_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_42837_, _42836_, _41941_);
  or (_42838_, _42837_, _42835_);
  and (_42839_, _42838_, _42231_);
  and (_42840_, _42839_, _42834_);
  or (_42841_, _42840_, _42830_);
  and (_42842_, _42841_, _42218_);
  or (_42843_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_42844_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_42845_, _42844_, _42843_);
  or (_42846_, _42845_, _41941_);
  or (_42847_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_42848_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_42849_, _42848_, _42847_);
  or (_42850_, _42849_, _42225_);
  and (_42851_, _42850_, _42091_);
  and (_42852_, _42851_, _42846_);
  and (_42853_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_42854_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_42855_, _42854_, _42225_);
  or (_42856_, _42855_, _42853_);
  and (_42857_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_42858_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_42859_, _42858_, _41941_);
  or (_42860_, _42859_, _42857_);
  and (_42861_, _42860_, _42231_);
  and (_42862_, _42861_, _42856_);
  or (_42863_, _42862_, _42852_);
  and (_42864_, _42863_, _42182_);
  or (_42865_, _42864_, _42192_);
  or (_42866_, _42865_, _42842_);
  or (_42867_, _42268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_39605_, _42357_, _42355_);
  or (_42868_, _39605_, _42272_);
  and (_42869_, _42868_, _42867_);
  and (_05064_, _42869_, _42866_);
  and (_42870_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_42871_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_42872_, _42871_, _42225_);
  or (_42873_, _42872_, _42870_);
  and (_42874_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_42875_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_42876_, _42875_, _41941_);
  or (_42877_, _42876_, _42874_);
  and (_42878_, _42877_, _42873_);
  or (_42879_, _42878_, _42218_);
  and (_42880_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_42881_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_42882_, _42881_, _41941_);
  or (_42883_, _42882_, _42880_);
  and (_42884_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_42885_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_42886_, _42885_, _42225_);
  or (_42887_, _42886_, _42884_);
  and (_42888_, _42887_, _42883_);
  or (_42889_, _42888_, _42182_);
  and (_42895_, _42889_, _42231_);
  and (_42899_, _42895_, _42879_);
  and (_42906_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_42914_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_42918_, _42914_, _41941_);
  or (_42923_, _42918_, _42906_);
  and (_42931_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_42937_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_42941_, _42937_, _42225_);
  or (_42948_, _42941_, _42931_);
  and (_42956_, _42948_, _42923_);
  or (_42960_, _42956_, _42218_);
  and (_42965_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_42973_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_42979_, _42973_, _41941_);
  or (_42982_, _42979_, _42965_);
  and (_42986_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_42997_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_43001_, _42997_, _42225_);
  or (_43008_, _43001_, _42986_);
  and (_43016_, _43008_, _42982_);
  or (_43020_, _43016_, _42182_);
  and (_43025_, _43020_, _42091_);
  and (_43033_, _43025_, _42960_);
  or (_43039_, _43033_, _42899_);
  and (_43043_, _43039_, _42270_);
  and (_43050_, _42370_, _42271_);
  and (_43058_, _42217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_43062_, _43058_, _43050_);
  or (_43067_, _43062_, _43043_);
  and (_05066_, _43067_, _42355_);
  and (_43080_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_43083_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_43084_, _43083_, _41941_);
  or (_43085_, _43084_, _43080_);
  and (_43086_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_43087_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_43088_, _43087_, _42225_);
  or (_43089_, _43088_, _43086_);
  and (_43090_, _43089_, _43085_);
  or (_43091_, _43090_, _42218_);
  and (_43092_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_43093_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_43094_, _43093_, _41941_);
  or (_43095_, _43094_, _43092_);
  and (_43096_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_43097_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_43098_, _43097_, _42225_);
  or (_43099_, _43098_, _43096_);
  and (_43100_, _43099_, _43095_);
  or (_43101_, _43100_, _42182_);
  and (_43102_, _43101_, _42231_);
  and (_43103_, _43102_, _43091_);
  or (_43104_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_43105_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_43106_, _43105_, _43104_);
  or (_43107_, _43106_, _42225_);
  or (_43108_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_43109_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_43110_, _43109_, _43108_);
  or (_43111_, _43110_, _41941_);
  and (_43112_, _43111_, _43107_);
  or (_43113_, _43112_, _42218_);
  or (_43114_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_43115_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_43116_, _43115_, _43114_);
  or (_43117_, _43116_, _42225_);
  or (_43118_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_43119_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_43120_, _43119_, _43118_);
  or (_43121_, _43120_, _41941_);
  and (_43122_, _43121_, _43117_);
  or (_43123_, _43122_, _42182_);
  and (_43124_, _43123_, _42091_);
  and (_43125_, _43124_, _43113_);
  or (_43126_, _43125_, _43103_);
  or (_43127_, _43126_, _42217_);
  or (_43128_, _42268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_43129_, _43128_, _42272_);
  and (_43130_, _43129_, _43127_);
  and (_39607_, _42379_, _42355_);
  and (_43131_, _39607_, _42271_);
  or (_05068_, _43131_, _43130_);
  and (_43132_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_43133_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_43134_, _43133_, _41941_);
  or (_43135_, _43134_, _43132_);
  and (_43136_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_43137_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_43138_, _43137_, _42225_);
  or (_43139_, _43138_, _43136_);
  and (_43140_, _43139_, _43135_);
  or (_43141_, _43140_, _42218_);
  and (_43142_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_43143_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_43144_, _43143_, _41941_);
  or (_43145_, _43144_, _43142_);
  and (_43146_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_43147_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_43148_, _43147_, _42225_);
  or (_43149_, _43148_, _43146_);
  and (_43150_, _43149_, _43145_);
  or (_43151_, _43150_, _42182_);
  and (_43152_, _43151_, _42231_);
  and (_43153_, _43152_, _43141_);
  or (_43154_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_43155_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_43156_, _43155_, _43154_);
  or (_43157_, _43156_, _42225_);
  or (_43158_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_43159_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_43160_, _43159_, _43158_);
  or (_43161_, _43160_, _41941_);
  and (_43162_, _43161_, _43157_);
  or (_43163_, _43162_, _42218_);
  or (_43164_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_43165_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_43166_, _43165_, _43164_);
  or (_43167_, _43166_, _42225_);
  or (_43168_, _42039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_43169_, _42219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_43170_, _43169_, _43168_);
  or (_43171_, _43170_, _41941_);
  and (_43172_, _43171_, _43167_);
  or (_43173_, _43172_, _42182_);
  and (_43174_, _43173_, _42091_);
  and (_43175_, _43174_, _43163_);
  or (_43176_, _43175_, _43153_);
  or (_43177_, _43176_, _42217_);
  or (_43178_, _42268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_43179_, _43178_, _42272_);
  and (_43180_, _43179_, _43177_);
  and (_39608_, _42390_, _42355_);
  and (_43181_, _39608_, _42271_);
  or (_05069_, _43181_, _43180_);
  or (_43182_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_43183_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_43184_, _43183_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_43185_, _43184_, _43182_);
  nand (_43186_, _43185_, _42355_);
  or (_43187_, \oc8051_gm_cxrom_1.cell0.data [7], _42355_);
  and (_05077_, _43187_, _43186_);
  or (_43188_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43189_, \oc8051_gm_cxrom_1.cell0.data [0], _43183_);
  nand (_43190_, _43189_, _43188_);
  nand (_43191_, _43190_, _42355_);
  or (_43192_, \oc8051_gm_cxrom_1.cell0.data [0], _42355_);
  and (_05084_, _43192_, _43191_);
  or (_43193_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43194_, \oc8051_gm_cxrom_1.cell0.data [1], _43183_);
  nand (_43195_, _43194_, _43193_);
  nand (_43196_, _43195_, _42355_);
  or (_43197_, \oc8051_gm_cxrom_1.cell0.data [1], _42355_);
  and (_05088_, _43197_, _43196_);
  or (_43198_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43199_, \oc8051_gm_cxrom_1.cell0.data [2], _43183_);
  nand (_43200_, _43199_, _43198_);
  nand (_43201_, _43200_, _42355_);
  or (_43202_, \oc8051_gm_cxrom_1.cell0.data [2], _42355_);
  and (_05092_, _43202_, _43201_);
  or (_43203_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43204_, \oc8051_gm_cxrom_1.cell0.data [3], _43183_);
  nand (_43205_, _43204_, _43203_);
  nand (_43206_, _43205_, _42355_);
  or (_43207_, \oc8051_gm_cxrom_1.cell0.data [3], _42355_);
  and (_05096_, _43207_, _43206_);
  or (_43208_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43209_, \oc8051_gm_cxrom_1.cell0.data [4], _43183_);
  nand (_43210_, _43209_, _43208_);
  nand (_43211_, _43210_, _42355_);
  or (_43212_, \oc8051_gm_cxrom_1.cell0.data [4], _42355_);
  and (_05100_, _43212_, _43211_);
  or (_43213_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43214_, \oc8051_gm_cxrom_1.cell0.data [5], _43183_);
  nand (_43215_, _43214_, _43213_);
  nand (_43216_, _43215_, _42355_);
  or (_43217_, \oc8051_gm_cxrom_1.cell0.data [5], _42355_);
  and (_05104_, _43217_, _43216_);
  or (_43218_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_43219_, \oc8051_gm_cxrom_1.cell0.data [6], _43183_);
  nand (_43220_, _43219_, _43218_);
  nand (_43221_, _43220_, _42355_);
  or (_43222_, \oc8051_gm_cxrom_1.cell0.data [6], _42355_);
  and (_05108_, _43222_, _43221_);
  or (_43223_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_43224_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_43225_, _43224_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_43226_, _43225_, _43223_);
  nand (_43227_, _43226_, _42355_);
  or (_43228_, \oc8051_gm_cxrom_1.cell1.data [7], _42355_);
  and (_05129_, _43228_, _43227_);
  or (_43229_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43230_, \oc8051_gm_cxrom_1.cell1.data [0], _43224_);
  nand (_43231_, _43230_, _43229_);
  nand (_43232_, _43231_, _42355_);
  or (_43233_, \oc8051_gm_cxrom_1.cell1.data [0], _42355_);
  and (_05136_, _43233_, _43232_);
  or (_43234_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43235_, \oc8051_gm_cxrom_1.cell1.data [1], _43224_);
  nand (_43236_, _43235_, _43234_);
  nand (_43237_, _43236_, _42355_);
  or (_43238_, \oc8051_gm_cxrom_1.cell1.data [1], _42355_);
  and (_05140_, _43238_, _43237_);
  or (_43239_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43240_, \oc8051_gm_cxrom_1.cell1.data [2], _43224_);
  nand (_43241_, _43240_, _43239_);
  nand (_43242_, _43241_, _42355_);
  or (_43243_, \oc8051_gm_cxrom_1.cell1.data [2], _42355_);
  and (_05143_, _43243_, _43242_);
  or (_43244_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43245_, \oc8051_gm_cxrom_1.cell1.data [3], _43224_);
  nand (_43246_, _43245_, _43244_);
  nand (_43247_, _43246_, _42355_);
  or (_43248_, \oc8051_gm_cxrom_1.cell1.data [3], _42355_);
  and (_05147_, _43248_, _43247_);
  or (_43249_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43250_, \oc8051_gm_cxrom_1.cell1.data [4], _43224_);
  nand (_43251_, _43250_, _43249_);
  nand (_43252_, _43251_, _42355_);
  or (_43253_, \oc8051_gm_cxrom_1.cell1.data [4], _42355_);
  and (_05151_, _43253_, _43252_);
  or (_43254_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43255_, \oc8051_gm_cxrom_1.cell1.data [5], _43224_);
  nand (_43256_, _43255_, _43254_);
  nand (_43257_, _43256_, _42355_);
  or (_43258_, \oc8051_gm_cxrom_1.cell1.data [5], _42355_);
  and (_05155_, _43258_, _43257_);
  or (_43259_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_43260_, \oc8051_gm_cxrom_1.cell1.data [6], _43224_);
  nand (_43261_, _43260_, _43259_);
  nand (_43262_, _43261_, _42355_);
  or (_43263_, \oc8051_gm_cxrom_1.cell1.data [6], _42355_);
  and (_05159_, _43263_, _43262_);
  or (_43264_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_43265_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_43266_, _43265_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_43267_, _43266_, _43264_);
  nand (_00002_, _43267_, _42355_);
  or (_00003_, \oc8051_gm_cxrom_1.cell2.data [7], _42355_);
  and (_05180_, _00003_, _00002_);
  or (_00004_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00005_, \oc8051_gm_cxrom_1.cell2.data [0], _43265_);
  nand (_00006_, _00005_, _00004_);
  nand (_00007_, _00006_, _42355_);
  or (_00008_, \oc8051_gm_cxrom_1.cell2.data [0], _42355_);
  and (_05187_, _00008_, _00007_);
  or (_00009_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00010_, \oc8051_gm_cxrom_1.cell2.data [1], _43265_);
  nand (_00011_, _00010_, _00009_);
  nand (_00012_, _00011_, _42355_);
  or (_00013_, \oc8051_gm_cxrom_1.cell2.data [1], _42355_);
  and (_05191_, _00013_, _00012_);
  or (_00014_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00015_, \oc8051_gm_cxrom_1.cell2.data [2], _43265_);
  nand (_00016_, _00015_, _00014_);
  nand (_00017_, _00016_, _42355_);
  or (_00018_, \oc8051_gm_cxrom_1.cell2.data [2], _42355_);
  and (_05195_, _00018_, _00017_);
  or (_00019_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00020_, \oc8051_gm_cxrom_1.cell2.data [3], _43265_);
  nand (_00021_, _00020_, _00019_);
  nand (_00022_, _00021_, _42355_);
  or (_00023_, \oc8051_gm_cxrom_1.cell2.data [3], _42355_);
  and (_05199_, _00023_, _00022_);
  or (_00024_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00025_, \oc8051_gm_cxrom_1.cell2.data [4], _43265_);
  nand (_00026_, _00025_, _00024_);
  nand (_00027_, _00026_, _42355_);
  or (_00028_, \oc8051_gm_cxrom_1.cell2.data [4], _42355_);
  and (_05203_, _00028_, _00027_);
  or (_00029_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00030_, \oc8051_gm_cxrom_1.cell2.data [5], _43265_);
  nand (_00031_, _00030_, _00029_);
  nand (_00032_, _00031_, _42355_);
  or (_00033_, \oc8051_gm_cxrom_1.cell2.data [5], _42355_);
  and (_05207_, _00033_, _00032_);
  or (_00034_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_00035_, \oc8051_gm_cxrom_1.cell2.data [6], _43265_);
  nand (_00036_, _00035_, _00034_);
  nand (_00037_, _00036_, _42355_);
  or (_00038_, \oc8051_gm_cxrom_1.cell2.data [6], _42355_);
  and (_05211_, _00038_, _00037_);
  or (_00039_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_00040_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_00041_, _00040_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_00042_, _00041_, _00039_);
  nand (_00043_, _00042_, _42355_);
  or (_00044_, \oc8051_gm_cxrom_1.cell3.data [7], _42355_);
  and (_05232_, _00044_, _00043_);
  or (_00045_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00046_, \oc8051_gm_cxrom_1.cell3.data [0], _00040_);
  nand (_00047_, _00046_, _00045_);
  nand (_00048_, _00047_, _42355_);
  or (_00049_, \oc8051_gm_cxrom_1.cell3.data [0], _42355_);
  and (_05239_, _00049_, _00048_);
  or (_00050_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00051_, \oc8051_gm_cxrom_1.cell3.data [1], _00040_);
  nand (_00052_, _00051_, _00050_);
  nand (_00053_, _00052_, _42355_);
  or (_00054_, \oc8051_gm_cxrom_1.cell3.data [1], _42355_);
  and (_05243_, _00054_, _00053_);
  or (_00055_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00056_, \oc8051_gm_cxrom_1.cell3.data [2], _00040_);
  nand (_00057_, _00056_, _00055_);
  nand (_00058_, _00057_, _42355_);
  or (_00059_, \oc8051_gm_cxrom_1.cell3.data [2], _42355_);
  and (_05247_, _00059_, _00058_);
  or (_00060_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00061_, \oc8051_gm_cxrom_1.cell3.data [3], _00040_);
  nand (_00062_, _00061_, _00060_);
  nand (_00063_, _00062_, _42355_);
  or (_00064_, \oc8051_gm_cxrom_1.cell3.data [3], _42355_);
  and (_05251_, _00064_, _00063_);
  or (_00065_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00066_, \oc8051_gm_cxrom_1.cell3.data [4], _00040_);
  nand (_00067_, _00066_, _00065_);
  nand (_00068_, _00067_, _42355_);
  or (_00069_, \oc8051_gm_cxrom_1.cell3.data [4], _42355_);
  and (_05254_, _00069_, _00068_);
  or (_00070_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00071_, \oc8051_gm_cxrom_1.cell3.data [5], _00040_);
  nand (_00072_, _00071_, _00070_);
  nand (_00073_, _00072_, _42355_);
  or (_00074_, \oc8051_gm_cxrom_1.cell3.data [5], _42355_);
  and (_05258_, _00074_, _00073_);
  or (_00075_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_00076_, \oc8051_gm_cxrom_1.cell3.data [6], _00040_);
  nand (_00077_, _00076_, _00075_);
  nand (_00078_, _00077_, _42355_);
  or (_00079_, \oc8051_gm_cxrom_1.cell3.data [6], _42355_);
  and (_05262_, _00079_, _00078_);
  or (_00080_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_00081_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_00082_, _00081_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_00083_, _00082_, _00080_);
  nand (_00084_, _00083_, _42355_);
  or (_00085_, \oc8051_gm_cxrom_1.cell4.data [7], _42355_);
  and (_05284_, _00085_, _00084_);
  or (_00086_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00087_, \oc8051_gm_cxrom_1.cell4.data [0], _00081_);
  nand (_00088_, _00087_, _00086_);
  nand (_00089_, _00088_, _42355_);
  or (_00090_, \oc8051_gm_cxrom_1.cell4.data [0], _42355_);
  and (_05290_, _00090_, _00089_);
  or (_00091_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00092_, \oc8051_gm_cxrom_1.cell4.data [1], _00081_);
  nand (_00093_, _00092_, _00091_);
  nand (_00094_, _00093_, _42355_);
  or (_00095_, \oc8051_gm_cxrom_1.cell4.data [1], _42355_);
  and (_05294_, _00095_, _00094_);
  or (_00096_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00097_, \oc8051_gm_cxrom_1.cell4.data [2], _00081_);
  nand (_00098_, _00097_, _00096_);
  nand (_00099_, _00098_, _42355_);
  or (_00100_, \oc8051_gm_cxrom_1.cell4.data [2], _42355_);
  and (_05298_, _00100_, _00099_);
  or (_00101_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00102_, \oc8051_gm_cxrom_1.cell4.data [3], _00081_);
  nand (_00103_, _00102_, _00101_);
  nand (_00104_, _00103_, _42355_);
  or (_00105_, \oc8051_gm_cxrom_1.cell4.data [3], _42355_);
  and (_05302_, _00105_, _00104_);
  or (_00106_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00107_, \oc8051_gm_cxrom_1.cell4.data [4], _00081_);
  nand (_00108_, _00107_, _00106_);
  nand (_00109_, _00108_, _42355_);
  or (_00110_, \oc8051_gm_cxrom_1.cell4.data [4], _42355_);
  and (_05306_, _00110_, _00109_);
  or (_00111_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00112_, \oc8051_gm_cxrom_1.cell4.data [5], _00081_);
  nand (_00113_, _00112_, _00111_);
  nand (_00114_, _00113_, _42355_);
  or (_00115_, \oc8051_gm_cxrom_1.cell4.data [5], _42355_);
  and (_05310_, _00115_, _00114_);
  or (_00116_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_00117_, \oc8051_gm_cxrom_1.cell4.data [6], _00081_);
  nand (_00118_, _00117_, _00116_);
  nand (_00119_, _00118_, _42355_);
  or (_00120_, \oc8051_gm_cxrom_1.cell4.data [6], _42355_);
  and (_05314_, _00120_, _00119_);
  or (_00121_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_00122_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_00123_, _00122_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_00124_, _00123_, _00121_);
  nand (_00125_, _00124_, _42355_);
  or (_00126_, \oc8051_gm_cxrom_1.cell5.data [7], _42355_);
  and (_05335_, _00126_, _00125_);
  or (_00127_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00128_, \oc8051_gm_cxrom_1.cell5.data [0], _00122_);
  nand (_00129_, _00128_, _00127_);
  nand (_00130_, _00129_, _42355_);
  or (_00132_, \oc8051_gm_cxrom_1.cell5.data [0], _42355_);
  and (_05342_, _00132_, _00130_);
  or (_00135_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00137_, \oc8051_gm_cxrom_1.cell5.data [1], _00122_);
  nand (_00139_, _00137_, _00135_);
  nand (_00141_, _00139_, _42355_);
  or (_00143_, \oc8051_gm_cxrom_1.cell5.data [1], _42355_);
  and (_05346_, _00143_, _00141_);
  or (_00146_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00148_, \oc8051_gm_cxrom_1.cell5.data [2], _00122_);
  nand (_00150_, _00148_, _00146_);
  nand (_00152_, _00150_, _42355_);
  or (_00154_, \oc8051_gm_cxrom_1.cell5.data [2], _42355_);
  and (_05350_, _00154_, _00152_);
  or (_00157_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00159_, \oc8051_gm_cxrom_1.cell5.data [3], _00122_);
  nand (_00161_, _00159_, _00157_);
  nand (_00163_, _00161_, _42355_);
  or (_00165_, \oc8051_gm_cxrom_1.cell5.data [3], _42355_);
  and (_05354_, _00165_, _00163_);
  or (_00168_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00170_, \oc8051_gm_cxrom_1.cell5.data [4], _00122_);
  nand (_00172_, _00170_, _00168_);
  nand (_00174_, _00172_, _42355_);
  or (_00176_, \oc8051_gm_cxrom_1.cell5.data [4], _42355_);
  and (_05358_, _00176_, _00174_);
  or (_00179_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00181_, \oc8051_gm_cxrom_1.cell5.data [5], _00122_);
  nand (_00183_, _00181_, _00179_);
  nand (_00185_, _00183_, _42355_);
  or (_00187_, \oc8051_gm_cxrom_1.cell5.data [5], _42355_);
  and (_05362_, _00187_, _00185_);
  or (_00188_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_00189_, \oc8051_gm_cxrom_1.cell5.data [6], _00122_);
  nand (_00190_, _00189_, _00188_);
  nand (_00191_, _00190_, _42355_);
  or (_00192_, \oc8051_gm_cxrom_1.cell5.data [6], _42355_);
  and (_05365_, _00192_, _00191_);
  or (_00193_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_00194_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_00195_, _00194_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_00196_, _00195_, _00193_);
  nand (_00197_, _00196_, _42355_);
  or (_00198_, \oc8051_gm_cxrom_1.cell6.data [7], _42355_);
  and (_05387_, _00198_, _00197_);
  or (_00199_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00200_, \oc8051_gm_cxrom_1.cell6.data [0], _00194_);
  nand (_00201_, _00200_, _00199_);
  nand (_00202_, _00201_, _42355_);
  or (_00203_, \oc8051_gm_cxrom_1.cell6.data [0], _42355_);
  and (_05394_, _00203_, _00202_);
  or (_00204_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00205_, \oc8051_gm_cxrom_1.cell6.data [1], _00194_);
  nand (_00206_, _00205_, _00204_);
  nand (_00207_, _00206_, _42355_);
  or (_00208_, \oc8051_gm_cxrom_1.cell6.data [1], _42355_);
  and (_05397_, _00208_, _00207_);
  or (_00209_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00210_, \oc8051_gm_cxrom_1.cell6.data [2], _00194_);
  nand (_00211_, _00210_, _00209_);
  nand (_00212_, _00211_, _42355_);
  or (_00213_, \oc8051_gm_cxrom_1.cell6.data [2], _42355_);
  and (_05401_, _00213_, _00212_);
  or (_00214_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00215_, \oc8051_gm_cxrom_1.cell6.data [3], _00194_);
  nand (_00216_, _00215_, _00214_);
  nand (_00217_, _00216_, _42355_);
  or (_00218_, \oc8051_gm_cxrom_1.cell6.data [3], _42355_);
  and (_05405_, _00218_, _00217_);
  or (_00219_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00220_, \oc8051_gm_cxrom_1.cell6.data [4], _00194_);
  nand (_00221_, _00220_, _00219_);
  nand (_00222_, _00221_, _42355_);
  or (_00223_, \oc8051_gm_cxrom_1.cell6.data [4], _42355_);
  and (_05409_, _00223_, _00222_);
  or (_00224_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00225_, \oc8051_gm_cxrom_1.cell6.data [5], _00194_);
  nand (_00226_, _00225_, _00224_);
  nand (_00227_, _00226_, _42355_);
  or (_00228_, \oc8051_gm_cxrom_1.cell6.data [5], _42355_);
  and (_05413_, _00228_, _00227_);
  or (_00229_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_00230_, \oc8051_gm_cxrom_1.cell6.data [6], _00194_);
  nand (_00231_, _00230_, _00229_);
  nand (_00232_, _00231_, _42355_);
  or (_00233_, \oc8051_gm_cxrom_1.cell6.data [6], _42355_);
  and (_05417_, _00233_, _00232_);
  or (_00234_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_00235_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_00236_, _00235_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_00237_, _00236_, _00234_);
  nand (_00238_, _00237_, _42355_);
  or (_00239_, \oc8051_gm_cxrom_1.cell7.data [7], _42355_);
  and (_05438_, _00239_, _00238_);
  or (_00240_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00241_, \oc8051_gm_cxrom_1.cell7.data [0], _00235_);
  nand (_00242_, _00241_, _00240_);
  nand (_00243_, _00242_, _42355_);
  or (_00244_, \oc8051_gm_cxrom_1.cell7.data [0], _42355_);
  and (_05445_, _00244_, _00243_);
  or (_00245_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00246_, \oc8051_gm_cxrom_1.cell7.data [1], _00235_);
  nand (_00247_, _00246_, _00245_);
  nand (_00248_, _00247_, _42355_);
  or (_00249_, \oc8051_gm_cxrom_1.cell7.data [1], _42355_);
  and (_05449_, _00249_, _00248_);
  or (_00250_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00251_, \oc8051_gm_cxrom_1.cell7.data [2], _00235_);
  nand (_00252_, _00251_, _00250_);
  nand (_00253_, _00252_, _42355_);
  or (_00254_, \oc8051_gm_cxrom_1.cell7.data [2], _42355_);
  and (_05453_, _00254_, _00253_);
  or (_00255_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00256_, \oc8051_gm_cxrom_1.cell7.data [3], _00235_);
  nand (_00257_, _00256_, _00255_);
  nand (_00258_, _00257_, _42355_);
  or (_00259_, \oc8051_gm_cxrom_1.cell7.data [3], _42355_);
  and (_05457_, _00259_, _00258_);
  or (_00260_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00261_, \oc8051_gm_cxrom_1.cell7.data [4], _00235_);
  nand (_00262_, _00261_, _00260_);
  nand (_00263_, _00262_, _42355_);
  or (_00264_, \oc8051_gm_cxrom_1.cell7.data [4], _42355_);
  and (_05461_, _00264_, _00263_);
  or (_00265_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00266_, \oc8051_gm_cxrom_1.cell7.data [5], _00235_);
  nand (_00267_, _00266_, _00265_);
  nand (_00268_, _00267_, _42355_);
  or (_00269_, \oc8051_gm_cxrom_1.cell7.data [5], _42355_);
  and (_05465_, _00269_, _00268_);
  or (_00270_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_00271_, \oc8051_gm_cxrom_1.cell7.data [6], _00235_);
  nand (_00272_, _00271_, _00270_);
  nand (_00273_, _00272_, _42355_);
  or (_00274_, \oc8051_gm_cxrom_1.cell7.data [6], _42355_);
  and (_05469_, _00274_, _00273_);
  or (_00275_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_00276_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_00277_, _00276_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_00278_, _00277_, _00275_);
  nand (_00279_, _00278_, _42355_);
  or (_00280_, \oc8051_gm_cxrom_1.cell8.data [7], _42355_);
  and (_05490_, _00280_, _00279_);
  or (_00281_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00282_, \oc8051_gm_cxrom_1.cell8.data [0], _00276_);
  nand (_00283_, _00282_, _00281_);
  nand (_00284_, _00283_, _42355_);
  or (_00285_, \oc8051_gm_cxrom_1.cell8.data [0], _42355_);
  and (_05497_, _00285_, _00284_);
  or (_00286_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00287_, \oc8051_gm_cxrom_1.cell8.data [1], _00276_);
  nand (_00288_, _00287_, _00286_);
  nand (_00289_, _00288_, _42355_);
  or (_00290_, \oc8051_gm_cxrom_1.cell8.data [1], _42355_);
  and (_05501_, _00290_, _00289_);
  or (_00291_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00292_, \oc8051_gm_cxrom_1.cell8.data [2], _00276_);
  nand (_00293_, _00292_, _00291_);
  nand (_00294_, _00293_, _42355_);
  or (_00295_, \oc8051_gm_cxrom_1.cell8.data [2], _42355_);
  and (_05505_, _00295_, _00294_);
  or (_00296_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00297_, \oc8051_gm_cxrom_1.cell8.data [3], _00276_);
  nand (_00298_, _00297_, _00296_);
  nand (_00299_, _00298_, _42355_);
  or (_00300_, \oc8051_gm_cxrom_1.cell8.data [3], _42355_);
  and (_05508_, _00300_, _00299_);
  or (_00301_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00302_, \oc8051_gm_cxrom_1.cell8.data [4], _00276_);
  nand (_00303_, _00302_, _00301_);
  nand (_00304_, _00303_, _42355_);
  or (_00305_, \oc8051_gm_cxrom_1.cell8.data [4], _42355_);
  and (_05512_, _00305_, _00304_);
  or (_00306_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00307_, \oc8051_gm_cxrom_1.cell8.data [5], _00276_);
  nand (_00308_, _00307_, _00306_);
  nand (_00309_, _00308_, _42355_);
  or (_00310_, \oc8051_gm_cxrom_1.cell8.data [5], _42355_);
  and (_05516_, _00310_, _00309_);
  or (_00311_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_00312_, \oc8051_gm_cxrom_1.cell8.data [6], _00276_);
  nand (_00313_, _00312_, _00311_);
  nand (_00314_, _00313_, _42355_);
  or (_00315_, \oc8051_gm_cxrom_1.cell8.data [6], _42355_);
  and (_05520_, _00315_, _00314_);
  or (_00316_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_00317_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_00318_, _00317_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_00319_, _00318_, _00316_);
  nand (_00320_, _00319_, _42355_);
  or (_00321_, \oc8051_gm_cxrom_1.cell9.data [7], _42355_);
  and (_05541_, _00321_, _00320_);
  or (_00322_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00323_, \oc8051_gm_cxrom_1.cell9.data [0], _00317_);
  nand (_00324_, _00323_, _00322_);
  nand (_00325_, _00324_, _42355_);
  or (_00326_, \oc8051_gm_cxrom_1.cell9.data [0], _42355_);
  and (_05548_, _00326_, _00325_);
  or (_00327_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00328_, \oc8051_gm_cxrom_1.cell9.data [1], _00317_);
  nand (_00329_, _00328_, _00327_);
  nand (_00330_, _00329_, _42355_);
  or (_00331_, \oc8051_gm_cxrom_1.cell9.data [1], _42355_);
  and (_05552_, _00331_, _00330_);
  or (_00332_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00333_, \oc8051_gm_cxrom_1.cell9.data [2], _00317_);
  nand (_00334_, _00333_, _00332_);
  nand (_00335_, _00334_, _42355_);
  or (_00336_, \oc8051_gm_cxrom_1.cell9.data [2], _42355_);
  and (_05556_, _00336_, _00335_);
  or (_00337_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00338_, \oc8051_gm_cxrom_1.cell9.data [3], _00317_);
  nand (_00339_, _00338_, _00337_);
  nand (_00340_, _00339_, _42355_);
  or (_00341_, \oc8051_gm_cxrom_1.cell9.data [3], _42355_);
  and (_05560_, _00341_, _00340_);
  or (_00342_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00343_, \oc8051_gm_cxrom_1.cell9.data [4], _00317_);
  nand (_00344_, _00343_, _00342_);
  nand (_00345_, _00344_, _42355_);
  or (_00346_, \oc8051_gm_cxrom_1.cell9.data [4], _42355_);
  and (_05564_, _00346_, _00345_);
  or (_00347_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00348_, \oc8051_gm_cxrom_1.cell9.data [5], _00317_);
  nand (_00349_, _00348_, _00347_);
  nand (_00350_, _00349_, _42355_);
  or (_00351_, \oc8051_gm_cxrom_1.cell9.data [5], _42355_);
  and (_05568_, _00351_, _00350_);
  or (_00352_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_00353_, \oc8051_gm_cxrom_1.cell9.data [6], _00317_);
  nand (_00354_, _00353_, _00352_);
  nand (_00355_, _00354_, _42355_);
  or (_00356_, \oc8051_gm_cxrom_1.cell9.data [6], _42355_);
  and (_05572_, _00356_, _00355_);
  or (_00357_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_00358_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_00359_, _00358_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_00360_, _00359_, _00357_);
  nand (_00361_, _00360_, _42355_);
  or (_00362_, \oc8051_gm_cxrom_1.cell10.data [7], _42355_);
  and (_05593_, _00362_, _00361_);
  or (_00363_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00364_, \oc8051_gm_cxrom_1.cell10.data [0], _00358_);
  nand (_00365_, _00364_, _00363_);
  nand (_00366_, _00365_, _42355_);
  or (_00367_, \oc8051_gm_cxrom_1.cell10.data [0], _42355_);
  and (_05600_, _00367_, _00366_);
  or (_00368_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00369_, \oc8051_gm_cxrom_1.cell10.data [1], _00358_);
  nand (_00370_, _00369_, _00368_);
  nand (_00371_, _00370_, _42355_);
  or (_00372_, \oc8051_gm_cxrom_1.cell10.data [1], _42355_);
  and (_05604_, _00372_, _00371_);
  or (_00373_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00374_, \oc8051_gm_cxrom_1.cell10.data [2], _00358_);
  nand (_00375_, _00374_, _00373_);
  nand (_00376_, _00375_, _42355_);
  or (_00377_, \oc8051_gm_cxrom_1.cell10.data [2], _42355_);
  and (_05608_, _00377_, _00376_);
  or (_00378_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00379_, \oc8051_gm_cxrom_1.cell10.data [3], _00358_);
  nand (_00380_, _00379_, _00378_);
  nand (_00381_, _00380_, _42355_);
  or (_00382_, \oc8051_gm_cxrom_1.cell10.data [3], _42355_);
  and (_05612_, _00382_, _00381_);
  or (_00383_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00384_, \oc8051_gm_cxrom_1.cell10.data [4], _00358_);
  nand (_00385_, _00384_, _00383_);
  nand (_00386_, _00385_, _42355_);
  or (_00387_, \oc8051_gm_cxrom_1.cell10.data [4], _42355_);
  and (_05616_, _00387_, _00386_);
  or (_00388_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00389_, \oc8051_gm_cxrom_1.cell10.data [5], _00358_);
  nand (_00390_, _00389_, _00388_);
  nand (_00391_, _00390_, _42355_);
  or (_00392_, \oc8051_gm_cxrom_1.cell10.data [5], _42355_);
  and (_05620_, _00392_, _00391_);
  or (_00393_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_00394_, \oc8051_gm_cxrom_1.cell10.data [6], _00358_);
  nand (_00395_, _00394_, _00393_);
  nand (_00396_, _00395_, _42355_);
  or (_00397_, \oc8051_gm_cxrom_1.cell10.data [6], _42355_);
  and (_05624_, _00397_, _00396_);
  or (_00398_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_00399_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_00400_, _00399_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_00401_, _00400_, _00398_);
  nand (_00402_, _00401_, _42355_);
  or (_00403_, \oc8051_gm_cxrom_1.cell11.data [7], _42355_);
  and (_05646_, _00403_, _00402_);
  or (_00404_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00405_, \oc8051_gm_cxrom_1.cell11.data [0], _00399_);
  nand (_00406_, _00405_, _00404_);
  nand (_00407_, _00406_, _42355_);
  or (_00408_, \oc8051_gm_cxrom_1.cell11.data [0], _42355_);
  and (_05653_, _00408_, _00407_);
  or (_00409_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00410_, \oc8051_gm_cxrom_1.cell11.data [1], _00399_);
  nand (_00411_, _00410_, _00409_);
  nand (_00412_, _00411_, _42355_);
  or (_00413_, \oc8051_gm_cxrom_1.cell11.data [1], _42355_);
  and (_05657_, _00413_, _00412_);
  or (_00414_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00415_, \oc8051_gm_cxrom_1.cell11.data [2], _00399_);
  nand (_00416_, _00415_, _00414_);
  nand (_00417_, _00416_, _42355_);
  or (_00418_, \oc8051_gm_cxrom_1.cell11.data [2], _42355_);
  and (_05661_, _00418_, _00417_);
  or (_00419_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00420_, \oc8051_gm_cxrom_1.cell11.data [3], _00399_);
  nand (_00421_, _00420_, _00419_);
  nand (_00422_, _00421_, _42355_);
  or (_00423_, \oc8051_gm_cxrom_1.cell11.data [3], _42355_);
  and (_05665_, _00423_, _00422_);
  or (_00424_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00425_, \oc8051_gm_cxrom_1.cell11.data [4], _00399_);
  nand (_00426_, _00425_, _00424_);
  nand (_00427_, _00426_, _42355_);
  or (_00428_, \oc8051_gm_cxrom_1.cell11.data [4], _42355_);
  and (_05669_, _00428_, _00427_);
  or (_00429_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00430_, \oc8051_gm_cxrom_1.cell11.data [5], _00399_);
  nand (_00431_, _00430_, _00429_);
  nand (_00432_, _00431_, _42355_);
  or (_00433_, \oc8051_gm_cxrom_1.cell11.data [5], _42355_);
  and (_05673_, _00433_, _00432_);
  or (_00434_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_00435_, \oc8051_gm_cxrom_1.cell11.data [6], _00399_);
  nand (_00436_, _00435_, _00434_);
  nand (_00437_, _00436_, _42355_);
  or (_00438_, \oc8051_gm_cxrom_1.cell11.data [6], _42355_);
  and (_05677_, _00438_, _00437_);
  or (_00439_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_00440_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_00441_, _00440_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_00442_, _00441_, _00439_);
  nand (_00443_, _00442_, _42355_);
  or (_00444_, \oc8051_gm_cxrom_1.cell12.data [7], _42355_);
  and (_05699_, _00444_, _00443_);
  or (_00445_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00446_, \oc8051_gm_cxrom_1.cell12.data [0], _00440_);
  nand (_00447_, _00446_, _00445_);
  nand (_00448_, _00447_, _42355_);
  or (_00449_, \oc8051_gm_cxrom_1.cell12.data [0], _42355_);
  and (_05706_, _00449_, _00448_);
  or (_00450_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00451_, \oc8051_gm_cxrom_1.cell12.data [1], _00440_);
  nand (_00452_, _00451_, _00450_);
  nand (_00453_, _00452_, _42355_);
  or (_00454_, \oc8051_gm_cxrom_1.cell12.data [1], _42355_);
  and (_05710_, _00454_, _00453_);
  or (_00455_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00456_, \oc8051_gm_cxrom_1.cell12.data [2], _00440_);
  nand (_00457_, _00456_, _00455_);
  nand (_00458_, _00457_, _42355_);
  or (_00459_, \oc8051_gm_cxrom_1.cell12.data [2], _42355_);
  and (_05714_, _00459_, _00458_);
  or (_00460_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00461_, \oc8051_gm_cxrom_1.cell12.data [3], _00440_);
  nand (_00462_, _00461_, _00460_);
  nand (_00463_, _00462_, _42355_);
  or (_00464_, \oc8051_gm_cxrom_1.cell12.data [3], _42355_);
  and (_05718_, _00464_, _00463_);
  or (_00465_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00466_, \oc8051_gm_cxrom_1.cell12.data [4], _00440_);
  nand (_00467_, _00466_, _00465_);
  nand (_00468_, _00467_, _42355_);
  or (_00469_, \oc8051_gm_cxrom_1.cell12.data [4], _42355_);
  and (_05722_, _00469_, _00468_);
  or (_00470_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00471_, \oc8051_gm_cxrom_1.cell12.data [5], _00440_);
  nand (_00472_, _00471_, _00470_);
  nand (_00473_, _00472_, _42355_);
  or (_00474_, \oc8051_gm_cxrom_1.cell12.data [5], _42355_);
  and (_05726_, _00474_, _00473_);
  or (_00475_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_00476_, \oc8051_gm_cxrom_1.cell12.data [6], _00440_);
  nand (_00477_, _00476_, _00475_);
  nand (_00478_, _00477_, _42355_);
  or (_00479_, \oc8051_gm_cxrom_1.cell12.data [6], _42355_);
  and (_05730_, _00479_, _00478_);
  or (_00480_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_00481_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_00482_, _00481_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_00483_, _00482_, _00480_);
  nand (_00484_, _00483_, _42355_);
  or (_00485_, \oc8051_gm_cxrom_1.cell13.data [7], _42355_);
  and (_05752_, _00485_, _00484_);
  or (_00486_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00487_, \oc8051_gm_cxrom_1.cell13.data [0], _00481_);
  nand (_00488_, _00487_, _00486_);
  nand (_00489_, _00488_, _42355_);
  or (_00490_, \oc8051_gm_cxrom_1.cell13.data [0], _42355_);
  and (_05759_, _00490_, _00489_);
  or (_00491_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00492_, \oc8051_gm_cxrom_1.cell13.data [1], _00481_);
  nand (_00493_, _00492_, _00491_);
  nand (_00494_, _00493_, _42355_);
  or (_00495_, \oc8051_gm_cxrom_1.cell13.data [1], _42355_);
  and (_05763_, _00495_, _00494_);
  or (_00496_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00497_, \oc8051_gm_cxrom_1.cell13.data [2], _00481_);
  nand (_00498_, _00497_, _00496_);
  nand (_00499_, _00498_, _42355_);
  or (_00500_, \oc8051_gm_cxrom_1.cell13.data [2], _42355_);
  and (_05767_, _00500_, _00499_);
  or (_00501_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00502_, \oc8051_gm_cxrom_1.cell13.data [3], _00481_);
  nand (_00503_, _00502_, _00501_);
  nand (_00504_, _00503_, _42355_);
  or (_00505_, \oc8051_gm_cxrom_1.cell13.data [3], _42355_);
  and (_05771_, _00505_, _00504_);
  or (_00506_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00507_, \oc8051_gm_cxrom_1.cell13.data [4], _00481_);
  nand (_00508_, _00507_, _00506_);
  nand (_00509_, _00508_, _42355_);
  or (_00510_, \oc8051_gm_cxrom_1.cell13.data [4], _42355_);
  and (_05775_, _00510_, _00509_);
  or (_00511_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00512_, \oc8051_gm_cxrom_1.cell13.data [5], _00481_);
  nand (_00513_, _00512_, _00511_);
  nand (_00514_, _00513_, _42355_);
  or (_00515_, \oc8051_gm_cxrom_1.cell13.data [5], _42355_);
  and (_05779_, _00515_, _00514_);
  or (_00516_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_00517_, \oc8051_gm_cxrom_1.cell13.data [6], _00481_);
  nand (_00518_, _00517_, _00516_);
  nand (_00519_, _00518_, _42355_);
  or (_00520_, \oc8051_gm_cxrom_1.cell13.data [6], _42355_);
  and (_05783_, _00520_, _00519_);
  or (_00521_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_00522_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_00523_, _00522_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_00524_, _00523_, _00521_);
  nand (_00525_, _00524_, _42355_);
  or (_00526_, \oc8051_gm_cxrom_1.cell14.data [7], _42355_);
  and (_05805_, _00526_, _00525_);
  or (_00527_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00528_, \oc8051_gm_cxrom_1.cell14.data [0], _00522_);
  nand (_00529_, _00528_, _00527_);
  nand (_00530_, _00529_, _42355_);
  or (_00531_, \oc8051_gm_cxrom_1.cell14.data [0], _42355_);
  and (_05812_, _00531_, _00530_);
  or (_00532_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00533_, \oc8051_gm_cxrom_1.cell14.data [1], _00522_);
  nand (_00534_, _00533_, _00532_);
  nand (_00535_, _00534_, _42355_);
  or (_00536_, \oc8051_gm_cxrom_1.cell14.data [1], _42355_);
  and (_05816_, _00536_, _00535_);
  or (_00537_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00538_, \oc8051_gm_cxrom_1.cell14.data [2], _00522_);
  nand (_00539_, _00538_, _00537_);
  nand (_00540_, _00539_, _42355_);
  or (_00541_, \oc8051_gm_cxrom_1.cell14.data [2], _42355_);
  and (_05820_, _00541_, _00540_);
  or (_00542_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00544_, \oc8051_gm_cxrom_1.cell14.data [3], _00522_);
  nand (_00545_, _00544_, _00542_);
  nand (_00547_, _00545_, _42355_);
  or (_00548_, \oc8051_gm_cxrom_1.cell14.data [3], _42355_);
  and (_05824_, _00548_, _00547_);
  or (_00550_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00552_, \oc8051_gm_cxrom_1.cell14.data [4], _00522_);
  nand (_00553_, _00552_, _00550_);
  nand (_00555_, _00553_, _42355_);
  or (_00556_, \oc8051_gm_cxrom_1.cell14.data [4], _42355_);
  and (_05828_, _00556_, _00555_);
  or (_00558_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00560_, \oc8051_gm_cxrom_1.cell14.data [5], _00522_);
  nand (_00561_, _00560_, _00558_);
  nand (_00563_, _00561_, _42355_);
  or (_00564_, \oc8051_gm_cxrom_1.cell14.data [5], _42355_);
  and (_05832_, _00564_, _00563_);
  or (_00566_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_00568_, \oc8051_gm_cxrom_1.cell14.data [6], _00522_);
  nand (_00569_, _00568_, _00566_);
  nand (_00571_, _00569_, _42355_);
  or (_00572_, \oc8051_gm_cxrom_1.cell14.data [6], _42355_);
  and (_05836_, _00572_, _00571_);
  or (_00574_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_00576_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_00577_, _00576_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_00579_, _00577_, _00574_);
  nand (_00580_, _00579_, _42355_);
  or (_00582_, \oc8051_gm_cxrom_1.cell15.data [7], _42355_);
  and (_05858_, _00582_, _00580_);
  or (_00584_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00585_, \oc8051_gm_cxrom_1.cell15.data [0], _00576_);
  nand (_00587_, _00585_, _00584_);
  nand (_00588_, _00587_, _42355_);
  or (_00590_, \oc8051_gm_cxrom_1.cell15.data [0], _42355_);
  and (_05865_, _00590_, _00588_);
  or (_00592_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00593_, \oc8051_gm_cxrom_1.cell15.data [1], _00576_);
  nand (_00594_, _00593_, _00592_);
  nand (_00595_, _00594_, _42355_);
  or (_00596_, \oc8051_gm_cxrom_1.cell15.data [1], _42355_);
  and (_05869_, _00596_, _00595_);
  or (_00597_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00598_, \oc8051_gm_cxrom_1.cell15.data [2], _00576_);
  nand (_00599_, _00598_, _00597_);
  nand (_00600_, _00599_, _42355_);
  or (_00601_, \oc8051_gm_cxrom_1.cell15.data [2], _42355_);
  and (_05873_, _00601_, _00600_);
  or (_00602_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00603_, \oc8051_gm_cxrom_1.cell15.data [3], _00576_);
  nand (_00604_, _00603_, _00602_);
  nand (_00605_, _00604_, _42355_);
  or (_00606_, \oc8051_gm_cxrom_1.cell15.data [3], _42355_);
  and (_05877_, _00606_, _00605_);
  or (_00607_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00608_, \oc8051_gm_cxrom_1.cell15.data [4], _00576_);
  nand (_00609_, _00608_, _00607_);
  nand (_00610_, _00609_, _42355_);
  or (_00611_, \oc8051_gm_cxrom_1.cell15.data [4], _42355_);
  and (_05881_, _00611_, _00610_);
  or (_00612_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00613_, \oc8051_gm_cxrom_1.cell15.data [5], _00576_);
  nand (_00614_, _00613_, _00612_);
  nand (_00615_, _00614_, _42355_);
  or (_00616_, \oc8051_gm_cxrom_1.cell15.data [5], _42355_);
  and (_05885_, _00616_, _00615_);
  or (_00617_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_00618_, \oc8051_gm_cxrom_1.cell15.data [6], _00576_);
  nand (_00619_, _00618_, _00617_);
  nand (_00620_, _00619_, _42355_);
  or (_00621_, \oc8051_gm_cxrom_1.cell15.data [6], _42355_);
  and (_05889_, _00621_, _00620_);
  nor (_09664_, _37738_, rst);
  and (_00622_, _37025_, _42355_);
  nand (_00623_, _00622_, _37797_);
  nor (_00624_, _37724_, _37704_);
  or (_09667_, _00624_, _00623_);
  and (_00625_, _37652_, _37675_);
  and (_00626_, _00625_, _37697_);
  and (_00627_, _00626_, _37628_);
  and (_00628_, _37603_, _37556_);
  and (_00629_, _37579_, _37429_);
  and (_00630_, _00629_, _00628_);
  and (_00631_, _00630_, _00627_);
  not (_00632_, _37628_);
  nor (_00633_, _37579_, _37429_);
  not (_00634_, _37603_);
  and (_00635_, _00634_, _37556_);
  and (_00636_, _00635_, _00633_);
  nor (_00637_, _00636_, _00632_);
  not (_00638_, _37652_);
  and (_00639_, _37697_, _37675_);
  and (_00640_, _00639_, _00638_);
  not (_00641_, _00640_);
  nor (_00642_, _00641_, _00637_);
  not (_00643_, _00642_);
  and (_00644_, _37628_, _00638_);
  and (_00645_, _00644_, _00639_);
  not (_00646_, _37579_);
  and (_00647_, _00646_, _37429_);
  and (_00648_, _00647_, _00628_);
  and (_00649_, _00648_, _00645_);
  not (_00650_, _37429_);
  and (_00651_, _37579_, _00650_);
  and (_00652_, _00651_, _00635_);
  and (_00653_, _00652_, _00645_);
  nor (_00654_, _00653_, _00649_);
  and (_00655_, _00654_, _00643_);
  nor (_00656_, _37603_, _37556_);
  and (_00657_, _00656_, _00646_);
  and (_00658_, _37429_, _37697_);
  and (_00659_, _00658_, _00625_);
  and (_00660_, _00659_, _00657_);
  not (_00661_, _37697_);
  and (_00662_, _00656_, _00629_);
  and (_00663_, _00662_, _00661_);
  nor (_00664_, _00661_, _37675_);
  and (_00665_, _00664_, _00638_);
  not (_00666_, _37556_);
  and (_00667_, _37603_, _00666_);
  and (_00668_, _00667_, _00647_);
  and (_00669_, _00668_, _00665_);
  or (_00670_, _00669_, _00663_);
  nor (_00671_, _00670_, _00660_);
  nand (_00672_, _00671_, _00655_);
  or (_00673_, _00672_, _00631_);
  nor (_00674_, _00651_, _00647_);
  and (_00675_, _00645_, _00628_);
  and (_00676_, _00675_, _00674_);
  and (_00677_, _00664_, _00644_);
  and (_00678_, _00677_, _00650_);
  and (_00679_, _00678_, _00667_);
  and (_00680_, _00627_, _00628_);
  not (_00681_, _00629_);
  and (_00682_, _00681_, _00680_);
  or (_00683_, _00682_, _00679_);
  or (_00684_, _00683_, _00676_);
  and (_00685_, _00650_, _37697_);
  and (_00686_, _00685_, _00625_);
  and (_00687_, _00686_, _00657_);
  and (_00688_, _00665_, _00632_);
  and (_00689_, _00688_, _00662_);
  or (_00690_, _00689_, _00687_);
  nor (_00691_, _00638_, _37675_);
  nor (_00692_, _00691_, _00661_);
  not (_00693_, _00692_);
  and (_00694_, _00693_, _00668_);
  and (_00695_, _00657_, _00645_);
  or (_00696_, _00695_, _00694_);
  or (_00697_, _00696_, _00690_);
  and (_00698_, _00667_, _37579_);
  and (_00699_, _00626_, _00632_);
  and (_00700_, _00699_, _00698_);
  and (_00701_, _00635_, _37429_);
  and (_00702_, _00701_, _00645_);
  or (_00703_, _00702_, _00700_);
  and (_00704_, _00647_, _00635_);
  and (_00705_, _00704_, _00699_);
  and (_00706_, _00667_, _00651_);
  and (_00707_, _00706_, _00645_);
  or (_00708_, _00707_, _00705_);
  or (_00709_, _00708_, _00703_);
  or (_00710_, _00709_, _00697_);
  or (_00711_, _00710_, _00684_);
  or (_00712_, _00711_, _00673_);
  and (_00713_, _00712_, _37036_);
  not (_00714_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_00715_, _37014_, _18787_);
  and (_00716_, _00715_, _37720_);
  nor (_00717_, _00716_, _00714_);
  or (_00718_, _00717_, rst);
  or (_09670_, _00718_, _00713_);
  nand (_00719_, _37556_, _36960_);
  or (_00720_, _36960_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_00721_, _00720_, _42355_);
  and (_09673_, _00721_, _00719_);
  and (_00722_, \oc8051_top_1.oc8051_sfr1.wait_data , _42355_);
  and (_00723_, _00722_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00724_, _37732_, _37798_);
  and (_00725_, _37705_, _37714_);
  and (_00726_, _00725_, _37505_);
  or (_00727_, _00726_, _00724_);
  and (_00728_, _37729_, _37724_);
  or (_00729_, _00728_, _37726_);
  or (_00730_, _00729_, _37757_);
  and (_00731_, _37765_, _37704_);
  and (_00732_, _37705_, _37756_);
  or (_00733_, _00732_, _00731_);
  nor (_00734_, _00733_, _00730_);
  nand (_00735_, _00734_, _37790_);
  or (_00736_, _00735_, _00727_);
  and (_00737_, _00736_, _00622_);
  or (_09676_, _00737_, _00723_);
  and (_00738_, _37505_, _37702_);
  and (_00739_, _00738_, _37755_);
  or (_00740_, _00739_, _37859_);
  and (_00741_, _37742_, _37731_);
  and (_00742_, _00741_, _37756_);
  or (_00743_, _00742_, _00740_);
  and (_00744_, _37715_, _37724_);
  or (_00745_, _00744_, _37706_);
  or (_00746_, _00745_, _00743_);
  and (_00747_, _00746_, _37025_);
  and (_00748_, _37833_, _00714_);
  not (_00749_, _37735_);
  and (_00750_, _00749_, _00748_);
  and (_00751_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00752_, _00751_, _00750_);
  or (_00753_, _00752_, _00747_);
  and (_09679_, _00753_, _42355_);
  and (_00754_, _00722_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_00755_, _37732_, _37815_);
  nor (_00756_, _37815_, _37765_);
  nor (_00757_, _00756_, _37809_);
  or (_00758_, _00757_, _00755_);
  and (_00759_, _00741_, _37747_);
  or (_00760_, _00759_, _00758_);
  nor (_00761_, _00756_, _37730_);
  and (_00762_, _37495_, _37702_);
  and (_00763_, _00762_, _37746_);
  or (_00764_, _00763_, _00761_);
  or (_00765_, _00764_, _37851_);
  and (_00766_, _37732_, _37805_);
  and (_00767_, _37752_, _37702_);
  or (_00768_, _00767_, _00766_);
  or (_00769_, _00768_, _00745_);
  or (_00770_, _00769_, _00765_);
  or (_00771_, _00770_, _00760_);
  and (_00772_, _00771_, _00622_);
  or (_09682_, _00772_, _00754_);
  and (_00773_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00774_, _37779_, _37025_);
  or (_00775_, _00774_, _00773_);
  or (_00776_, _00775_, _00750_);
  and (_09685_, _00776_, _42355_);
  and (_00777_, _37751_, _37747_);
  and (_00778_, _37703_, _37743_);
  and (_00779_, _00778_, _37495_);
  or (_00780_, _00779_, _00777_);
  or (_00781_, _00780_, _00726_);
  and (_00782_, _00780_, _37722_);
  or (_00783_, _00782_, _36971_);
  and (_00784_, _00783_, _00781_);
  not (_00785_, _37798_);
  nor (_00786_, _00624_, _00785_);
  nor (_00787_, _00786_, _00725_);
  not (_00788_, _00787_);
  and (_00789_, _00788_, _00748_);
  or (_00790_, _00789_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00791_, _00790_, _00784_);
  or (_00792_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18787_);
  and (_00793_, _00792_, _42355_);
  and (_09688_, _00793_, _00791_);
  and (_00794_, _00722_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_00795_, _00763_, _37706_);
  and (_00796_, _00762_, _37755_);
  or (_00797_, _00796_, _37766_);
  or (_00798_, _00797_, _00795_);
  and (_00799_, _37609_, _37751_);
  or (_00800_, _00759_, _00731_);
  or (_00801_, _00800_, _00799_);
  or (_00802_, _37756_, _37747_);
  and (_00803_, _00802_, _37802_);
  or (_00804_, _00739_, _37822_);
  or (_00805_, _00804_, _00803_);
  or (_00806_, _00805_, _00801_);
  or (_00807_, _00806_, _00798_);
  and (_00808_, _00807_, _00622_);
  or (_09691_, _00808_, _00794_);
  and (_00809_, _00722_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_00810_, _00741_, _37792_);
  and (_00811_, _37705_, _37745_);
  or (_00812_, _00811_, _00742_);
  or (_00813_, _00812_, _00810_);
  or (_00814_, _00813_, _00764_);
  nand (_00815_, _37732_, _37762_);
  nand (_00816_, _00815_, _37770_);
  and (_00817_, _37803_, _37754_);
  or (_00818_, _00817_, _37863_);
  and (_00819_, _37802_, _37765_);
  or (_00820_, _00819_, _00818_);
  or (_00821_, _00820_, _00816_);
  or (_00822_, _00821_, _00814_);
  and (_00823_, _00738_, _37754_);
  and (_00824_, _00738_, _37710_);
  or (_00825_, _00824_, _00823_);
  nor (_00826_, _37850_, _37793_);
  nand (_00827_, _00826_, _37764_);
  or (_00828_, _00827_, _00825_);
  or (_00829_, _00828_, _00760_);
  or (_00830_, _00829_, _00822_);
  and (_00831_, _00830_, _00622_);
  or (_09694_, _00831_, _00809_);
  and (_00832_, _00741_, _37782_);
  or (_00833_, _00832_, _37860_);
  and (_00834_, _00762_, _37713_);
  and (_00835_, _00834_, _37561_);
  or (_00836_, _00835_, _37844_);
  and (_00837_, _37782_, _37702_);
  or (_00838_, _00837_, _00836_);
  or (_00839_, _00838_, _00833_);
  and (_00840_, _00741_, _37715_);
  or (_00841_, _00840_, _00749_);
  or (_00842_, _00841_, _00839_);
  and (_00843_, _00842_, _00622_);
  nor (_00844_, _37735_, _36971_);
  and (_00845_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_00846_, _00845_, _00844_);
  and (_00847_, _00846_, _42355_);
  or (_09697_, _00847_, _00843_);
  nand (_00848_, _37794_, _37780_);
  or (_00849_, _37824_, _37822_);
  or (_00850_, _00849_, _00757_);
  or (_00851_, _00850_, _00848_);
  and (_00852_, _37709_, _37495_);
  and (_00853_, _00852_, _37744_);
  or (_00854_, _00853_, _37769_);
  or (_00855_, _00854_, _00777_);
  or (_00856_, _00855_, _37759_);
  or (_00857_, _00856_, _00851_);
  and (_00858_, _00738_, _37714_);
  or (_00859_, _00858_, _37847_);
  or (_00860_, _00859_, _00779_);
  or (_00861_, _00860_, _37776_);
  and (_00862_, _00852_, _37802_);
  or (_00863_, _00862_, _37850_);
  or (_00864_, _00863_, _37804_);
  and (_00865_, _00762_, _37709_);
  or (_00866_, _00865_, _37817_);
  or (_00867_, _00866_, _00740_);
  or (_00868_, _00867_, _00864_);
  or (_00869_, _00868_, _00764_);
  or (_00870_, _00869_, _00861_);
  or (_00871_, _00870_, _00857_);
  and (_00872_, _00871_, _37025_);
  or (_00873_, _00782_, _00750_);
  and (_00874_, _37722_, _37788_);
  or (_00875_, _00874_, _00873_);
  and (_00876_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00877_, _00876_, _00875_);
  or (_00878_, _00877_, _00872_);
  and (_09700_, _00878_, _42355_);
  nor (_09759_, _37872_, rst);
  nor (_09761_, _37837_, rst);
  nand (_09764_, _00788_, _00622_);
  nand (_00879_, _00725_, _00622_);
  not (_00880_, _37724_);
  or (_00881_, _00623_, _00880_);
  and (_09767_, _00881_, _00879_);
  and (_00882_, _00680_, _00646_);
  or (_00883_, _00700_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_00884_, _00883_, _00679_);
  or (_00885_, _00884_, _00882_);
  and (_00886_, _00885_, _00716_);
  nor (_00887_, _00715_, _37720_);
  or (_00888_, _00887_, rst);
  or (_09770_, _00888_, _00886_);
  nand (_00889_, _37628_, _36960_);
  or (_00890_, _36960_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_00891_, _00890_, _42355_);
  and (_09773_, _00891_, _00889_);
  not (_00892_, _36960_);
  or (_00893_, _37652_, _00892_);
  or (_00894_, _36960_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_00895_, _00894_, _42355_);
  and (_09776_, _00895_, _00893_);
  nand (_00896_, _37675_, _36960_);
  or (_00897_, _36960_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_00898_, _00897_, _42355_);
  and (_09779_, _00898_, _00896_);
  nand (_00899_, _37697_, _36960_);
  or (_00900_, _36960_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_00901_, _00900_, _42355_);
  and (_09782_, _00901_, _00899_);
  or (_00902_, _37429_, _00892_);
  or (_00903_, _36960_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_00904_, _00903_, _42355_);
  and (_09785_, _00904_, _00902_);
  nand (_00905_, _37579_, _36960_);
  or (_00906_, _36960_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_00907_, _00906_, _42355_);
  and (_09788_, _00907_, _00905_);
  nand (_00908_, _37603_, _36960_);
  or (_00909_, _36960_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_00910_, _00909_, _42355_);
  and (_09791_, _00910_, _00908_);
  or (_00911_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _18787_);
  and (_00912_, _00911_, _42355_);
  and (_00913_, _00912_, _00790_);
  and (_00914_, _00741_, _37762_);
  or (_00915_, _00914_, _00744_);
  and (_00916_, _37802_, _37715_);
  or (_00917_, _00832_, _00916_);
  and (_00918_, _00738_, _37761_);
  or (_00919_, _00840_, _00918_);
  or (_00920_, _00919_, _00917_);
  or (_00921_, _37706_, _37853_);
  or (_00922_, _00921_, _00920_);
  or (_00923_, _00922_, _00915_);
  and (_00924_, _00741_, _37775_);
  and (_00926_, _37802_, _37775_);
  or (_00927_, _00926_, _00924_);
  and (_00928_, _00738_, _37797_);
  and (_00929_, _00741_, _37798_);
  or (_00930_, _00929_, _00928_);
  or (_00931_, _00930_, _00927_);
  or (_00932_, _00824_, _37863_);
  or (_00933_, _00836_, _00810_);
  or (_00934_, _00933_, _00932_);
  or (_00935_, _00934_, _00931_);
  or (_00936_, _37765_, _37746_);
  or (_00937_, _00936_, _00852_);
  and (_00938_, _00937_, _37732_);
  and (_00939_, _37761_, _37702_);
  and (_00940_, _00939_, _37495_);
  or (_00941_, _00940_, _00837_);
  or (_00942_, _00941_, _00811_);
  or (_00943_, _00942_, _00938_);
  or (_00944_, _00943_, _00935_);
  or (_00945_, _00944_, _00923_);
  and (_00946_, _00945_, _00622_);
  or (_09794_, _00946_, _00913_);
  and (_00947_, _00722_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_00948_, _37792_, _37762_);
  and (_00949_, _00948_, _37751_);
  or (_00950_, _00915_, _00825_);
  or (_00951_, _00950_, _00949_);
  and (_00952_, _00762_, _37608_);
  and (_00953_, _00952_, _37561_);
  nor (_00954_, _00953_, _37849_);
  not (_00956_, _00954_);
  nor (_00957_, _00956_, _00766_);
  nand (_00958_, _00957_, _37823_);
  or (_00959_, _00958_, _00727_);
  not (_00960_, _37792_);
  nand (_00961_, _37810_, _00960_);
  and (_00962_, _00961_, _37732_);
  or (_00963_, _00962_, _00820_);
  or (_00964_, _00963_, _00959_);
  or (_00965_, _00964_, _00951_);
  and (_00966_, _00965_, _00622_);
  or (_34183_, _00966_, _00947_);
  or (_00967_, _00861_, _00857_);
  and (_00968_, _00967_, _37025_);
  and (_00969_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00970_, _00969_, _00875_);
  or (_00971_, _00970_, _00968_);
  and (_34185_, _00971_, _42355_);
  and (_00972_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00973_, _00972_, _00873_);
  and (_00975_, _00973_, _42355_);
  and (_00976_, _37791_, _37505_);
  or (_00977_, _00976_, _37859_);
  or (_00978_, _00977_, _00864_);
  or (_00979_, _00978_, _00780_);
  and (_00980_, _00979_, _00622_);
  or (_34188_, _00980_, _00975_);
  or (_00981_, _00836_, _37843_);
  or (_00982_, _00948_, _37711_);
  and (_00983_, _00982_, _37732_);
  or (_00984_, _00725_, _37734_);
  and (_00985_, _00832_, _37495_);
  or (_00986_, _00985_, _00924_);
  or (_00987_, _00986_, _00984_);
  or (_00988_, _00987_, _00983_);
  or (_00989_, _00988_, _00981_);
  or (_00990_, _00936_, _37756_);
  and (_00991_, _00990_, _37732_);
  and (_00992_, _37797_, _37495_);
  and (_00993_, _00992_, _37732_);
  or (_00994_, _00993_, _37733_);
  and (_00995_, _00741_, _37752_);
  or (_00996_, _00995_, _00840_);
  or (_00997_, _00996_, _00724_);
  or (_00998_, _00997_, _00994_);
  or (_00999_, _00998_, _00991_);
  and (_01000_, _00832_, _37505_);
  or (_01001_, _01000_, _37712_);
  or (_01002_, _00865_, _00916_);
  or (_01003_, _01002_, _00862_);
  and (_01004_, _00992_, _37744_);
  and (_01005_, _37775_, _37751_);
  or (_01006_, _01005_, _01004_);
  or (_01007_, _01006_, _01003_);
  or (_01008_, _01007_, _01001_);
  or (_01009_, _00942_, _00780_);
  or (_01010_, _01009_, _01008_);
  or (_01011_, _01010_, _00999_);
  or (_01012_, _01011_, _00989_);
  and (_01013_, _01012_, _37025_);
  and (_01014_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01015_, _00789_, _00844_);
  or (_01016_, _01015_, _01014_);
  or (_01017_, _01016_, _01013_);
  and (_34190_, _01017_, _42355_);
  and (_01018_, _00992_, _37802_);
  or (_01019_, _37734_, _00916_);
  or (_01020_, _01019_, _37776_);
  or (_01021_, _01020_, _01018_);
  or (_01022_, _01021_, _00942_);
  or (_01023_, _01022_, _00981_);
  and (_01024_, _00762_, _37797_);
  or (_01025_, _00853_, _00744_);
  nor (_01026_, _01025_, _01024_);
  nand (_01027_, _01026_, _37717_);
  and (_01028_, _00948_, _37705_);
  or (_01029_, _01028_, _37811_);
  or (_01030_, _01029_, _01027_);
  or (_01031_, _01030_, _00999_);
  or (_01032_, _01031_, _01023_);
  and (_01033_, _01032_, _37025_);
  and (_01034_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01035_, _01034_, _01015_);
  or (_01036_, _01035_, _01033_);
  and (_34192_, _01036_, _42355_);
  and (_01037_, _00722_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_01038_, _41835_);
  or (_01039_, _00840_, _01038_);
  or (_01040_, _01039_, _00798_);
  and (_01041_, _37705_, _37746_);
  and (_01042_, _01041_, _37495_);
  and (_01043_, _00731_, _37633_);
  or (_01044_, _01043_, _01042_);
  or (_01045_, _01044_, _01040_);
  not (_01046_, _41833_);
  or (_01047_, _00803_, _01046_);
  and (_01048_, _37732_, _37765_);
  or (_01049_, _01048_, _00759_);
  or (_01050_, _01049_, _00849_);
  or (_01051_, _01050_, _01047_);
  and (_01052_, _37842_, _37782_);
  or (_01053_, _00835_, _00739_);
  and (_01054_, _37705_, _37752_);
  or (_01055_, _01054_, _01053_);
  or (_01056_, _01055_, _01052_);
  and (_01057_, _00952_, _37708_);
  or (_01058_, _01057_, _00916_);
  or (_01059_, _01058_, _37778_);
  and (_01060_, _37705_, _37783_);
  or (_01061_, _01060_, _00985_);
  or (_01062_, _01061_, _01059_);
  or (_01063_, _01062_, _01056_);
  or (_01064_, _01063_, _01051_);
  or (_01065_, _01064_, _01045_);
  and (_01066_, _01065_, _00622_);
  or (_34194_, _01066_, _01037_);
  or (_01067_, _00742_, _37763_);
  or (_01068_, _00819_, _00817_);
  or (_01069_, _01068_, _01067_);
  or (_01070_, _01069_, _00816_);
  or (_01071_, _01070_, _00987_);
  or (_01072_, _01060_, _01048_);
  or (_01073_, _01042_, _01001_);
  or (_01074_, _01073_, _01072_);
  or (_01075_, _00823_, _37706_);
  or (_01076_, _01075_, _37845_);
  not (_01077_, _37777_);
  or (_01078_, _00941_, _01077_);
  or (_01079_, _01078_, _01076_);
  or (_01080_, _01079_, _01074_);
  or (_01081_, _01080_, _01071_);
  and (_01082_, _01081_, _00622_);
  and (_01083_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01084_, _37734_, _36982_);
  or (_01085_, _01084_, _01083_);
  and (_01086_, _01085_, _42355_);
  or (_34196_, _01086_, _01082_);
  or (_01087_, _00767_, _37862_);
  or (_01088_, _01087_, _00997_);
  or (_01089_, _00940_, _00926_);
  and (_01090_, _37752_, _37704_);
  or (_01091_, _01090_, _00993_);
  or (_01092_, _01091_, _01089_);
  or (_01093_, _01092_, _01088_);
  or (_01094_, _00924_, _37776_);
  or (_01095_, _01094_, _37774_);
  or (_01096_, _00742_, _41832_);
  and (_01097_, _37705_, _37782_);
  or (_01098_, _01097_, _01053_);
  or (_01099_, _01098_, _01096_);
  or (_01100_, _01099_, _01095_);
  or (_01101_, _01100_, _01093_);
  or (_01102_, _00765_, _00760_);
  or (_01103_, _01102_, _01101_);
  and (_01104_, _01103_, _37025_);
  and (_01105_, _37734_, _18787_);
  and (_01106_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01107_, _01106_, _01105_);
  or (_01108_, _01107_, _01104_);
  and (_34198_, _01108_, _42355_);
  or (_01109_, _37733_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_01110_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18787_);
  and (_01111_, _01110_, _42355_);
  and (_01112_, _01111_, _01109_);
  or (_01113_, _01094_, _01092_);
  or (_01114_, _37859_, _37850_);
  nor (_01115_, _01114_, _01041_);
  nand (_01116_, _01115_, _41835_);
  or (_01117_, _01049_, _00804_);
  or (_01118_, _01117_, _01116_);
  or (_01119_, _00764_, _00758_);
  or (_01120_, _01119_, _01118_);
  or (_01121_, _01120_, _01113_);
  and (_01122_, _01121_, _00622_);
  or (_34200_, _01122_, _01112_);
  and (_01123_, _00722_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_01124_, _00732_, _37825_);
  nand (_01125_, _01124_, _41833_);
  not (_01126_, _37703_);
  or (_01127_, _37705_, _01126_);
  and (_01128_, _01127_, _37752_);
  or (_01129_, _01128_, _01072_);
  or (_01130_, _01129_, _01125_);
  or (_01131_, _01039_, _00839_);
  or (_01132_, _01131_, _01044_);
  or (_01133_, _01132_, _01130_);
  and (_01134_, _01133_, _00622_);
  or (_34202_, _01134_, _01123_);
  nor (_38381_, _37556_, rst);
  nor (_38382_, _41767_, rst);
  and (_01135_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_01136_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_01137_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01138_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_01139_, _01138_, _01137_);
  and (_01140_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_01141_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_01142_, _01141_, _01140_);
  and (_01143_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_01144_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_01145_, _01144_, _01143_);
  and (_01146_, _01145_, _01142_);
  and (_01147_, _01146_, _01139_);
  nor (_01148_, _01147_, _37156_);
  nor (_01149_, _01148_, _01136_);
  nor (_01150_, _01149_, _41751_);
  nor (_01151_, _01150_, _01135_);
  nor (_38384_, _01151_, rst);
  nor (_38395_, _37628_, rst);
  and (_38397_, _37652_, _42355_);
  nor (_38398_, _37675_, rst);
  nor (_38399_, _37697_, rst);
  and (_38400_, _37429_, _42355_);
  nor (_38401_, _37579_, rst);
  nor (_38402_, _37603_, rst);
  nor (_38403_, _42011_, rst);
  nor (_38404_, _41933_, rst);
  nor (_38406_, _42154_, rst);
  nor (_38407_, _41968_, rst);
  nor (_38408_, _41864_, rst);
  nor (_38409_, _42128_, rst);
  nor (_38410_, _42084_, rst);
  and (_01152_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_01153_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_01154_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_01155_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01156_, _01155_, _01154_);
  and (_01157_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_01158_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01159_, _01158_, _01157_);
  and (_01160_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01161_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_01162_, _01161_, _01160_);
  and (_01163_, _01162_, _01159_);
  and (_01164_, _01163_, _01156_);
  nor (_01165_, _01164_, _37156_);
  nor (_01166_, _01165_, _01153_);
  nor (_01167_, _01166_, _41751_);
  nor (_01168_, _01167_, _01152_);
  nor (_38412_, _01168_, rst);
  and (_01169_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_01170_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_01171_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_01172_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01173_, _01172_, _01171_);
  and (_01174_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_01175_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01176_, _01175_, _01174_);
  and (_01177_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01178_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_01179_, _01178_, _01177_);
  and (_01180_, _01179_, _01176_);
  and (_01181_, _01180_, _01173_);
  nor (_01182_, _01181_, _37156_);
  nor (_01183_, _01182_, _01170_);
  nor (_01184_, _01183_, _41751_);
  nor (_01185_, _01184_, _01169_);
  nor (_38413_, _01185_, rst);
  and (_01186_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_01187_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_01188_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_01189_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01190_, _01189_, _01188_);
  and (_01191_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_01192_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01193_, _01192_, _01191_);
  and (_01194_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_01195_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_01196_, _01195_, _01194_);
  and (_01197_, _01196_, _01193_);
  and (_01198_, _01197_, _01190_);
  nor (_01199_, _01198_, _37156_);
  nor (_01200_, _01199_, _01187_);
  nor (_01201_, _01200_, _41751_);
  nor (_01202_, _01201_, _01186_);
  nor (_38414_, _01202_, rst);
  and (_01203_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_01204_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_01205_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_01206_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01207_, _01206_, _01205_);
  and (_01208_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_01210_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01212_, _01210_, _01208_);
  and (_01214_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_01216_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_01218_, _01216_, _01214_);
  and (_01220_, _01218_, _01212_);
  and (_01222_, _01220_, _01207_);
  nor (_01224_, _01222_, _37156_);
  nor (_01226_, _01224_, _01204_);
  nor (_01228_, _01226_, _41751_);
  nor (_01230_, _01228_, _01203_);
  nor (_38415_, _01230_, rst);
  and (_01233_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_01235_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_01237_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_01239_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01241_, _01239_, _01237_);
  and (_01243_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_01245_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_01247_, _01245_, _01243_);
  and (_01249_, _01247_, _01241_);
  and (_01251_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_01253_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01255_, _01253_, _01251_);
  and (_01257_, _01255_, _01249_);
  nor (_01259_, _01257_, _37156_);
  nor (_01261_, _01259_, _01235_);
  nor (_01263_, _01261_, _41751_);
  nor (_01265_, _01263_, _01233_);
  nor (_38416_, _01265_, rst);
  and (_01268_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_01270_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_01272_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_01274_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01276_, _01274_, _01272_);
  and (_01278_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_01280_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_01282_, _01280_, _01278_);
  and (_01284_, _01282_, _01276_);
  and (_01286_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_01288_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01290_, _01288_, _01286_);
  and (_01292_, _01290_, _01284_);
  nor (_01294_, _01292_, _37156_);
  nor (_01296_, _01294_, _01270_);
  nor (_01298_, _01296_, _41751_);
  nor (_01300_, _01298_, _01268_);
  nor (_38418_, _01300_, rst);
  and (_01303_, _41751_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_01304_, _37156_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_01305_, _37309_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_01306_, _37254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01307_, _01306_, _01305_);
  and (_01308_, _37091_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_01309_, _37287_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01310_, _01309_, _01308_);
  and (_01311_, _37123_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_01312_, _37189_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_01313_, _01312_, _01311_);
  and (_01314_, _01313_, _01310_);
  and (_01315_, _01314_, _01307_);
  nor (_01316_, _01315_, _37156_);
  nor (_01317_, _01316_, _01304_);
  nor (_01318_, _01317_, _41751_);
  nor (_01319_, _01318_, _01303_);
  nor (_38419_, _01319_, rst);
  and (_01320_, _37036_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_01321_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_01322_, _01320_, _38050_);
  and (_01323_, _01322_, _42355_);
  and (_38444_, _01323_, _01321_);
  not (_01324_, _01320_);
  or (_01325_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _01320_, _42355_);
  and (_01326_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _42355_);
  or (_01327_, _01326_, _00000_);
  and (_38445_, _01327_, _01325_);
  nor (_38480_, _41829_, rst);
  and (_38483_, _41825_, _42355_);
  nor (_01328_, _41994_, _28290_);
  and (_01329_, _41994_, _28290_);
  nor (_01330_, _01329_, _01328_);
  not (_01331_, _01330_);
  nor (_01332_, _42088_, _27830_);
  and (_01333_, _42088_, _27830_);
  nor (_01334_, _01333_, _01332_);
  nor (_01335_, _01334_, _42212_);
  nor (_01336_, _42138_, _27961_);
  and (_01337_, _42138_, _27961_);
  nor (_01338_, _01337_, _01336_);
  nor (_01339_, _41894_, _28433_);
  and (_01340_, _41894_, _28433_);
  nor (_01341_, _01340_, _01339_);
  nor (_01342_, _01341_, _01338_);
  and (_01343_, _01342_, _01335_);
  and (_01344_, _01343_, _01331_);
  and (_01345_, _42037_, _33206_);
  nor (_01346_, _42037_, _33206_);
  or (_01347_, _01346_, _01345_);
  nor (_01348_, _01347_, _38681_);
  nor (_01349_, _41939_, _27490_);
  and (_01350_, _41939_, _27490_);
  nor (_01351_, _01350_, _01349_);
  nor (_01352_, _42180_, _27369_);
  and (_01353_, _42180_, _27369_);
  nor (_01354_, _01353_, _01352_);
  nor (_01355_, _01354_, _01351_);
  and (_01356_, _01355_, _01348_);
  and (_01357_, _01356_, _01344_);
  nor (_01358_, _28137_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_01359_, _01358_, _01357_);
  not (_01360_, _01359_);
  nor (_01361_, _37790_, _37833_);
  nor (_01362_, _31922_, _39283_);
  and (_01363_, _01362_, _01344_);
  and (_01364_, _01363_, _01361_);
  and (_01365_, _37751_, _37746_);
  nor (_01366_, _01365_, _00778_);
  nor (_01367_, _01366_, _36982_);
  nor (_01368_, _37742_, _37679_);
  and (_01369_, _37633_, _37730_);
  and (_01370_, _01369_, _01368_);
  and (_01371_, _01370_, _37711_);
  nor (_01372_, _01371_, _00728_);
  or (_01373_, _34174_, _32073_);
  or (_01374_, _01373_, _29617_);
  nor (_01375_, _01374_, _34815_);
  and (_01376_, _01375_, _35567_);
  and (_01377_, _01376_, _29157_);
  nor (_01378_, _01361_, _37727_);
  and (_01379_, _01378_, _01377_);
  and (_01380_, _01379_, _36306_);
  and (_01381_, _01380_, _29803_);
  and (_01382_, _01361_, _29518_);
  nor (_01383_, _01361_, _37585_);
  nor (_01384_, _01383_, _37728_);
  and (_01385_, _01384_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_01386_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_01387_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01388_, _01387_, _01386_);
  nor (_01389_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_01390_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01391_, _01390_, _01389_);
  and (_01392_, _01391_, _01388_);
  and (_01393_, _01392_, _37870_);
  or (_01394_, _01393_, _01385_);
  or (_01395_, _01394_, _01382_);
  nor (_01396_, _01395_, _01381_);
  not (_01397_, _00796_);
  nor (_01398_, _00995_, _37766_);
  and (_01399_, _01398_, _01397_);
  or (_01400_, _37783_, _37711_);
  or (_01401_, _01400_, _37775_);
  and (_01402_, _01401_, _37724_);
  nor (_01403_, _01402_, _00956_);
  and (_01404_, _01403_, _01399_);
  not (_01405_, _01404_);
  and (_01406_, _01405_, _01396_);
  and (_01407_, _37726_, _37505_);
  not (_01408_, _01407_);
  and (_01409_, _01408_, _37789_);
  nor (_01410_, _01409_, _01396_);
  nor (_01411_, _01410_, _01406_);
  and (_01412_, _01411_, _01372_);
  and (_01413_, _01412_, _37814_);
  nor (_01414_, _37835_, _37722_);
  nor (_01415_, _01414_, _01413_);
  nor (_01416_, _01415_, _01367_);
  and (_01417_, _38539_, _38659_);
  not (_01418_, _01417_);
  and (_01419_, _01418_, _37870_);
  nor (_01420_, _38365_, _38356_);
  and (_01421_, _01420_, _38448_);
  not (_01422_, _01421_);
  and (_01423_, _01422_, _01384_);
  nor (_01424_, _01423_, _01419_);
  not (_01425_, _01424_);
  nor (_01426_, _01425_, _01416_);
  not (_01427_, _01426_);
  nor (_01428_, _01427_, _01364_);
  and (_01429_, _01428_, _01360_);
  nor (_01430_, _37835_, rst);
  and (_38487_, _01430_, _01429_);
  and (_38488_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _42355_);
  and (_38489_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _42355_);
  nor (_01431_, _41842_, _37790_);
  and (_01432_, _37782_, _37724_);
  and (_01433_, _01432_, _36971_);
  nor (_01434_, _01433_, _01431_);
  and (_01435_, _01398_, _00954_);
  nor (_01436_, _01435_, _41842_);
  and (_01437_, _01365_, _36971_);
  nor (_01438_, _01437_, _37835_);
  not (_01439_, _01438_);
  nor (_01440_, _01439_, _01436_);
  and (_01441_, _01440_, _01434_);
  and (_01442_, _01441_, _01367_);
  and (_01443_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01444_, _01443_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01445_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01446_, _01445_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01447_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01448_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01449_, _01448_, _01447_);
  and (_01450_, _01449_, _01446_);
  and (_01451_, _01450_, _01444_);
  and (_01452_, _01451_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01453_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01454_, _01453_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_01455_, _01454_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_01456_, _01455_, _38050_);
  or (_01457_, _01455_, _38050_);
  and (_01458_, _01457_, _01456_);
  and (_01459_, _01458_, _01442_);
  and (_01460_, _37835_, _31235_);
  not (_01461_, _01434_);
  nor (_01462_, _00956_, _37726_);
  and (_01463_, _01462_, _01372_);
  nand (_01464_, _01463_, _01399_);
  and (_01465_, _01464_, _37722_);
  nor (_01466_, _01465_, _01461_);
  and (_01467_, _37712_, _37722_);
  nor (_01468_, _01467_, _01367_);
  and (_01469_, _01468_, _01441_);
  and (_01470_, _01469_, _01466_);
  and (_01471_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01472_, _01437_, _41768_);
  or (_01473_, _01472_, _01471_);
  not (_01474_, _38098_);
  and (_01475_, _01371_, _37722_);
  and (_01476_, _01475_, _01474_);
  or (_01477_, _01476_, _01473_);
  or (_01478_, _01477_, _01460_);
  or (_01479_, _01478_, _01459_);
  not (_01480_, _01429_);
  and (_01481_, _01441_, _41768_);
  nor (_01482_, _01441_, _01151_);
  nor (_01483_, _01482_, _01481_);
  not (_01484_, _01483_);
  not (_01485_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_01486_, _01483_, _01485_);
  and (_01487_, _01483_, _01485_);
  not (_01488_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01489_, _01441_, _42085_);
  nor (_01490_, _01441_, _01319_);
  nor (_01491_, _01490_, _01489_);
  nor (_01492_, _01491_, _01488_);
  and (_01493_, _01491_, _01488_);
  nor (_01494_, _01493_, _01492_);
  not (_01495_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01496_, _01441_, _42129_);
  nor (_01497_, _01441_, _01300_);
  nor (_01498_, _01497_, _01496_);
  nor (_01499_, _01498_, _01495_);
  and (_01500_, _01498_, _01495_);
  and (_01501_, _01441_, _41865_);
  nor (_01502_, _01441_, _01265_);
  nor (_01503_, _01502_, _01501_);
  not (_01504_, _01503_);
  nand (_01505_, _01504_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_01506_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01507_, _01441_, _41969_);
  nor (_01508_, _01441_, _01230_);
  nor (_01509_, _01508_, _01507_);
  nor (_01510_, _01509_, _01506_);
  and (_01511_, _01509_, _01506_);
  not (_01512_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01513_, _01441_, _42155_);
  nor (_01514_, _01441_, _01202_);
  nor (_01515_, _01514_, _01513_);
  nor (_01516_, _01515_, _01512_);
  not (_01517_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01518_, _01441_, _41934_);
  nor (_01519_, _01441_, _01185_);
  nor (_01520_, _01519_, _01518_);
  nor (_01521_, _01520_, _01517_);
  and (_01522_, _01441_, _42012_);
  nor (_01523_, _01441_, _01168_);
  nor (_01524_, _01523_, _01522_);
  not (_01525_, _01524_);
  and (_01526_, _01525_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_01527_, _01520_, _01517_);
  nor (_01528_, _01527_, _01521_);
  and (_01529_, _01528_, _01526_);
  nor (_01530_, _01529_, _01521_);
  not (_01531_, _01530_);
  and (_01532_, _01515_, _01512_);
  nor (_01533_, _01532_, _01516_);
  and (_01534_, _01533_, _01531_);
  nor (_01535_, _01534_, _01516_);
  nor (_01536_, _01535_, _01511_);
  or (_01537_, _01536_, _01510_);
  or (_01538_, _01504_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01539_, _01538_, _01505_);
  nand (_01540_, _01539_, _01537_);
  and (_01541_, _01540_, _01505_);
  nor (_01542_, _01541_, _01500_);
  or (_01543_, _01542_, _01499_);
  and (_01544_, _01543_, _01494_);
  nor (_01545_, _01544_, _01492_);
  nor (_01546_, _01545_, _01487_);
  or (_01547_, _01546_, _01486_);
  and (_01548_, _01444_, _01547_);
  and (_01549_, _01548_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01550_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01551_, _01550_, _01549_);
  nor (_01552_, _01551_, _01484_);
  nor (_01553_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01554_, _01553_, _38024_);
  and (_01555_, _01554_, _38029_);
  and (_01556_, _01555_, _38014_);
  and (_01557_, _01556_, _38035_);
  and (_01558_, _01557_, _38040_);
  nor (_01559_, _01558_, _01483_);
  nor (_01560_, _01559_, _01552_);
  or (_01561_, _01483_, _38045_);
  nand (_01562_, _01483_, _38045_);
  and (_01563_, _01562_, _01561_);
  and (_01564_, _01563_, _01560_);
  nand (_01565_, _01564_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_01566_, _01564_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_01567_, _01441_);
  or (_01568_, _01468_, _01567_);
  and (_01569_, _37724_, _36971_);
  and (_01570_, _01569_, _37782_);
  or (_01571_, _01570_, _01431_);
  or (_01572_, _01571_, _01465_);
  and (_01573_, _01572_, _01568_);
  and (_01574_, _01573_, _01566_);
  and (_01575_, _01574_, _01565_);
  or (_01576_, _01575_, _01480_);
  or (_01577_, _01576_, _01479_);
  and (_01578_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01579_, _37080_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01580_, _01579_, _41751_);
  nor (_01581_, _01580_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_01582_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_01583_, _01582_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_01584_, _01583_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_01585_, _01584_);
  nor (_01586_, _01585_, _01581_);
  and (_01587_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_01588_, _01587_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01589_, _01588_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01590_, _01589_, _01586_);
  and (_01591_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01592_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01593_, _01592_, _01578_);
  and (_01594_, _01593_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01595_, _01594_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_01596_, _01594_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_01597_, _01596_, _01595_);
  or (_01598_, _01597_, _01429_);
  and (_01599_, _01598_, _42355_);
  and (_38490_, _01599_, _01577_);
  and (_01600_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _42355_);
  and (_01601_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01602_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_01603_, _37025_, _01602_);
  not (_01604_, _01603_);
  not (_01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_01609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_01612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_01615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01616_, _01615_, _01614_);
  and (_01617_, _01616_, _01613_);
  and (_01618_, _01617_, _01612_);
  and (_01619_, _01618_, _01611_);
  and (_01620_, _01619_, _01610_);
  and (_01621_, _01620_, _01609_);
  and (_01622_, _01621_, _01608_);
  and (_01623_, _01622_, _01607_);
  and (_01624_, _01623_, _01606_);
  nor (_01625_, _01624_, _01605_);
  and (_01626_, _01624_, _01605_);
  nor (_01627_, _01626_, _01625_);
  nor (_01628_, _01623_, _01606_);
  nor (_01630_, _01628_, _01624_);
  and (_01631_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01634_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01636_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_01637_, _01636_, _01633_);
  and (_01639_, _01637_, _01634_);
  nor (_01640_, _01639_, _01633_);
  nor (_01642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_01643_, _01642_, _01631_);
  not (_01645_, _01643_);
  nor (_01646_, _01645_, _01640_);
  nor (_01648_, _01646_, _01631_);
  not (_01649_, _01648_);
  and (_01651_, _01649_, _01621_);
  and (_01652_, _01651_, _01608_);
  and (_01654_, _01652_, _01607_);
  not (_01655_, _01654_);
  nor (_01657_, _01655_, _01630_);
  and (_01658_, _01655_, _01630_);
  or (_01660_, _01658_, _01657_);
  not (_01661_, _01660_);
  and (_01662_, _01648_, _01623_);
  and (_01663_, _01648_, _01622_);
  nor (_01664_, _01663_, _01607_);
  nor (_01665_, _01664_, _01662_);
  not (_01666_, _01665_);
  and (_01667_, _01648_, _01621_);
  nor (_01668_, _01667_, _01608_);
  nor (_01669_, _01668_, _01663_);
  not (_01670_, _01669_);
  and (_01671_, _01648_, _01619_);
  and (_01672_, _01671_, _01610_);
  nor (_01673_, _01672_, _01609_);
  nor (_01674_, _01673_, _01667_);
  not (_01675_, _01674_);
  nor (_01676_, _01671_, _01610_);
  nor (_01677_, _01676_, _01672_);
  not (_01678_, _01677_);
  not (_01679_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_01680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01681_, _01648_, _01618_);
  and (_01682_, _01681_, _01680_);
  nor (_01683_, _01682_, _01679_);
  nor (_01684_, _01683_, _01671_);
  not (_01685_, _01684_);
  and (_01686_, _01648_, _01616_);
  and (_01687_, _01686_, _01613_);
  nor (_01688_, _01687_, _01612_);
  nor (_01689_, _01688_, _01681_);
  not (_01690_, _01689_);
  nor (_01691_, _01686_, _01613_);
  or (_01692_, _01691_, _01687_);
  and (_01693_, _01648_, _01615_);
  nor (_01694_, _01693_, _01614_);
  nor (_01695_, _01694_, _01686_);
  not (_01696_, _01695_);
  not (_01697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01698_, _01648_, _01697_);
  nor (_01699_, _01648_, _01697_);
  nor (_01700_, _01699_, _01698_);
  not (_01701_, _01700_);
  and (_01702_, _00635_, _00629_);
  not (_01703_, _01702_);
  nor (_01704_, _00665_, _00627_);
  nor (_01705_, _01704_, _01703_);
  not (_01706_, _00645_);
  and (_01707_, _00656_, _37579_);
  and (_01708_, _00667_, _00633_);
  nor (_01709_, _01708_, _01707_);
  nor (_01710_, _01709_, _01706_);
  nor (_01711_, _01710_, _01705_);
  nor (_01712_, _00704_, _01708_);
  nor (_01713_, _01712_, _37697_);
  not (_01714_, _00627_);
  and (_01715_, _00656_, _00651_);
  nor (_01716_, _01715_, _00668_);
  nor (_01717_, _01716_, _01714_);
  nor (_01718_, _01717_, _01713_);
  and (_01719_, _01718_, _01711_);
  and (_01720_, _00667_, _00627_);
  and (_01721_, _01720_, _00674_);
  not (_01722_, _00665_);
  and (_01723_, _00667_, _00629_);
  nor (_01724_, _01723_, _00636_);
  nor (_01725_, _01724_, _01722_);
  nor (_01726_, _01725_, _01721_);
  and (_01727_, _00628_, _00646_);
  and (_01728_, _00678_, _01727_);
  and (_01729_, _00667_, _00645_);
  and (_01730_, _01729_, _37429_);
  nor (_01731_, _01730_, _01728_);
  and (_01732_, _01731_, _01726_);
  and (_01733_, _01732_, _01719_);
  and (_01734_, _00677_, _00668_);
  not (_01735_, _01734_);
  nor (_01736_, _00689_, _00676_);
  and (_01737_, _01736_, _01735_);
  not (_01738_, _00688_);
  and (_01739_, _00656_, _00633_);
  nor (_01740_, _01739_, _00628_);
  nor (_01741_, _01740_, _01738_);
  not (_01742_, _01741_);
  or (_01743_, _00704_, _00706_);
  and (_01744_, _01743_, _00688_);
  not (_01745_, _00691_);
  and (_01746_, _00635_, _00646_);
  and (_01747_, _00658_, _01746_);
  and (_01748_, _00685_, _00667_);
  nor (_01749_, _01748_, _01747_);
  nor (_01750_, _01749_, _01745_);
  nor (_01751_, _01750_, _01744_);
  and (_01752_, _01751_, _01742_);
  and (_01753_, _01752_, _01737_);
  and (_01754_, _01753_, _01733_);
  and (_01755_, _00688_, _00668_);
  and (_01756_, _01702_, _00699_);
  or (_01757_, _01756_, _01755_);
  not (_01758_, _01757_);
  and (_01759_, _00677_, _00652_);
  nor (_01760_, _01759_, _00627_);
  not (_01761_, _00652_);
  nor (_01762_, _00704_, _00662_);
  and (_01763_, _01762_, _01761_);
  nor (_01764_, _01763_, _01760_);
  not (_01765_, _01764_);
  and (_01766_, _01765_, _00655_);
  and (_01767_, _01766_, _01758_);
  and (_01768_, _00680_, _37579_);
  not (_01769_, _01768_);
  nor (_01770_, _00707_, _00702_);
  and (_01771_, _01770_, _01769_);
  and (_01772_, _00706_, _00627_);
  and (_01773_, _00656_, _00647_);
  nor (_01774_, _01773_, _00652_);
  nor (_01775_, _01774_, _01738_);
  nor (_01776_, _01775_, _01772_);
  and (_01777_, _01776_, _01771_);
  and (_01778_, _00636_, _00626_);
  and (_01779_, _00704_, _00677_);
  nor (_01780_, _01779_, _01778_);
  and (_01781_, _00699_, _00652_);
  and (_01782_, _00706_, _00661_);
  nor (_01783_, _01782_, _01781_);
  and (_01784_, _01783_, _01780_);
  nor (_01785_, _00694_, _00663_);
  and (_01786_, _01715_, _00688_);
  and (_01787_, _00677_, _00648_);
  nor (_01788_, _01787_, _01786_);
  and (_01789_, _01788_, _01785_);
  and (_01790_, _01789_, _01784_);
  and (_01791_, _01790_, _01777_);
  and (_01792_, _01791_, _01767_);
  and (_01793_, _01792_, _01754_);
  nor (_01794_, _01637_, _01634_);
  nor (_01795_, _01794_, _01639_);
  not (_01796_, _01795_);
  nor (_01797_, _01796_, _01793_);
  not (_01798_, _01797_);
  nand (_01799_, _01758_, _01737_);
  or (_01800_, _00694_, _01768_);
  nor (_01801_, _01800_, _01744_);
  nand (_01802_, _01729_, _00629_);
  nand (_01803_, _00699_, _00636_);
  and (_01804_, _01803_, _01802_);
  nor (_01805_, _01781_, _00649_);
  and (_01806_, _01805_, _01804_);
  nand (_01807_, _01806_, _01801_);
  or (_01808_, _01807_, _01799_);
  nor (_01809_, _01808_, _01793_);
  not (_01810_, _01809_);
  nor (_01811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01812_, _01811_, _01634_);
  and (_01813_, _01812_, _01810_);
  and (_01814_, _01796_, _01793_);
  nor (_01815_, _01814_, _01797_);
  nand (_01816_, _01815_, _01813_);
  and (_01817_, _01816_, _01798_);
  not (_01818_, _01817_);
  and (_01819_, _01645_, _01640_);
  nor (_01820_, _01819_, _01646_);
  and (_01821_, _01820_, _01818_);
  and (_01822_, _01821_, _01701_);
  not (_01823_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_01824_, _01698_, _01823_);
  or (_01825_, _01824_, _01693_);
  and (_01826_, _01825_, _01822_);
  and (_01827_, _01826_, _01696_);
  and (_01828_, _01827_, _01692_);
  and (_01829_, _01828_, _01690_);
  nor (_01830_, _01681_, _01680_);
  or (_01831_, _01830_, _01682_);
  and (_01832_, _01831_, _01829_);
  and (_01833_, _01832_, _01685_);
  and (_01834_, _01833_, _01678_);
  and (_01835_, _01834_, _01675_);
  and (_01836_, _01835_, _01670_);
  and (_01837_, _01836_, _01666_);
  and (_01838_, _01837_, _01661_);
  nor (_01839_, _01838_, _01657_);
  not (_01840_, _01839_);
  nor (_01841_, _01840_, _01627_);
  and (_01842_, _01840_, _01627_);
  or (_01843_, _01842_, _01841_);
  or (_01844_, _01843_, _01604_);
  or (_01845_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_01846_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01847_, _01846_, _01845_);
  and (_01848_, _01847_, _01844_);
  or (_38492_, _01848_, _01601_);
  nor (_01849_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_38493_, _01849_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_38494_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _42355_);
  nor (_01850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_01851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01852_, _01851_, _01850_);
  nor (_01853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_01854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_01855_, _01854_, _01853_);
  and (_01856_, _01855_, _01852_);
  nor (_01857_, _01856_, rst);
  and (_01858_, \oc8051_top_1.oc8051_rom1.ea_int , _36993_);
  nand (_01859_, _01858_, _37025_);
  and (_01860_, _01859_, _38494_);
  or (_38495_, _01860_, _01857_);
  and (_01861_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_01862_, _01861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_38497_, _01862_, _42355_);
  nor (_01863_, _01581_, _41751_);
  or (_01864_, _01793_, _37232_);
  nor (_01865_, _01809_, _37167_);
  nand (_01866_, _01793_, _37232_);
  and (_01867_, _01866_, _01864_);
  nand (_01868_, _01867_, _01865_);
  and (_01869_, _01868_, _01864_);
  nor (_01870_, _01869_, _41751_);
  and (_01871_, _01870_, _37069_);
  nor (_01872_, _01870_, _37069_);
  nor (_01873_, _01872_, _01871_);
  nor (_01874_, _01873_, _01863_);
  and (_01875_, _37243_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_01876_, _01875_, _01863_);
  and (_01877_, _01876_, _01808_);
  or (_01878_, _01877_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01879_, _01878_, _01874_);
  and (_38498_, _01879_, _42355_);
  not (_01880_, _37646_);
  and (_01881_, _37551_, _01880_);
  not (_01882_, _37352_);
  and (_01883_, _37598_, _01882_);
  and (_01884_, _01883_, _01881_);
  and (_01885_, _37036_, _42355_);
  nand (_01886_, _01885_, _37670_);
  nor (_01887_, _01886_, _37693_);
  not (_01888_, _37575_);
  nor (_01889_, _01888_, _37624_);
  and (_01890_, _01889_, _01887_);
  and (_38501_, _01890_, _01884_);
  nor (_01891_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_01892_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_01893_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_38503_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _42355_);
  and (_01894_, _38503_, _01893_);
  or (_38502_, _01894_, _01892_);
  not (_01895_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01896_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01897_, _01896_, _01895_);
  and (_01898_, _01896_, _01895_);
  nor (_01899_, _01898_, _01897_);
  not (_01900_, _01899_);
  and (_01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01902_, _01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01903_, _01901_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01904_, _01903_, _01902_);
  or (_01905_, _01904_, _01896_);
  and (_01906_, _01905_, _01900_);
  nor (_01907_, _01897_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01908_, _01897_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01909_, _01908_, _01907_);
  or (_01910_, _01902_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_38505_, _01910_, _42355_);
  and (_01911_, _38505_, _01909_);
  and (_38504_, _01911_, _01906_);
  not (_01912_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_01913_, _01581_, _01912_);
  and (_01914_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_01915_, _01913_);
  and (_01916_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_01917_, _01916_, _01914_);
  and (_38506_, _01917_, _42355_);
  and (_01918_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_01919_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_01920_, _01919_, _01918_);
  and (_38507_, _01920_, _42355_);
  and (_01921_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_01922_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01923_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01922_);
  and (_01924_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01925_, _01924_, _01921_);
  and (_38508_, _01925_, _42355_);
  and (_01926_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01927_, _01926_, _01923_);
  and (_38509_, _01927_, _42355_);
  or (_01928_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_38511_, _01928_, _42355_);
  not (_01929_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_01930_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01931_, _01930_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_01932_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_01933_, _01932_, _42355_);
  and (_38512_, _01933_, _01931_);
  or (_01934_, _01922_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_38513_, _01934_, _42355_);
  nor (_01935_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_01936_, _01935_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_01937_, _01936_, _42355_);
  and (_01938_, _38503_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_38514_, _01938_, _01937_);
  and (_01939_, _01912_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_01940_, _01939_, _01936_);
  and (_38515_, _01940_, _42355_);
  nand (_01941_, _01936_, _38098_);
  or (_01942_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_01943_, _01942_, _42355_);
  and (_38516_, _01943_, _01941_);
  nand (_01944_, _37740_, _42355_);
  nor (_38517_, _01944_, _37874_);
  and (_01945_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_01946_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_01947_, _01946_, _01945_);
  and (_38555_, _01947_, _42355_);
  or (_01948_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_01949_, _01320_, _01517_);
  and (_01950_, _01949_, _42355_);
  and (_38556_, _01950_, _01948_);
  or (_01951_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_01952_, _01320_, _01512_);
  and (_01953_, _01952_, _42355_);
  and (_38557_, _01953_, _01951_);
  or (_01954_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_01955_, _01320_, _01506_);
  and (_01956_, _01955_, _42355_);
  and (_38558_, _01956_, _01954_);
  and (_01957_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01958_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_01959_, _01958_, _01957_);
  and (_38559_, _01959_, _42355_);
  or (_01960_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_01961_, _01320_, _01495_);
  and (_01962_, _01961_, _42355_);
  and (_38561_, _01962_, _01960_);
  or (_01963_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_01964_, _01320_, _01488_);
  and (_01965_, _01964_, _42355_);
  and (_38562_, _01965_, _01963_);
  or (_01966_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_01967_, _01320_, _01485_);
  and (_01968_, _01967_, _42355_);
  and (_38563_, _01968_, _01966_);
  or (_01969_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01970_, _01320_, _38018_);
  and (_01971_, _01970_, _42355_);
  and (_38564_, _01971_, _01969_);
  or (_01972_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01973_, _01320_, _38024_);
  and (_01974_, _01973_, _42355_);
  and (_38565_, _01974_, _01972_);
  or (_01975_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_01976_, _01320_, _38029_);
  and (_01977_, _01976_, _42355_);
  and (_38566_, _01977_, _01975_);
  or (_01978_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_01979_, _01320_, _38014_);
  and (_01980_, _01979_, _42355_);
  and (_38567_, _01980_, _01978_);
  or (_01981_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_01982_, _01320_, _38035_);
  and (_01983_, _01982_, _42355_);
  and (_38568_, _01983_, _01981_);
  or (_01984_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_01985_, _01320_, _38040_);
  and (_01986_, _01985_, _42355_);
  and (_38569_, _01986_, _01984_);
  or (_01987_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_01988_, _01320_, _38045_);
  and (_01989_, _01988_, _42355_);
  and (_38570_, _01989_, _01987_);
  and (_01990_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_01991_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_01992_, _01991_, _01990_);
  and (_38575_, _01992_, _42355_);
  and (_01993_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_01994_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_01995_, _01994_, _01993_);
  and (_38576_, _01995_, _42355_);
  and (_01996_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_01997_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_01998_, _01997_, _01996_);
  and (_38577_, _01998_, _42355_);
  and (_01999_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_02000_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_02001_, _02000_, _01999_);
  and (_38578_, _02001_, _42355_);
  and (_02002_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_02003_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_02004_, _02003_, _02002_);
  and (_38579_, _02004_, _42355_);
  and (_02005_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_02006_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or (_02007_, _02006_, _02005_);
  and (_38580_, _02007_, _42355_);
  and (_02008_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_02009_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or (_02010_, _02009_, _02008_);
  and (_38581_, _02010_, _42355_);
  and (_02011_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_02012_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or (_02013_, _02012_, _02011_);
  and (_38582_, _02013_, _42355_);
  and (_02014_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_02015_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or (_02016_, _02015_, _02014_);
  and (_38583_, _02016_, _42355_);
  and (_02017_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02018_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02019_, _02018_, _02017_);
  and (_38584_, _02019_, _42355_);
  and (_02020_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_02021_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02022_, _02021_, _02020_);
  and (_38586_, _02022_, _42355_);
  and (_02023_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_02024_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or (_02025_, _02024_, _02023_);
  and (_38587_, _02025_, _42355_);
  and (_02026_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_02027_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or (_02028_, _02027_, _02026_);
  and (_38588_, _02028_, _42355_);
  and (_02029_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_02030_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or (_02031_, _02030_, _02029_);
  and (_38589_, _02031_, _42355_);
  and (_02032_, _01320_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_02033_, _01324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_02034_, _02033_, _02032_);
  and (_38590_, _02034_, _42355_);
  and (_38766_, _37633_, _42355_);
  and (_38767_, _37657_, _42355_);
  and (_38768_, _37679_, _42355_);
  nor (_38769_, _41774_, rst);
  and (_02035_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02036_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_02037_, _02036_, _02035_);
  and (_38770_, _02037_, _42355_);
  and (_02038_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02039_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_02040_, _02039_, _02038_);
  and (_38771_, _02040_, _42355_);
  and (_02041_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02042_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_02043_, _02042_, _02041_);
  and (_38772_, _02043_, _42355_);
  and (_02044_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02045_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_02046_, _02045_, _01913_);
  or (_02047_, _02046_, _02044_);
  and (_38773_, _02047_, _42355_);
  and (_02048_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02049_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_02050_, _02049_, _02048_);
  and (_38775_, _02050_, _42355_);
  and (_02051_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02052_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_02053_, _02052_, _02051_);
  and (_38776_, _02053_, _42355_);
  and (_02054_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02055_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_02056_, _02055_, _02054_);
  and (_38777_, _02056_, _42355_);
  and (_02057_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02058_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_02059_, _02058_, _02057_);
  and (_38778_, _02059_, _42355_);
  and (_02060_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_02061_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_02062_, _02061_, _02060_);
  and (_38779_, _02062_, _42355_);
  and (_02063_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_02064_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_02065_, _02064_, _02063_);
  and (_38780_, _02065_, _42355_);
  and (_02066_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_02067_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_02068_, _02067_, _02066_);
  and (_38781_, _02068_, _42355_);
  and (_02069_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_02070_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_02071_, _02070_, _02069_);
  and (_38782_, _02071_, _42355_);
  and (_02072_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_02073_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_02074_, _02073_, _02072_);
  and (_38783_, _02074_, _42355_);
  and (_02075_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_02076_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_02077_, _02076_, _02075_);
  and (_38784_, _02077_, _42355_);
  and (_02078_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_02079_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_02080_, _02079_, _02078_);
  and (_38786_, _02080_, _42355_);
  and (_02081_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_02082_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_02083_, _02082_, _02081_);
  and (_38787_, _02083_, _42355_);
  and (_02084_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_02085_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_02086_, _02085_, _02084_);
  and (_38788_, _02086_, _42355_);
  and (_02087_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_02088_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_02089_, _02088_, _02087_);
  and (_38789_, _02089_, _42355_);
  and (_02090_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_02091_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_02092_, _02091_, _02090_);
  and (_38790_, _02092_, _42355_);
  and (_02093_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_02094_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_02095_, _02094_, _02093_);
  and (_38791_, _02095_, _42355_);
  and (_02096_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_02097_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_02098_, _02097_, _02096_);
  and (_38792_, _02098_, _42355_);
  and (_02099_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_02100_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_02101_, _02100_, _02099_);
  and (_38793_, _02101_, _42355_);
  and (_02102_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_02103_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_02104_, _02103_, _02102_);
  and (_38794_, _02104_, _42355_);
  and (_02105_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_02106_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_02107_, _02106_, _02105_);
  and (_38795_, _02107_, _42355_);
  and (_02108_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_02109_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_02111_, _02109_, _02108_);
  and (_38797_, _02111_, _42355_);
  and (_02114_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_02116_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_02118_, _02116_, _02114_);
  and (_38798_, _02118_, _42355_);
  and (_02121_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_02123_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_02125_, _02123_, _02121_);
  and (_38799_, _02125_, _42355_);
  and (_02128_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_02130_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_02132_, _02130_, _02128_);
  and (_38800_, _02132_, _42355_);
  and (_02135_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_02137_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_02139_, _02137_, _02135_);
  and (_38801_, _02139_, _42355_);
  and (_02142_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_02144_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_02146_, _02144_, _02142_);
  and (_38802_, _02146_, _42355_);
  and (_02149_, _01913_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_02151_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_02153_, _02151_, _02149_);
  and (_38803_, _02153_, _42355_);
  and (_38804_, _42034_, _42355_);
  and (_38806_, _41914_, _42355_);
  and (_38807_, _42177_, _42355_);
  and (_38808_, _41991_, _42355_);
  and (_38809_, _41886_, _42355_);
  and (_38810_, _42113_, _42355_);
  and (_38812_, _42066_, _42355_);
  and (_38828_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _42355_);
  and (_38829_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _42355_);
  and (_38830_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _42355_);
  and (_38831_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _42355_);
  and (_38832_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _42355_);
  and (_38834_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _42355_);
  and (_38835_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _42355_);
  or (_02164_, _01470_, _01467_);
  and (_02165_, _02164_, _32455_);
  and (_02166_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not (_02167_, _01168_);
  and (_02168_, _01437_, _02167_);
  and (_02169_, _01522_, _01367_);
  or (_02170_, _02169_, _02168_);
  or (_02171_, _01525_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02172_, _01526_);
  and (_02173_, _01573_, _02172_);
  and (_02174_, _02173_, _02171_);
  or (_02175_, _02174_, _02170_);
  nor (_02176_, _02175_, _02166_);
  nand (_02177_, _02176_, _01429_);
  or (_02178_, _02177_, _02165_);
  or (_02179_, _01429_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_02180_, _02179_, _42355_);
  and (_38836_, _02180_, _02178_);
  and (_02181_, _02164_, _33130_);
  and (_02182_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  not (_02183_, _01185_);
  and (_02184_, _01437_, _02183_);
  and (_02185_, _01518_, _01367_);
  or (_02186_, _02185_, _02184_);
  or (_02187_, _02186_, _02182_);
  or (_02188_, _01528_, _01526_);
  not (_02189_, _01529_);
  and (_02190_, _01573_, _02189_);
  and (_02191_, _02190_, _02188_);
  nor (_02192_, _02191_, _02187_);
  nand (_02193_, _02192_, _01429_);
  or (_02194_, _02193_, _02181_);
  or (_02195_, _01429_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_02196_, _02195_, _42355_);
  and (_38837_, _02196_, _02194_);
  and (_02197_, _02164_, _33848_);
  and (_02198_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not (_02199_, _01202_);
  and (_02200_, _01437_, _02199_);
  and (_02201_, _01513_, _01367_);
  or (_02202_, _02201_, _02200_);
  or (_02203_, _01533_, _01531_);
  not (_02204_, _01534_);
  and (_02205_, _01573_, _02204_);
  and (_02206_, _02205_, _02203_);
  or (_02207_, _02206_, _02202_);
  nor (_02208_, _02207_, _02198_);
  nand (_02209_, _02208_, _01429_);
  or (_02210_, _02209_, _02197_);
  not (_02211_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02212_, _01581_, _02211_);
  and (_02213_, _01581_, _02211_);
  nor (_02214_, _02213_, _02212_);
  or (_02215_, _02214_, _01429_);
  and (_02216_, _02215_, _42355_);
  and (_38838_, _02216_, _02210_);
  and (_02217_, _02164_, _34566_);
  and (_02218_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not (_02219_, _01230_);
  and (_02220_, _01437_, _02219_);
  and (_02221_, _01507_, _01367_);
  or (_02222_, _02221_, _02220_);
  or (_02223_, _02222_, _02218_);
  or (_02224_, _02223_, _02217_);
  or (_02225_, _01511_, _01510_);
  or (_02226_, _02225_, _01535_);
  nand (_02227_, _02225_, _01535_);
  and (_02228_, _02227_, _02226_);
  nand (_02229_, _02228_, _01573_);
  nand (_02230_, _02229_, _01429_);
  or (_02231_, _02230_, _02224_);
  and (_02232_, _02212_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02233_, _02212_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02234_, _02233_, _02232_);
  or (_02235_, _02234_, _01429_);
  and (_02236_, _02235_, _42355_);
  and (_38839_, _02236_, _02231_);
  and (_02237_, _02164_, _35229_);
  and (_02238_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  not (_02239_, _01265_);
  and (_02240_, _01437_, _02239_);
  and (_02241_, _01442_, _41865_);
  or (_02242_, _02241_, _02240_);
  or (_02243_, _01539_, _01537_);
  and (_02244_, _01573_, _01540_);
  and (_02245_, _02244_, _02243_);
  or (_02246_, _02245_, _02242_);
  nor (_02247_, _02246_, _02238_);
  nand (_02248_, _02247_, _01429_);
  or (_02249_, _02248_, _02237_);
  not (_02250_, _01581_);
  and (_02251_, _01583_, _02250_);
  nor (_02252_, _02232_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02253_, _02252_, _02251_);
  or (_02254_, _02253_, _01429_);
  and (_02255_, _02254_, _42355_);
  and (_38840_, _02255_, _02249_);
  and (_02256_, _02164_, _36035_);
  and (_02257_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_02258_, _01300_);
  and (_02259_, _01437_, _02258_);
  and (_02260_, _01496_, _01367_);
  or (_02261_, _02260_, _02259_);
  or (_02262_, _01500_, _01499_);
  or (_02263_, _02262_, _01541_);
  nand (_02264_, _02262_, _01541_);
  and (_02265_, _02264_, _01573_);
  and (_02266_, _02265_, _02263_);
  or (_02267_, _02266_, _02261_);
  nor (_02268_, _02267_, _02257_);
  nand (_02269_, _02268_, _01429_);
  or (_02270_, _02269_, _02256_);
  nor (_02271_, _02251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_02272_, _02271_, _01586_);
  or (_02273_, _02272_, _01429_);
  and (_02274_, _02273_, _42355_);
  and (_38841_, _02274_, _02270_);
  nor (_02275_, _01586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02276_, _01586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02277_, _02276_, _02275_);
  or (_02278_, _02277_, _01429_);
  and (_02279_, _02278_, _42355_);
  and (_02280_, _02164_, _36763_);
  and (_02281_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_02282_, _01319_);
  and (_02283_, _01437_, _02282_);
  and (_02284_, _01489_, _01367_);
  or (_02285_, _02284_, _02283_);
  or (_02286_, _02285_, _02281_);
  or (_02287_, _01543_, _01494_);
  not (_02288_, _01544_);
  and (_02289_, _01573_, _02288_);
  and (_02290_, _02289_, _02287_);
  nor (_02291_, _02290_, _02286_);
  nand (_02292_, _02291_, _01429_);
  or (_02293_, _02292_, _02280_);
  and (_38842_, _02293_, _02279_);
  or (_02294_, _01486_, _01487_);
  or (_02295_, _02294_, _01545_);
  nand (_02296_, _02294_, _01545_);
  and (_02297_, _02296_, _02295_);
  and (_02298_, _02297_, _01573_);
  and (_02299_, _02164_, _31235_);
  and (_02300_, _37835_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_02301_, _01151_);
  and (_02302_, _01437_, _02301_);
  and (_02303_, _01442_, _41768_);
  or (_02304_, _02303_, _02302_);
  or (_02305_, _02304_, _02300_);
  or (_02306_, _02305_, _02299_);
  or (_02307_, _02306_, _02298_);
  or (_02308_, _02307_, _01480_);
  nor (_02309_, _02276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02310_, _02276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_02311_, _02310_, _02309_);
  or (_02312_, _02311_, _01429_);
  and (_02313_, _02312_, _42355_);
  and (_38843_, _02313_, _02308_);
  and (_02314_, _37835_, _32455_);
  and (_02315_, _01547_, _38018_);
  nor (_02316_, _01547_, _38018_);
  nor (_02317_, _02316_, _02315_);
  nor (_02318_, _02317_, _01484_);
  and (_02319_, _02317_, _01484_);
  or (_02320_, _02319_, _02318_);
  and (_02321_, _02320_, _01573_);
  and (_02322_, _01442_, _00646_);
  and (_02323_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_02324_, _01437_, _42012_);
  or (_02325_, _02324_, _02323_);
  or (_02326_, _02325_, _02322_);
  not (_02327_, _38137_);
  and (_02328_, _01475_, _02327_);
  or (_02329_, _02328_, _02326_);
  or (_02330_, _02329_, _02321_);
  or (_02331_, _02330_, _02314_);
  or (_02332_, _02331_, _01480_);
  or (_02333_, _02310_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_02334_, _01588_, _01586_);
  and (_02335_, _02334_, _02333_);
  or (_02336_, _02335_, _01429_);
  and (_02337_, _02336_, _42355_);
  and (_38845_, _02337_, _02332_);
  and (_02338_, _37835_, _33130_);
  not (_02339_, _38168_);
  and (_02340_, _01467_, _02339_);
  and (_02341_, _01442_, _00634_);
  and (_02342_, _01437_, _41934_);
  or (_02343_, _02342_, _02341_);
  and (_02344_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_02345_, _02344_, _02343_);
  or (_02346_, _02345_, _02340_);
  or (_02347_, _02346_, _02338_);
  and (_02348_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02349_, _02348_, _01483_);
  and (_02350_, _01553_, _01484_);
  nor (_02351_, _02350_, _02349_);
  nand (_02352_, _02351_, _38024_);
  or (_02353_, _02351_, _38024_);
  and (_02354_, _02353_, _02352_);
  and (_02355_, _02354_, _01573_);
  or (_02356_, _02355_, _01480_);
  or (_02357_, _02356_, _02347_);
  nand (_02359_, _02334_, _01679_);
  or (_02360_, _02334_, _01679_);
  and (_02361_, _02360_, _02359_);
  or (_02362_, _02361_, _01429_);
  and (_02363_, _02362_, _42355_);
  and (_38846_, _02363_, _02357_);
  and (_02364_, _01554_, _01484_);
  and (_02365_, _02349_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02366_, _02365_, _02364_);
  nor (_02367_, _02366_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_02368_, _02366_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_02369_, _02368_, _02367_);
  and (_02370_, _02369_, _01573_);
  and (_02371_, _37835_, _33848_);
  not (_02372_, _38198_);
  and (_02373_, _01467_, _02372_);
  and (_02374_, _01437_, _42155_);
  and (_02375_, _01442_, _00666_);
  and (_02376_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_02377_, _02376_, _02375_);
  or (_02378_, _02377_, _02374_);
  or (_02379_, _02378_, _02373_);
  or (_02380_, _02379_, _02371_);
  or (_02381_, _02380_, _02370_);
  or (_02382_, _02381_, _01480_);
  nor (_02383_, _01590_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_02384_, _02383_, _01591_);
  or (_02385_, _02384_, _01429_);
  and (_02386_, _02385_, _42355_);
  and (_38847_, _02386_, _02382_);
  and (_02387_, _01548_, _01483_);
  and (_02388_, _01555_, _01484_);
  nor (_02389_, _02388_, _02387_);
  nor (_02390_, _02389_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02391_, _02389_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_02392_, _02391_, _02390_);
  and (_02393_, _02392_, _01573_);
  and (_02394_, _37835_, _34566_);
  and (_02395_, _01467_, _38226_);
  and (_02396_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02397_, _01451_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02398_, _02397_, _01452_);
  and (_02399_, _02398_, _01442_);
  and (_02400_, _01437_, _41969_);
  or (_02401_, _02400_, _02399_);
  or (_02402_, _02401_, _02396_);
  or (_02403_, _02402_, _02395_);
  or (_02404_, _02403_, _02394_);
  or (_02405_, _02404_, _02393_);
  or (_02406_, _02405_, _01480_);
  nor (_02407_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02408_, _02407_, _01592_);
  or (_02409_, _02408_, _01429_);
  and (_02410_, _02409_, _42355_);
  and (_38848_, _02410_, _02406_);
  and (_02411_, _37835_, _35229_);
  and (_02412_, _01467_, _38256_);
  and (_02413_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02414_, _01452_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02415_, _02414_, _01453_);
  and (_02416_, _02415_, _01442_);
  and (_02417_, _01437_, _41865_);
  or (_02418_, _02417_, _02416_);
  or (_02419_, _02418_, _02413_);
  or (_02420_, _02419_, _02412_);
  and (_02421_, _01549_, _01483_);
  and (_02422_, _01556_, _01484_);
  nor (_02423_, _02422_, _02421_);
  nand (_02424_, _02423_, _38035_);
  or (_02425_, _02423_, _38035_);
  and (_02426_, _02425_, _02424_);
  and (_02427_, _02426_, _01573_);
  or (_02428_, _02427_, _02420_);
  or (_02429_, _02428_, _02411_);
  or (_02430_, _02429_, _01480_);
  nor (_02431_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02432_, _01584_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02433_, _02432_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02434_, _02433_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_02435_, _02434_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_02436_, _02435_, _02250_);
  and (_02437_, _02436_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_02438_, _02437_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_02439_, _02438_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_02440_, _02439_, _02431_);
  or (_02441_, _02440_, _01429_);
  and (_02442_, _02441_, _42355_);
  and (_38849_, _02442_, _02430_);
  and (_02443_, _37835_, _36035_);
  and (_02444_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02445_, _01437_, _42129_);
  or (_02446_, _02445_, _02444_);
  not (_02447_, _38291_);
  and (_02448_, _01475_, _02447_);
  or (_02449_, _02448_, _02446_);
  nor (_02450_, _01453_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_02451_, _02450_, _01454_);
  and (_02452_, _02451_, _01442_);
  and (_02453_, _01483_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02454_, _02453_, _01549_);
  and (_02455_, _01557_, _01484_);
  nor (_02456_, _02455_, _02454_);
  or (_02457_, _02456_, _38040_);
  nand (_02458_, _02456_, _38040_);
  and (_02459_, _02458_, _01573_);
  and (_02460_, _02459_, _02457_);
  or (_02461_, _02460_, _02452_);
  or (_02462_, _02461_, _02449_);
  or (_02463_, _02462_, _02443_);
  and (_02464_, _02463_, _01429_);
  nor (_02465_, _02439_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_02466_, _02465_, _01593_);
  nor (_02467_, _02466_, _01429_);
  or (_02468_, _02467_, _02464_);
  and (_38850_, _02468_, _42355_);
  and (_02469_, _37835_, _36763_);
  and (_02470_, _01470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_02471_, _01437_, _42085_);
  or (_02472_, _02471_, _02470_);
  and (_02473_, _01475_, _38317_);
  or (_02474_, _02473_, _02472_);
  or (_02475_, _01454_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02476_, _02475_, _01455_);
  and (_02477_, _02476_, _01442_);
  nand (_02478_, _01560_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_02479_, _01560_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02480_, _02479_, _01573_);
  and (_02481_, _02480_, _02478_);
  or (_02482_, _02481_, _02477_);
  or (_02483_, _02482_, _02474_);
  or (_02484_, _02483_, _02469_);
  or (_02485_, _02484_, _01480_);
  nor (_02486_, _01593_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02487_, _02486_, _01594_);
  or (_02488_, _02487_, _01429_);
  and (_02489_, _02488_, _42355_);
  and (_38851_, _02489_, _02485_);
  and (_02490_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_02491_, _01812_, _01810_);
  nor (_02492_, _02491_, _01813_);
  or (_02493_, _02492_, _01604_);
  or (_02494_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02495_, _02494_, _01846_);
  and (_02496_, _02495_, _02493_);
  or (_38852_, _02496_, _02490_);
  or (_02497_, _01815_, _01813_);
  and (_02498_, _02497_, _01816_);
  or (_02499_, _02498_, _01604_);
  or (_02500_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02501_, _02500_, _01846_);
  and (_02502_, _02501_, _02499_);
  and (_02503_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_38853_, _02503_, _02502_);
  and (_02504_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_02505_, _01820_, _01818_);
  nor (_02506_, _02505_, _01821_);
  or (_02507_, _02506_, _01604_);
  or (_02508_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_02509_, _02508_, _01846_);
  and (_02510_, _02509_, _02507_);
  or (_38854_, _02510_, _02504_);
  and (_02511_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_02512_, _01821_, _01701_);
  nor (_02513_, _02512_, _01822_);
  or (_02514_, _02513_, _01604_);
  or (_02515_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_02516_, _02515_, _01846_);
  and (_02517_, _02516_, _02514_);
  or (_38855_, _02517_, _02511_);
  and (_02518_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_02519_, _01825_, _01822_);
  nor (_02520_, _02519_, _01826_);
  or (_02521_, _02520_, _01604_);
  or (_02522_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_02523_, _02522_, _01846_);
  and (_02524_, _02523_, _02521_);
  or (_38856_, _02524_, _02518_);
  nor (_02525_, _01826_, _01696_);
  nor (_02526_, _02525_, _01827_);
  or (_02527_, _02526_, _01604_);
  or (_02528_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_02529_, _02528_, _01846_);
  and (_02530_, _02529_, _02527_);
  and (_02531_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_38857_, _02531_, _02530_);
  nor (_02532_, _01827_, _01692_);
  nor (_02533_, _02532_, _01828_);
  or (_02534_, _02533_, _01604_);
  or (_02535_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02536_, _02535_, _01846_);
  and (_02537_, _02536_, _02534_);
  and (_02538_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_38858_, _02538_, _02537_);
  nor (_02539_, _01828_, _01690_);
  nor (_02540_, _02539_, _01829_);
  or (_02541_, _02540_, _01604_);
  or (_02542_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_02543_, _02542_, _01846_);
  and (_02544_, _02543_, _02541_);
  and (_02545_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_38859_, _02545_, _02544_);
  nor (_02547_, _01831_, _01829_);
  nor (_02548_, _02547_, _01832_);
  or (_02549_, _02548_, _01604_);
  or (_02550_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_02551_, _02550_, _01846_);
  and (_02552_, _02551_, _02549_);
  and (_02553_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_38860_, _02553_, _02552_);
  nor (_02554_, _01832_, _01685_);
  nor (_02555_, _02554_, _01833_);
  or (_02556_, _02555_, _01604_);
  or (_02557_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_02558_, _02557_, _01846_);
  and (_02559_, _02558_, _02556_);
  and (_02560_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_38861_, _02560_, _02559_);
  or (_02561_, _01833_, _01678_);
  nor (_02562_, _01604_, _01834_);
  and (_02563_, _02562_, _02561_);
  nor (_02564_, _01603_, _38029_);
  or (_02565_, _02564_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02566_, _02565_, _02563_);
  or (_02568_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _36993_);
  and (_02569_, _02568_, _42355_);
  and (_38862_, _02569_, _02566_);
  and (_02570_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_02571_, _01834_, _01675_);
  nor (_02572_, _02571_, _01835_);
  or (_02573_, _02572_, _01604_);
  or (_02574_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_02575_, _02574_, _01846_);
  and (_02576_, _02575_, _02573_);
  or (_38863_, _02576_, _02570_);
  nor (_02578_, _01835_, _01670_);
  nor (_02579_, _02578_, _01836_);
  or (_02580_, _02579_, _01604_);
  or (_02581_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_02582_, _02581_, _01846_);
  and (_02583_, _02582_, _02580_);
  and (_02584_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_38864_, _02584_, _02583_);
  nor (_02585_, _01836_, _01666_);
  nor (_02586_, _02585_, _01837_);
  or (_02587_, _02586_, _01604_);
  or (_02588_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_02589_, _02588_, _01846_);
  and (_02590_, _02589_, _02587_);
  and (_02591_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_38866_, _02591_, _02590_);
  and (_02592_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_02593_, _01837_, _01661_);
  nor (_02594_, _02593_, _01838_);
  or (_02595_, _02594_, _01604_);
  or (_02596_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02597_, _02596_, _01846_);
  and (_02598_, _02597_, _02595_);
  or (_38867_, _02598_, _02592_);
  and (_02599_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_02600_, _02599_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_38868_, _02600_, _42355_);
  and (_02601_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_02602_, _02601_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_38869_, _02602_, _42355_);
  and (_02603_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_02604_, _02603_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_38870_, _02604_, _42355_);
  and (_02605_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_02606_, _02605_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_38871_, _02606_, _42355_);
  and (_02607_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_02608_, _02607_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_38872_, _02608_, _42355_);
  and (_02609_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_02610_, _02609_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_38873_, _02610_, _42355_);
  and (_02611_, _01856_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_02612_, _02611_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_38874_, _02612_, _42355_);
  nor (_02613_, _01809_, _41751_);
  nand (_02614_, _02613_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_02615_, _02613_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_02616_, _02615_, _01846_);
  and (_38875_, _02616_, _02614_);
  or (_02617_, _01867_, _01865_);
  and (_02618_, _02617_, _01868_);
  or (_02619_, _02618_, _41751_);
  or (_02620_, _37025_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_02621_, _02620_, _01846_);
  and (_38877_, _02621_, _02619_);
  and (_02622_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_02623_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_02624_, _02623_, _38503_);
  or (_38893_, _02624_, _02622_);
  and (_02625_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_02626_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_02627_, _02626_, _38503_);
  or (_38894_, _02627_, _02625_);
  and (_02628_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_02629_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_02630_, _02629_, _38503_);
  or (_38895_, _02630_, _02628_);
  and (_02631_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_02632_, _02045_, _38503_);
  or (_38896_, _02632_, _02631_);
  and (_02633_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_02634_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_02635_, _02634_, _38503_);
  or (_38897_, _02635_, _02633_);
  and (_02636_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_02637_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_02638_, _02637_, _38503_);
  or (_38899_, _02638_, _02636_);
  and (_02639_, _01891_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_02640_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_02641_, _02640_, _38503_);
  or (_38900_, _02641_, _02639_);
  and (_38901_, _01899_, _42355_);
  nor (_38902_, _01909_, rst);
  and (_38903_, _01905_, _42355_);
  and (_02642_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_02643_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_02644_, _02643_, _02642_);
  and (_38904_, _02644_, _42355_);
  and (_02645_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_02646_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_02647_, _02646_, _02645_);
  and (_38905_, _02647_, _42355_);
  and (_02648_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_02649_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_02650_, _02649_, _02648_);
  and (_38906_, _02650_, _42355_);
  and (_02651_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_02652_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_02653_, _02652_, _02651_);
  and (_38907_, _02653_, _42355_);
  and (_02654_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_02655_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_02656_, _02655_, _02654_);
  and (_38908_, _02656_, _42355_);
  and (_02657_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_02658_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_02659_, _02658_, _02657_);
  and (_38910_, _02659_, _42355_);
  and (_02660_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_02661_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_02662_, _02661_, _02660_);
  and (_38911_, _02662_, _42355_);
  and (_02663_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_02664_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_02665_, _02664_, _02663_);
  and (_38912_, _02665_, _42355_);
  and (_02666_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_02667_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_02668_, _02667_, _02666_);
  and (_38913_, _02668_, _42355_);
  and (_02669_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_02670_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_02671_, _02670_, _02669_);
  and (_38914_, _02671_, _42355_);
  and (_02672_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_02673_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_02674_, _02673_, _02672_);
  and (_38915_, _02674_, _42355_);
  and (_02675_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_02676_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_02677_, _02676_, _02675_);
  and (_38916_, _02677_, _42355_);
  and (_02678_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_02679_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_02680_, _02679_, _02678_);
  and (_38917_, _02680_, _42355_);
  and (_02681_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_02682_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_02683_, _02682_, _02681_);
  and (_38918_, _02683_, _42355_);
  and (_02684_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_02685_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_02686_, _02685_, _02684_);
  and (_38919_, _02686_, _42355_);
  and (_02687_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_02688_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_02689_, _02688_, _02687_);
  and (_38921_, _02689_, _42355_);
  and (_02690_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_02691_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_02692_, _02691_, _02690_);
  and (_38922_, _02692_, _42355_);
  and (_02693_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_02694_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_02695_, _02694_, _02693_);
  and (_38923_, _02695_, _42355_);
  and (_02696_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_02697_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_02698_, _02697_, _02696_);
  and (_38924_, _02698_, _42355_);
  and (_02699_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_02700_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_02701_, _02700_, _02699_);
  and (_38925_, _02701_, _42355_);
  and (_02703_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02704_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_02705_, _02704_, _02703_);
  and (_38926_, _02705_, _42355_);
  and (_02706_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02707_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_02708_, _02707_, _02706_);
  and (_38927_, _02708_, _42355_);
  and (_02709_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_02710_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_02711_, _02710_, _02709_);
  and (_38928_, _02711_, _42355_);
  and (_02712_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_02713_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_02714_, _02713_, _02712_);
  and (_38929_, _02714_, _42355_);
  and (_02715_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_02716_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_02717_, _02716_, _02715_);
  and (_38930_, _02717_, _42355_);
  and (_02718_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_02719_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_02720_, _02719_, _02718_);
  and (_38932_, _02720_, _42355_);
  and (_02721_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_02722_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_02723_, _02722_, _02721_);
  and (_38933_, _02723_, _42355_);
  and (_02724_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_02725_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_02726_, _02725_, _02724_);
  and (_38934_, _02726_, _42355_);
  and (_02727_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_02728_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_02729_, _02728_, _02727_);
  and (_38935_, _02729_, _42355_);
  and (_02730_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_02731_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_02732_, _02731_, _02730_);
  and (_38936_, _02732_, _42355_);
  and (_02733_, _01913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_02734_, _01915_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_02735_, _02734_, _02733_);
  and (_38937_, _02735_, _42355_);
  and (_02736_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02737_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_02738_, _02737_, _02736_);
  and (_38938_, _02738_, _42355_);
  and (_02739_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02740_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_02741_, _02740_, _02739_);
  and (_38939_, _02741_, _42355_);
  and (_02742_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02743_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_02744_, _02743_, _02742_);
  and (_38940_, _02744_, _42355_);
  and (_02745_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02746_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_02747_, _02746_, _02745_);
  and (_38941_, _02747_, _42355_);
  and (_02748_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02749_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_02750_, _02749_, _02748_);
  and (_38943_, _02750_, _42355_);
  and (_02751_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02752_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_02753_, _02752_, _02751_);
  and (_38944_, _02753_, _42355_);
  and (_02754_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_02755_, _01923_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_02756_, _02755_, _02754_);
  and (_38945_, _02756_, _42355_);
  and (_02757_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02758_, _42034_, _01929_);
  or (_02759_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_02760_, _02759_, _01922_);
  and (_02761_, _02760_, _02758_);
  or (_02762_, _02761_, _02757_);
  and (_38946_, _02762_, _42355_);
  and (_02763_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02764_, _41914_, _01929_);
  or (_02765_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_02766_, _02765_, _01922_);
  and (_02767_, _02766_, _02764_);
  or (_02768_, _02767_, _02763_);
  and (_38947_, _02768_, _42355_);
  and (_02769_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02770_, _42177_, _01929_);
  or (_02771_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_02772_, _02771_, _01922_);
  and (_02773_, _02772_, _02770_);
  or (_02774_, _02773_, _02769_);
  and (_38948_, _02774_, _42355_);
  and (_02775_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02776_, _41991_, _01929_);
  or (_02777_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_02778_, _02777_, _01922_);
  and (_02779_, _02778_, _02776_);
  or (_02780_, _02779_, _02775_);
  and (_38949_, _02780_, _42355_);
  and (_02781_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02782_, _41886_, _01929_);
  or (_02783_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_02784_, _02783_, _01922_);
  and (_02785_, _02784_, _02782_);
  or (_02786_, _02785_, _02781_);
  and (_38950_, _02786_, _42355_);
  and (_02787_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02788_, _42113_, _01929_);
  or (_02789_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_02790_, _02789_, _01922_);
  and (_02791_, _02790_, _02788_);
  or (_02792_, _02791_, _02787_);
  and (_38951_, _02792_, _42355_);
  and (_02793_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02794_, _42066_, _01929_);
  or (_02795_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02796_, _02795_, _01922_);
  and (_02797_, _02796_, _02794_);
  or (_02798_, _02797_, _02793_);
  and (_38952_, _02798_, _42355_);
  and (_02799_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02800_, _41825_, _01929_);
  or (_02802_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_02803_, _02802_, _01922_);
  and (_02804_, _02803_, _02800_);
  or (_02805_, _02804_, _02799_);
  and (_38954_, _02805_, _42355_);
  and (_02807_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_02808_, _02807_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02809_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01922_);
  and (_02810_, _02809_, _42355_);
  and (_38955_, _02810_, _02808_);
  and (_02812_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_02813_, _02812_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02814_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01922_);
  and (_02815_, _02814_, _42355_);
  and (_38956_, _02815_, _02813_);
  and (_02817_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_02818_, _02817_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02819_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01922_);
  and (_02820_, _02819_, _42355_);
  and (_38957_, _02820_, _02818_);
  and (_02822_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_02823_, _02822_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02824_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01922_);
  and (_02825_, _02824_, _42355_);
  and (_38958_, _02825_, _02823_);
  and (_02827_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_02828_, _02827_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02829_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01922_);
  and (_02830_, _02829_, _42355_);
  and (_38959_, _02830_, _02828_);
  and (_02832_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_02833_, _02832_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02835_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01922_);
  and (_02836_, _02835_, _42355_);
  and (_38960_, _02836_, _02833_);
  and (_02837_, _01929_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_02838_, _02837_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02840_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01922_);
  and (_02841_, _02840_, _42355_);
  and (_38961_, _02841_, _02838_);
  nand (_02843_, _01936_, _32444_);
  or (_02844_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02846_, _02844_, _42355_);
  and (_38962_, _02846_, _02843_);
  nand (_02847_, _01936_, _33119_);
  or (_02849_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02850_, _02849_, _42355_);
  and (_38963_, _02850_, _02847_);
  nand (_02853_, _01936_, _33837_);
  or (_02854_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_02855_, _02854_, _42355_);
  and (_38965_, _02855_, _02853_);
  not (_02857_, _01936_);
  or (_02858_, _02857_, _34566_);
  or (_02860_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_02861_, _02860_, _42355_);
  and (_38966_, _02861_, _02858_);
  or (_02863_, _02857_, _35229_);
  or (_02864_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_02866_, _02864_, _42355_);
  and (_38967_, _02866_, _02863_);
  nand (_02867_, _01936_, _36025_);
  or (_02868_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_02869_, _02868_, _42355_);
  and (_38968_, _02869_, _02867_);
  nand (_02870_, _01936_, _36752_);
  or (_02872_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_02874_, _02872_, _42355_);
  and (_38969_, _02874_, _02870_);
  nand (_02876_, _01936_, _31234_);
  or (_02877_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_02878_, _02877_, _42355_);
  and (_38970_, _02878_, _02876_);
  nand (_02880_, _01936_, _38137_);
  or (_02881_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_02883_, _02881_, _42355_);
  and (_38971_, _02883_, _02880_);
  nand (_02885_, _01936_, _38168_);
  or (_02887_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_02888_, _02887_, _42355_);
  and (_38972_, _02888_, _02885_);
  nand (_02890_, _01936_, _38198_);
  or (_02891_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_02892_, _02891_, _42355_);
  and (_38973_, _02892_, _02890_);
  or (_02894_, _02857_, _38226_);
  or (_02896_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_02898_, _02896_, _42355_);
  and (_38974_, _02898_, _02894_);
  or (_02899_, _02857_, _38256_);
  or (_02900_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_02902_, _02900_, _42355_);
  and (_38976_, _02902_, _02899_);
  nand (_02903_, _01936_, _38291_);
  or (_02905_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_02906_, _02905_, _42355_);
  and (_38977_, _02906_, _02903_);
  or (_02908_, _02857_, _38317_);
  or (_02909_, _01936_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_02910_, _02909_, _42355_);
  and (_38978_, _02910_, _02908_);
  nor (_39196_, _41844_, rst);
  and (_02912_, _41797_, _37879_);
  and (_02914_, _02912_, _38522_);
  and (_02915_, _02914_, _41799_);
  nand (_02916_, _02915_, _37963_);
  or (_02918_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02920_, _02918_, _42355_);
  and (_39197_, _02920_, _02916_);
  and (_02922_, _02912_, _38746_);
  not (_02923_, _02922_);
  nor (_02925_, _02923_, _37963_);
  not (_02926_, _41799_);
  and (_02927_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_02928_, _02927_, _02926_);
  or (_02929_, _02928_, _02925_);
  or (_02930_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02932_, _02930_, _42355_);
  and (_39198_, _02932_, _02929_);
  and (_02934_, _27633_, _28301_);
  and (_02935_, _02912_, _02934_);
  and (_02937_, _02935_, _41799_);
  nand (_02938_, _02937_, _37963_);
  or (_02939_, _02937_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_02941_, _02939_, _42355_);
  and (_39199_, _02941_, _02938_);
  and (_02942_, _02912_, _40897_);
  and (_02945_, _02942_, _41799_);
  not (_02946_, _02945_);
  nor (_02947_, _02946_, _37963_);
  and (_02949_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_02950_, _02949_, _02947_);
  and (_39201_, _02950_, _42355_);
  nor (_02952_, _02922_, _02914_);
  not (_02953_, _02935_);
  and (_02954_, _02953_, _02952_);
  and (_02956_, _41797_, _38361_);
  and (_02958_, _02956_, _38522_);
  nor (_02960_, _02958_, _02942_);
  and (_02961_, _02960_, _02954_);
  nand (_02962_, _02954_, _41799_);
  or (_02963_, _02962_, _02942_);
  or (_02965_, _02963_, _02961_);
  and (_02966_, _02965_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_02967_, _02958_, _41799_);
  not (_02969_, _02967_);
  nor (_02970_, _02969_, _37963_);
  or (_02972_, _02970_, _02966_);
  and (_39202_, _02972_, _42355_);
  and (_02974_, _02956_, _38746_);
  not (_02975_, _02974_);
  and (_02977_, _02975_, _02960_);
  and (_02978_, _02977_, _02954_);
  nand (_02979_, _02960_, _02953_);
  and (_02981_, _02979_, _41799_);
  nand (_02982_, _02952_, _41799_);
  or (_02983_, _02982_, _02981_);
  or (_02986_, _02983_, _02978_);
  and (_02987_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_02988_, _02974_, _41799_);
  and (_02990_, _02988_, _40030_);
  or (_02991_, _02990_, _02987_);
  and (_39203_, _02991_, _42355_);
  and (_02993_, _02956_, _02934_);
  and (_02994_, _02993_, _41799_);
  not (_02995_, _02994_);
  nor (_02997_, _02995_, _37963_);
  and (_02999_, _02995_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_03000_, _02999_, _02997_);
  and (_39204_, _03000_, _42355_);
  and (_03002_, _02956_, _40897_);
  not (_03003_, _03002_);
  nor (_03005_, _03003_, _37963_);
  and (_03006_, _03003_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_03007_, _03006_, _02926_);
  or (_03009_, _03007_, _03005_);
  or (_03010_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_03012_, _03010_, _42355_);
  and (_39205_, _03012_, _03009_);
  nand (_03014_, _02915_, _37941_);
  or (_03015_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03017_, _03015_, _42355_);
  and (_39294_, _03017_, _03014_);
  nand (_03018_, _02915_, _37934_);
  or (_03020_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03021_, _03020_, _42355_);
  and (_39295_, _03021_, _03018_);
  nand (_03024_, _02915_, _37927_);
  or (_03025_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_03026_, _03025_, _42355_);
  and (_39296_, _03026_, _03024_);
  nand (_03028_, _02915_, _37920_);
  or (_03029_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_03031_, _03029_, _42355_);
  and (_39297_, _03031_, _03028_);
  nand (_03032_, _02915_, _37912_);
  or (_03034_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_03035_, _03034_, _42355_);
  and (_39298_, _03035_, _03032_);
  nand (_03037_, _02915_, _37904_);
  or (_03038_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03039_, _03038_, _42355_);
  and (_39299_, _03039_, _03037_);
  nand (_03041_, _02915_, _37896_);
  or (_03042_, _02915_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03044_, _03042_, _42355_);
  and (_39300_, _03044_, _03041_);
  and (_03045_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_03047_, _02923_, _37941_);
  or (_03048_, _03047_, _02926_);
  or (_03050_, _03048_, _03045_);
  or (_03051_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_03052_, _03051_, _42355_);
  and (_39301_, _03052_, _03050_);
  nor (_03053_, _02923_, _37934_);
  and (_03054_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_03055_, _03054_, _02926_);
  or (_03057_, _03055_, _03053_);
  or (_03058_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03059_, _03058_, _42355_);
  and (_39302_, _03059_, _03057_);
  nor (_03061_, _02923_, _37927_);
  and (_03062_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03064_, _03062_, _02926_);
  or (_03065_, _03064_, _03061_);
  or (_03066_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03068_, _03066_, _42355_);
  and (_39303_, _03068_, _03065_);
  nor (_03069_, _02923_, _37920_);
  and (_03071_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03072_, _03071_, _02926_);
  or (_03073_, _03072_, _03069_);
  or (_03075_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03076_, _03075_, _42355_);
  and (_39305_, _03076_, _03073_);
  nor (_03078_, _02923_, _37912_);
  and (_03079_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_03081_, _03079_, _02926_);
  or (_03082_, _03081_, _03078_);
  or (_03083_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_03084_, _03083_, _42355_);
  and (_39306_, _03084_, _03082_);
  nor (_03086_, _02923_, _37904_);
  and (_03087_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_03089_, _03087_, _02926_);
  or (_03090_, _03089_, _03086_);
  or (_03091_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_03093_, _03091_, _42355_);
  and (_39307_, _03093_, _03090_);
  nor (_03094_, _02923_, _37896_);
  and (_03096_, _02923_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03097_, _03096_, _02926_);
  or (_03098_, _03097_, _03094_);
  or (_03100_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03101_, _03100_, _42355_);
  and (_39308_, _03101_, _03098_);
  nand (_03103_, _02937_, _37941_);
  or (_03104_, _02937_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_03105_, _03104_, _42355_);
  and (_39309_, _03105_, _03103_);
  not (_03107_, _02937_);
  nor (_03109_, _03107_, _37934_);
  nor (_03110_, _02954_, _02926_);
  nand (_03111_, _03110_, _02952_);
  and (_03112_, _03111_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_03114_, _03112_, _03109_);
  and (_39310_, _03114_, _42355_);
  nor (_03115_, _03107_, _37927_);
  and (_03117_, _03111_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_03118_, _03117_, _03115_);
  and (_39311_, _03118_, _42355_);
  nor (_03120_, _03107_, _37920_);
  and (_03121_, _03111_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_03122_, _03121_, _03120_);
  and (_39312_, _03122_, _42355_);
  nand (_03124_, _02937_, _37912_);
  or (_03125_, _02937_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_03128_, _03125_, _42355_);
  and (_39313_, _03128_, _03124_);
  nor (_03129_, _03107_, _37904_);
  and (_03131_, _03111_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_03132_, _03131_, _03129_);
  and (_39314_, _03132_, _42355_);
  nor (_03134_, _03107_, _37896_);
  and (_03135_, _03111_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_03137_, _03135_, _03134_);
  and (_39316_, _03137_, _42355_);
  and (_03138_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_03139_, _02945_, _37942_);
  or (_03141_, _03139_, _03138_);
  and (_39317_, _03141_, _42355_);
  and (_03142_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_03144_, _02946_, _37934_);
  or (_03145_, _03144_, _03142_);
  and (_39318_, _03145_, _42355_);
  nor (_03147_, _02946_, _37927_);
  and (_03148_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_03149_, _03148_, _03147_);
  and (_39319_, _03149_, _42355_);
  nor (_03151_, _02946_, _37920_);
  and (_03152_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_03154_, _03152_, _03151_);
  and (_39320_, _03154_, _42355_);
  and (_03155_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_03157_, _02946_, _37912_);
  or (_03158_, _03157_, _03155_);
  and (_39321_, _03158_, _42355_);
  nor (_03160_, _02946_, _37904_);
  and (_03161_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_03163_, _03161_, _03160_);
  and (_39322_, _03163_, _42355_);
  nor (_03164_, _02946_, _37896_);
  and (_03165_, _02946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03166_, _03165_, _03164_);
  and (_39323_, _03166_, _42355_);
  and (_03168_, _02965_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_03169_, _02967_, _37942_);
  or (_03171_, _03169_, _03168_);
  and (_39324_, _03171_, _42355_);
  nor (_03172_, _02969_, _37934_);
  and (_03174_, _02969_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or (_03175_, _03174_, _03172_);
  and (_39325_, _03175_, _42355_);
  nor (_03177_, _02969_, _37927_);
  and (_03178_, _02965_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_03179_, _03178_, _03177_);
  and (_39327_, _03179_, _42355_);
  nor (_03181_, _02969_, _37920_);
  and (_03182_, _02965_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_03184_, _03182_, _03181_);
  and (_39328_, _03184_, _42355_);
  and (_03185_, _02969_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_03187_, _02969_, _37912_);
  or (_03188_, _03187_, _03185_);
  and (_39329_, _03188_, _42355_);
  nor (_03190_, _02969_, _37904_);
  and (_03191_, _02969_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_03192_, _03191_, _03190_);
  and (_39330_, _03192_, _42355_);
  nor (_03194_, _02969_, _37896_);
  and (_03195_, _02965_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_03197_, _03195_, _03194_);
  and (_39331_, _03197_, _42355_);
  and (_03198_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_03200_, _02926_, _37941_);
  and (_03201_, _03200_, _02974_);
  or (_03202_, _03201_, _03198_);
  and (_39332_, _03202_, _42355_);
  and (_03204_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_03205_, _02988_, _40709_);
  or (_03207_, _03205_, _03204_);
  and (_39333_, _03207_, _42355_);
  and (_03208_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  not (_03210_, _37927_);
  and (_03211_, _02988_, _03210_);
  or (_03212_, _03211_, _03208_);
  and (_39334_, _03212_, _42355_);
  and (_03214_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_03216_, _02988_, _40726_);
  or (_03217_, _03216_, _03214_);
  and (_39335_, _03217_, _42355_);
  and (_03218_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_03220_, _02988_, _40734_);
  or (_03221_, _03220_, _03218_);
  and (_39336_, _03221_, _42355_);
  and (_03223_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03224_, _02988_, _40742_);
  or (_03225_, _03224_, _03223_);
  and (_39338_, _03225_, _42355_);
  and (_03227_, _02986_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_03228_, _02988_, _41687_);
  or (_03230_, _03228_, _03227_);
  and (_39339_, _03230_, _42355_);
  not (_03231_, _02993_);
  and (_03233_, _03231_, _02978_);
  or (_03234_, _03233_, _02962_);
  and (_03235_, _03234_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_03237_, _02994_, _37942_);
  nand (_03238_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_03239_, _03238_, _02977_);
  or (_03241_, _03239_, _03237_);
  or (_03242_, _03241_, _03235_);
  and (_39340_, _03242_, _42355_);
  and (_03244_, _03234_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03245_, _02995_, _37934_);
  nand (_03246_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03248_, _03246_, _02977_);
  or (_03249_, _03248_, _03245_);
  or (_03250_, _03249_, _03244_);
  and (_39341_, _03250_, _42355_);
  and (_03252_, _02995_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_03253_, _02995_, _37927_);
  or (_03255_, _03253_, _03252_);
  and (_39342_, _03255_, _42355_);
  nor (_03256_, _02995_, _37920_);
  nor (_03258_, _02977_, _02926_);
  or (_03259_, _03258_, _03234_);
  and (_03260_, _03259_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or (_03262_, _03260_, _03256_);
  and (_39343_, _03262_, _42355_);
  and (_03263_, _02995_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_03265_, _02995_, _37912_);
  or (_03266_, _03265_, _03263_);
  and (_39344_, _03266_, _42355_);
  nor (_03268_, _02995_, _37904_);
  and (_03269_, _03259_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_03270_, _03269_, _03268_);
  and (_39345_, _03270_, _42355_);
  nor (_03271_, _02995_, _37896_);
  and (_03272_, _03259_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_03273_, _03272_, _03271_);
  and (_39346_, _03273_, _42355_);
  and (_03274_, _03003_, _03233_);
  or (_03275_, _03274_, _02963_);
  or (_03276_, _38746_, _27633_);
  and (_03277_, _03276_, _02956_);
  and (_03278_, _03277_, _41799_);
  or (_03279_, _03278_, _03275_);
  and (_03280_, _03279_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03281_, _03200_, _03002_);
  or (_03282_, _03281_, _03280_);
  and (_39347_, _03282_, _42355_);
  and (_03283_, _03003_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_03284_, _03003_, _37934_);
  or (_03285_, _03284_, _02926_);
  or (_03286_, _03285_, _03283_);
  or (_03287_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_03288_, _03287_, _42355_);
  and (_39349_, _03288_, _03286_);
  and (_03289_, _03003_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_03290_, _03003_, _37927_);
  or (_03291_, _03290_, _03289_);
  or (_03292_, _03291_, _02926_);
  or (_03293_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_03294_, _03293_, _42355_);
  and (_39350_, _03294_, _03292_);
  and (_03295_, _03275_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_03296_, _03003_, _37920_);
  and (_03297_, _03277_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or (_03298_, _03297_, _03296_);
  and (_03299_, _03298_, _41799_);
  or (_03300_, _03299_, _03295_);
  and (_39351_, _03300_, _42355_);
  nor (_03301_, _03003_, _37912_);
  nand (_03302_, _03002_, _41799_);
  and (_03303_, _03302_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_03304_, _03303_, _03301_);
  or (_03305_, _41799_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_03306_, _03305_, _42355_);
  and (_39352_, _03306_, _03304_);
  and (_03307_, _03275_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_03308_, _03003_, _37904_);
  and (_03309_, _03277_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  or (_03310_, _03309_, _03308_);
  and (_03311_, _03310_, _41799_);
  or (_03312_, _03311_, _03307_);
  and (_39353_, _03312_, _42355_);
  and (_03313_, _03275_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_03314_, _03003_, _37896_);
  and (_03315_, _03277_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_03316_, _03315_, _03314_);
  and (_03317_, _03316_, _41799_);
  or (_03318_, _03317_, _03313_);
  and (_39354_, _03318_, _42355_);
  not (_03319_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03320_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_03321_, _03320_, _03319_);
  and (_03322_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _42355_);
  and (_39418_, _03322_, _03321_);
  nor (_03323_, _03321_, rst);
  nand (_03324_, _03320_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03325_, _03320_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03326_, _03325_, _03324_);
  and (_39420_, _03326_, _03323_);
  and (_03327_, _01357_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not (_03328_, _42088_);
  and (_03329_, _03328_, _42138_);
  not (_03331_, _41829_);
  and (_03332_, _41894_, _03331_);
  and (_03333_, _03332_, _03329_);
  and (_03334_, _03333_, _41995_);
  nor (_03335_, _42037_, _41939_);
  not (_03336_, _42180_);
  and (_03337_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03338_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_03339_, _03338_, _03337_);
  and (_03340_, _03339_, _03335_);
  or (_03341_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03342_, _42037_, _41939_);
  nand (_03343_, _42180_, _41317_);
  and (_03344_, _03343_, _03342_);
  and (_03345_, _03344_, _03341_);
  not (_03346_, _42037_);
  nor (_03347_, _03346_, _41939_);
  and (_03348_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_03349_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03350_, _03349_, _03348_);
  and (_03351_, _03350_, _03347_);
  or (_03352_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_03353_, _03346_, _41939_);
  nand (_03354_, _42180_, _41284_);
  and (_03355_, _03354_, _03353_);
  and (_03356_, _03355_, _03352_);
  or (_03357_, _03356_, _03351_);
  or (_03358_, _03357_, _03345_);
  or (_03359_, _03358_, _03340_);
  and (_03360_, _03359_, _03334_);
  and (_03361_, _03332_, _41995_);
  and (_03362_, _42088_, _42138_);
  and (_03363_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03364_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_03365_, _03364_, _03363_);
  and (_03366_, _03365_, _03335_);
  or (_03367_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand (_03368_, _42180_, _40135_);
  and (_03369_, _03368_, _03342_);
  and (_03370_, _03369_, _03367_);
  or (_03371_, _03370_, _03366_);
  and (_03372_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03373_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03374_, _03373_, _03372_);
  and (_03375_, _03374_, _03347_);
  or (_03376_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03377_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_03378_, _03377_, _03353_);
  and (_03379_, _03378_, _03376_);
  or (_03380_, _03379_, _03375_);
  or (_03381_, _03380_, _03371_);
  and (_03382_, _03381_, _03362_);
  nor (_03383_, _03328_, _42138_);
  nor (_03384_, _42180_, _40177_);
  and (_03385_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03386_, _03385_, _03384_);
  and (_03387_, _03386_, _03342_);
  or (_03388_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03389_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03390_, _03389_, _03335_);
  and (_03391_, _03390_, _03388_);
  or (_03392_, _03391_, _03387_);
  and (_03393_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03394_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03395_, _03394_, _03393_);
  and (_03396_, _03395_, _03347_);
  or (_03397_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_03398_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03399_, _03398_, _03353_);
  and (_03400_, _03399_, _03397_);
  or (_03401_, _03400_, _03396_);
  or (_03402_, _03401_, _03392_);
  and (_03403_, _03402_, _03383_);
  or (_03404_, _03403_, _03382_);
  and (_03405_, _03404_, _03361_);
  or (_03406_, _03405_, _03360_);
  and (_03407_, _03342_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03408_, _03407_, _03336_);
  and (_03409_, _03335_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03410_, _03353_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03411_, _03347_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03412_, _03411_, _03410_);
  or (_03413_, _03412_, _03409_);
  or (_03414_, _03413_, _03408_);
  nor (_03415_, _42088_, _42138_);
  and (_03416_, _03415_, _03332_);
  and (_03417_, _03416_, _41994_);
  and (_03418_, _03342_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03419_, _03418_, _42180_);
  and (_03420_, _03335_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03421_, _03353_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03422_, _03347_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03423_, _03422_, _03421_);
  or (_03424_, _03423_, _03420_);
  or (_03425_, _03424_, _03419_);
  and (_03426_, _03425_, _03417_);
  and (_03427_, _03426_, _03414_);
  nor (_03428_, _00924_, _01077_);
  and (_03429_, _37803_, _37725_);
  or (_03430_, _03429_, _37821_);
  nor (_03431_, _03430_, _37843_);
  and (_03432_, _03431_, _00826_);
  or (_03433_, _00939_, _00763_);
  nor (_03434_, _03433_, _00824_);
  or (_03435_, _37824_, _37816_);
  nor (_03436_, _03435_, _00761_);
  and (_03437_, _03436_, _03434_);
  and (_03438_, _03437_, _03432_);
  and (_03439_, _03438_, _37773_);
  and (_03440_, _03439_, _03428_);
  nor (_03441_, _03440_, _36982_);
  or (_03442_, _03441_, p1_in[1]);
  not (_03443_, _03441_);
  or (_03444_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03445_, _03444_, _03442_);
  and (_03446_, _03445_, _03353_);
  nor (_03447_, _03441_, p1_in[0]);
  and (_03448_, _03441_, _39029_);
  nor (_03449_, _03448_, _03447_);
  and (_03450_, _03449_, _03342_);
  or (_03451_, _03450_, _03446_);
  or (_03452_, _03441_, p1_in[3]);
  or (_03453_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03454_, _03453_, _03452_);
  and (_03455_, _03454_, _03335_);
  or (_03456_, _03441_, p1_in[2]);
  or (_03457_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03458_, _03457_, _03456_);
  and (_03459_, _03458_, _03347_);
  or (_03460_, _03459_, _03455_);
  or (_03461_, _03460_, _03451_);
  and (_03462_, _03461_, _42180_);
  or (_03463_, _03441_, p1_in[5]);
  or (_03464_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03465_, _03464_, _03463_);
  and (_03466_, _03465_, _03353_);
  or (_03467_, _03441_, p1_in[4]);
  or (_03468_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03469_, _03468_, _03467_);
  and (_03470_, _03469_, _03342_);
  or (_03471_, _03470_, _03466_);
  or (_03472_, _03441_, p1_in[7]);
  or (_03473_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03474_, _03473_, _03472_);
  and (_03475_, _03474_, _03335_);
  or (_03476_, _03441_, p1_in[6]);
  or (_03477_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03478_, _03477_, _03476_);
  and (_03479_, _03478_, _03347_);
  or (_03480_, _03479_, _03475_);
  or (_03481_, _03480_, _03471_);
  and (_03482_, _03481_, _03336_);
  or (_03483_, _03482_, _03462_);
  nor (_03484_, _41995_, _41894_);
  and (_03485_, _03484_, _03331_);
  and (_03486_, _03362_, _03485_);
  and (_03487_, _03486_, _03483_);
  and (_03488_, _03332_, _03362_);
  and (_03489_, _03488_, _41994_);
  or (_03490_, _03441_, p0_in[7]);
  or (_03491_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03492_, _03491_, _03490_);
  and (_03493_, _03492_, _03336_);
  or (_03494_, _03441_, p0_in[3]);
  or (_03495_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03496_, _03495_, _03494_);
  and (_03497_, _03496_, _42180_);
  or (_03498_, _03497_, _03493_);
  and (_03499_, _03498_, _03335_);
  nor (_03500_, _03441_, p0_in[0]);
  and (_03501_, _03441_, _38742_);
  nor (_03502_, _03501_, _03500_);
  or (_03503_, _03502_, _03336_);
  or (_03504_, _03441_, p0_in[4]);
  or (_03505_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03506_, _03505_, _03504_);
  or (_03507_, _03506_, _42180_);
  and (_03508_, _03507_, _03342_);
  and (_03509_, _03508_, _03503_);
  or (_03510_, _03441_, p0_in[6]);
  or (_03511_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03512_, _03511_, _03510_);
  and (_03513_, _03512_, _03336_);
  or (_03514_, _03441_, p0_in[2]);
  or (_03515_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03516_, _03515_, _03514_);
  and (_03517_, _03516_, _42180_);
  or (_03518_, _03517_, _03513_);
  and (_03519_, _03518_, _03347_);
  or (_03520_, _03441_, p0_in[1]);
  or (_03521_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03522_, _03521_, _03520_);
  or (_03523_, _03522_, _03336_);
  or (_03524_, _03441_, p0_in[5]);
  or (_03525_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03526_, _03525_, _03524_);
  or (_03527_, _03526_, _42180_);
  and (_03528_, _03527_, _03353_);
  and (_03529_, _03528_, _03523_);
  or (_03530_, _03529_, _03519_);
  or (_03532_, _03530_, _03509_);
  or (_03533_, _03532_, _03499_);
  and (_03534_, _03533_, _03489_);
  and (_03535_, _42088_, _03331_);
  nand (_03536_, _03535_, _41995_);
  nor (_03537_, _03485_, _29200_);
  nand (_03538_, _03537_, _03536_);
  nor (_03539_, _03538_, _03489_);
  and (_03540_, _03383_, _03332_);
  and (_03541_, _03540_, _41994_);
  or (_03542_, _03417_, _03541_);
  nor (_03543_, _03542_, _03334_);
  and (_03544_, _03543_, _03539_);
  or (_03545_, _03544_, _03534_);
  or (_03546_, _03545_, _03487_);
  or (_03547_, _03546_, _03427_);
  or (_03548_, _03547_, _03406_);
  and (_03549_, _03485_, _03329_);
  not (_03550_, _38618_);
  and (_03551_, _38630_, _03550_);
  nor (_03552_, _38630_, _03550_);
  nor (_03553_, _03552_, _03551_);
  nor (_03554_, _38606_, _38595_);
  and (_03555_, _38606_, _38595_);
  nor (_03556_, _03555_, _03554_);
  nor (_03557_, _03556_, _03553_);
  and (_03558_, _03556_, _03553_);
  or (_03559_, _03558_, _03557_);
  and (_03560_, _38667_, _38547_);
  nor (_03561_, _38667_, _38547_);
  or (_03562_, _03561_, _03560_);
  not (_03563_, _38652_);
  and (_03564_, _03563_, _38640_);
  nor (_03565_, _03563_, _38640_);
  nor (_03566_, _03565_, _03564_);
  and (_03567_, _03566_, _03562_);
  nor (_03568_, _03566_, _03562_);
  or (_03569_, _03568_, _03567_);
  nor (_03570_, _03569_, _03559_);
  and (_03571_, _03569_, _03559_);
  nor (_03572_, _03571_, _03570_);
  nand (_03573_, _03572_, _42180_);
  or (_03574_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03575_, _03574_, _03342_);
  and (_03576_, _03575_, _03573_);
  nor (_03577_, _42180_, _38351_);
  and (_03578_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03579_, _03578_, _03577_);
  and (_03580_, _03579_, _03335_);
  or (_03581_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_03582_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03583_, _03582_, _03353_);
  and (_03584_, _03583_, _03581_);
  or (_03585_, _03584_, _03580_);
  or (_03586_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03587_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_03588_, _03587_, _03347_);
  and (_03589_, _03588_, _03586_);
  or (_03590_, _03589_, _03585_);
  or (_03591_, _03590_, _03576_);
  and (_03592_, _03591_, _03549_);
  and (_03593_, _03383_, _03485_);
  or (_03594_, _03441_, p3_in[7]);
  or (_03595_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03596_, _03595_, _03594_);
  and (_03597_, _03596_, _03336_);
  or (_03598_, _03441_, p3_in[3]);
  or (_03599_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03600_, _03599_, _03598_);
  and (_03601_, _03600_, _42180_);
  or (_03602_, _03601_, _03597_);
  and (_03603_, _03602_, _03335_);
  nor (_03604_, _03441_, p3_in[0]);
  and (_03605_, _03441_, _39195_);
  nor (_03606_, _03605_, _03604_);
  or (_03607_, _03606_, _03336_);
  or (_03608_, _03441_, p3_in[4]);
  or (_03609_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03610_, _03609_, _03608_);
  or (_03611_, _03610_, _42180_);
  and (_03612_, _03611_, _03342_);
  and (_03613_, _03612_, _03607_);
  or (_03614_, _03613_, _03603_);
  or (_03615_, _03441_, p3_in[6]);
  or (_03616_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03617_, _03616_, _03615_);
  and (_03618_, _03617_, _03336_);
  or (_03619_, _03441_, p3_in[2]);
  or (_03620_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03621_, _03620_, _03619_);
  and (_03622_, _03621_, _42180_);
  or (_03623_, _03622_, _03618_);
  and (_03624_, _03623_, _03347_);
  or (_03625_, _03441_, p3_in[1]);
  or (_03626_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03627_, _03626_, _03625_);
  or (_03628_, _03627_, _03336_);
  or (_03629_, _03441_, p3_in[5]);
  or (_03630_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03631_, _03630_, _03629_);
  or (_03632_, _03631_, _42180_);
  and (_03633_, _03632_, _03353_);
  and (_03634_, _03633_, _03628_);
  or (_03635_, _03634_, _03624_);
  or (_03636_, _03635_, _03614_);
  and (_03637_, _03636_, _03593_);
  or (_03638_, _41994_, _41829_);
  nor (_03639_, _03638_, _41894_);
  and (_03640_, _03383_, _03639_);
  and (_03641_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03642_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03643_, _03642_, _03641_);
  and (_03644_, _03643_, _03335_);
  or (_03645_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nand (_03646_, _42180_, _40196_);
  and (_03647_, _03646_, _03342_);
  and (_03648_, _03647_, _03645_);
  or (_03649_, _03648_, _03644_);
  and (_03650_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03651_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03652_, _03651_, _03650_);
  and (_03653_, _03652_, _03347_);
  or (_03654_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  nand (_03655_, _42180_, _40199_);
  and (_03656_, _03655_, _03353_);
  and (_03657_, _03656_, _03654_);
  or (_03658_, _03657_, _03653_);
  or (_03659_, _03658_, _03649_);
  and (_03660_, _03659_, _03640_);
  and (_03661_, _03415_, _03485_);
  nor (_03662_, _42180_, _31321_);
  and (_03663_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03664_, _03663_, _03662_);
  and (_03665_, _03664_, _03335_);
  or (_03666_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_03667_, _42180_, _32477_);
  and (_03668_, _03667_, _03342_);
  and (_03669_, _03668_, _03666_);
  or (_03670_, _03669_, _03665_);
  nor (_03671_, _42180_, _36057_);
  and (_03672_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03673_, _03672_, _03671_);
  and (_03674_, _03673_, _03353_);
  nand (_03675_, _42180_, _33870_);
  or (_03676_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03677_, _03676_, _03347_);
  and (_03678_, _03677_, _03675_);
  or (_03679_, _03678_, _03674_);
  or (_03680_, _03679_, _03670_);
  and (_03681_, _03680_, _03661_);
  or (_03682_, _03681_, _03660_);
  or (_03683_, _03682_, _03637_);
  nor (_03684_, _42180_, _40756_);
  and (_03685_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03686_, _03685_, _03684_);
  and (_03687_, _03686_, _03335_);
  or (_03688_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand (_03689_, _42180_, _40773_);
  and (_03690_, _03689_, _03342_);
  and (_03691_, _03690_, _03688_);
  or (_03692_, _03691_, _03687_);
  and (_03693_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03694_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03695_, _03694_, _03693_);
  and (_03696_, _03695_, _03347_);
  or (_03697_, _42180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_03698_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_03699_, _03698_, _03353_);
  and (_03700_, _03699_, _03697_);
  or (_03701_, _03700_, _03696_);
  or (_03702_, _03701_, _03692_);
  and (_03703_, _03639_, _03362_);
  and (_03704_, _03703_, _03702_);
  or (_03705_, _03441_, p2_in[1]);
  or (_03706_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03707_, _03706_, _03705_);
  or (_03708_, _03707_, _03336_);
  or (_03709_, _03441_, p2_in[5]);
  or (_03710_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03711_, _03710_, _03709_);
  or (_03712_, _03711_, _42180_);
  and (_03713_, _03712_, _03353_);
  and (_03714_, _03713_, _03708_);
  or (_03715_, _03441_, p2_in[2]);
  or (_03716_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03717_, _03716_, _03715_);
  or (_03718_, _03717_, _03336_);
  or (_03719_, _03441_, p2_in[6]);
  or (_03720_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03721_, _03720_, _03719_);
  or (_03722_, _03721_, _42180_);
  and (_03723_, _03722_, _03347_);
  and (_03724_, _03723_, _03718_);
  nor (_03725_, _03441_, p2_in[0]);
  and (_03726_, _03441_, _39110_);
  nor (_03727_, _03726_, _03725_);
  or (_03728_, _03727_, _03336_);
  or (_03729_, _03441_, p2_in[4]);
  or (_03730_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03731_, _03730_, _03729_);
  or (_03733_, _03731_, _42180_);
  and (_03734_, _03733_, _03342_);
  and (_03735_, _03734_, _03728_);
  or (_03736_, _03441_, p2_in[3]);
  or (_03737_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03738_, _03737_, _03736_);
  or (_03739_, _03738_, _03336_);
  or (_03740_, _03441_, p2_in[7]);
  or (_03741_, _03443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03742_, _03741_, _03740_);
  or (_03743_, _03742_, _42180_);
  and (_03744_, _03743_, _03335_);
  and (_03745_, _03744_, _03739_);
  or (_03746_, _03745_, _03735_);
  or (_03747_, _03746_, _03724_);
  or (_03748_, _03747_, _03714_);
  and (_03749_, _03748_, _03541_);
  or (_03750_, _03749_, _03704_);
  or (_03751_, _03750_, _03683_);
  or (_03752_, _03751_, _03592_);
  or (_03753_, _03752_, _03548_);
  or (_03754_, _03753_, _03327_);
  and (_03755_, _03417_, _38521_);
  nor (_03756_, _03755_, _01363_);
  nand (_03757_, _03327_, _31889_);
  and (_03758_, _03757_, _03756_);
  and (_03759_, _03758_, _03754_);
  nand (_03760_, _42180_, _37934_);
  or (_03761_, _42180_, _40742_);
  and (_03762_, _03761_, _03353_);
  and (_03763_, _03762_, _03760_);
  nor (_03764_, _42180_, _37963_);
  and (_03765_, _42180_, _40726_);
  or (_03766_, _03765_, _03764_);
  and (_03767_, _03766_, _03335_);
  nor (_03768_, _42180_, _37912_);
  and (_03769_, _42180_, _37942_);
  or (_03770_, _03769_, _03768_);
  and (_03771_, _03770_, _03342_);
  or (_03772_, _03771_, _03767_);
  or (_03773_, _42180_, _41687_);
  nand (_03774_, _42180_, _37927_);
  and (_03775_, _03774_, _03347_);
  and (_03776_, _03775_, _03773_);
  or (_03777_, _03776_, _03772_);
  nor (_03778_, _03777_, _03763_);
  nor (_03779_, _03778_, _03756_);
  or (_03780_, _03779_, _03759_);
  and (_39421_, _03780_, _42355_);
  and (_03781_, _42138_, _41895_);
  nor (_03782_, _42088_, _41829_);
  and (_03783_, _41994_, _42180_);
  and (_03784_, _03783_, _03342_);
  and (_03785_, _03784_, _03782_);
  and (_03786_, _03785_, _03781_);
  and (_03787_, _03786_, _38356_);
  and (_03788_, _03488_, _03335_);
  and (_03789_, _03788_, _03783_);
  and (_03790_, _03789_, _38011_);
  nor (_03791_, _03790_, _03787_);
  nor (_03792_, _03791_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_03793_, _03792_);
  and (_03794_, _03784_, _03416_);
  and (_03795_, _03794_, _38538_);
  not (_03796_, _38532_);
  and (_03797_, _03335_, _03336_);
  nor (_03798_, _03797_, _03796_);
  and (_03799_, _03798_, _01344_);
  nor (_03800_, _03799_, _03795_);
  and (_03801_, _03800_, _01360_);
  and (_03802_, _03801_, _03793_);
  and (_03803_, _03783_, _03347_);
  and (_03804_, _03803_, _03488_);
  and (_03805_, _03804_, _38011_);
  or (_03806_, _03805_, rst);
  nor (_39422_, _03806_, _03802_);
  nand (_03807_, _03805_, _31234_);
  and (_03808_, _41995_, _42180_);
  and (_03809_, _03808_, _03342_);
  and (_03810_, _03809_, _03333_);
  and (_03811_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_03812_, _41994_, _42180_);
  and (_03813_, _03812_, _03342_);
  and (_03814_, _03813_, _03333_);
  and (_03815_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_03816_, _03815_, _03811_);
  and (_03817_, _03808_, _03347_);
  and (_03818_, _03817_, _03333_);
  and (_03819_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_03820_, _03812_, _03353_);
  and (_03821_, _03820_, _03333_);
  and (_03822_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_03823_, _03822_, _03819_);
  or (_03824_, _03823_, _03816_);
  and (_03825_, _03808_, _03335_);
  and (_03826_, _03825_, _03333_);
  and (_03827_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_03828_, _03809_, _03488_);
  and (_03829_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03830_, _03829_, _03827_);
  and (_03831_, _03809_, _03540_);
  and (_03832_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03833_, _03797_, _41994_);
  nor (_03834_, _42138_, _41894_);
  and (_03835_, _03834_, _03535_);
  and (_03836_, _03835_, _03833_);
  and (_03837_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03838_, _03837_, _03832_);
  or (_03839_, _03838_, _03830_);
  or (_03840_, _03839_, _03824_);
  and (_03841_, _03825_, _03488_);
  and (_03842_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_03843_, _03808_, _03353_);
  and (_03844_, _03843_, _03488_);
  and (_03845_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_03846_, _03845_, _03842_);
  and (_03847_, _03820_, _03488_);
  and (_03848_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_03849_, _03817_, _03488_);
  and (_03850_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_03851_, _03850_, _03848_);
  or (_03852_, _03851_, _03846_);
  and (_03853_, _03781_, _03535_);
  and (_03854_, _03843_, _03853_);
  and (_03855_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03856_, _03853_, _03809_);
  and (_03857_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03858_, _03857_, _03855_);
  and (_03859_, _03813_, _03488_);
  and (_03860_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03861_, _03797_, _03489_);
  and (_03862_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03863_, _03862_, _03860_);
  or (_03864_, _03863_, _03858_);
  or (_03865_, _03864_, _03852_);
  or (_03866_, _03865_, _03840_);
  and (_03867_, _03488_, _03353_);
  and (_03868_, _03867_, _03783_);
  and (_03869_, _03868_, _37965_);
  and (_03870_, _03834_, _03785_);
  and (_03871_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_03872_, _03871_, _03869_);
  and (_03873_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_03874_, _03783_, _03335_);
  and (_03875_, _03874_, _03488_);
  and (_03876_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_03877_, _03876_, _03873_);
  or (_03878_, _03877_, _03872_);
  and (_03879_, _03853_, _03784_);
  and (_03880_, _03879_, _03474_);
  and (_03881_, _03784_, _03488_);
  and (_03882_, _03881_, _03492_);
  or (_03883_, _03882_, _03880_);
  and (_03884_, _03784_, _03540_);
  and (_03885_, _03884_, _03742_);
  and (_03886_, _03835_, _03784_);
  and (_03887_, _03886_, _03596_);
  or (_03888_, _03887_, _03885_);
  or (_03889_, _03888_, _03883_);
  or (_03890_, _03889_, _03878_);
  and (_03891_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03892_, _03786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03893_, _03892_, _03891_);
  or (_03894_, _03893_, _03890_);
  or (_03895_, _03894_, _03866_);
  and (_03896_, _03895_, _03802_);
  not (_03897_, _03802_);
  nand (_03898_, _03334_, _03342_);
  nor (_03899_, _03821_, _03818_);
  and (_03900_, _03899_, _03898_);
  nor (_03901_, _03828_, _03826_);
  nor (_03902_, _03836_, _03831_);
  and (_03903_, _03902_, _03901_);
  and (_03904_, _03903_, _03900_);
  nor (_03905_, _03844_, _03841_);
  nor (_03906_, _03849_, _03847_);
  and (_03907_, _03906_, _03905_);
  nor (_03908_, _03856_, _03854_);
  nor (_03909_, _03861_, _03859_);
  and (_03910_, _03909_, _03908_);
  and (_03911_, _03910_, _03907_);
  and (_03912_, _03911_, _03904_);
  nand (_03913_, _03784_, _03535_);
  nor (_03914_, _03875_, _03804_);
  and (_03915_, _03783_, _03353_);
  and (_03916_, _03915_, _03488_);
  nor (_03917_, _03916_, _03870_);
  and (_03918_, _03917_, _03914_);
  and (_03919_, _03918_, _03913_);
  nor (_03920_, _03794_, _03786_);
  and (_03921_, _03920_, _03919_);
  and (_03922_, _03921_, _03912_);
  nor (_03923_, _03922_, _03897_);
  nor (_03924_, _03923_, _20647_);
  or (_03925_, _03924_, _03896_);
  or (_03926_, _03925_, _03805_);
  and (_03927_, _03926_, _42355_);
  and (_39423_, _03927_, _03807_);
  nor (_39502_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_03928_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_03930_, _03320_, rst);
  and (_39503_, _03930_, _03928_);
  nor (_03931_, _03320_, _03319_);
  or (_03932_, _03931_, _03321_);
  and (_03933_, _03324_, _42355_);
  and (_39504_, _03933_, _03932_);
  nand (_03934_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_03935_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_03936_, _03935_, _03934_);
  nand (_03937_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_03938_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_03939_, _03938_, _03937_);
  and (_03940_, _03939_, _03936_);
  nand (_03941_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_03942_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_03943_, _03942_, _03941_);
  nand (_03944_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_03945_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_03946_, _03945_, _03944_);
  and (_03947_, _03946_, _03943_);
  and (_03948_, _03947_, _03940_);
  nand (_03949_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_03950_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_03951_, _03950_, _03949_);
  nand (_03952_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_03953_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_03954_, _03953_, _03952_);
  and (_03955_, _03954_, _03951_);
  nand (_03956_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_03957_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_03958_, _03957_, _03956_);
  nand (_03959_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_03960_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_03961_, _03960_, _03959_);
  and (_03962_, _03961_, _03958_);
  and (_03963_, _03962_, _03955_);
  and (_03964_, _03963_, _03948_);
  nand (_03965_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_03966_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_03967_, _03966_, _03965_);
  nand (_03968_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_03969_, _03868_, _42015_);
  and (_03970_, _03969_, _03968_);
  and (_03971_, _03970_, _03967_);
  nand (_03972_, _03884_, _03727_);
  nand (_03973_, _03886_, _03606_);
  and (_03974_, _03973_, _03972_);
  nand (_03975_, _03879_, _03449_);
  nand (_03976_, _03881_, _03502_);
  and (_03977_, _03976_, _03975_);
  and (_03978_, _03977_, _03974_);
  and (_03979_, _03978_, _03971_);
  not (_03980_, _03786_);
  or (_03981_, _03980_, _03572_);
  nand (_03982_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_03983_, _03982_, _03981_);
  and (_03984_, _03983_, _03979_);
  and (_03985_, _03984_, _03964_);
  nor (_03986_, _03985_, _03897_);
  not (_03987_, _03805_);
  or (_03988_, _03923_, _19488_);
  nand (_03989_, _03988_, _03987_);
  or (_03990_, _03989_, _03986_);
  nand (_03991_, _03805_, _32444_);
  and (_03992_, _03991_, _42355_);
  and (_39506_, _03992_, _03990_);
  nand (_03993_, _03805_, _33119_);
  and (_03994_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_03995_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_03996_, _03995_, _03994_);
  and (_03997_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_03998_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_03999_, _03998_, _03997_);
  or (_04000_, _03999_, _03996_);
  and (_04001_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_04002_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_04003_, _04002_, _04001_);
  and (_04004_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04005_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_04006_, _04005_, _04004_);
  or (_04007_, _04006_, _04003_);
  or (_04008_, _04007_, _04000_);
  and (_04009_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_04010_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_04011_, _04010_, _04009_);
  and (_04012_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_04013_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_04014_, _04013_, _04012_);
  or (_04015_, _04014_, _04011_);
  and (_04016_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_04017_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_04018_, _04017_, _04016_);
  and (_04019_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_04020_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_04021_, _04020_, _04019_);
  or (_04022_, _04021_, _04018_);
  or (_04023_, _04022_, _04015_);
  or (_04024_, _04023_, _04008_);
  and (_04025_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_04026_, _03868_, _41917_);
  or (_04028_, _04026_, _04025_);
  and (_04029_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_04030_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_04031_, _04030_, _04029_);
  or (_04032_, _04031_, _04028_);
  and (_04033_, _03881_, _03522_);
  and (_04034_, _03879_, _03445_);
  or (_04035_, _04034_, _04033_);
  and (_04036_, _03884_, _03707_);
  and (_04037_, _03886_, _03627_);
  or (_04038_, _04037_, _04036_);
  or (_04039_, _04038_, _04035_);
  or (_04040_, _04039_, _04032_);
  and (_04041_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_04042_, _03786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_04043_, _04042_, _04041_);
  or (_04044_, _04043_, _04040_);
  or (_04045_, _04044_, _04024_);
  or (_04046_, _03802_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_04047_, _04046_, _04045_);
  nor (_04048_, _03923_, _20473_);
  or (_04049_, _04048_, _03805_);
  or (_04050_, _04049_, _04047_);
  and (_04051_, _04050_, _42355_);
  and (_39507_, _04051_, _03993_);
  and (_04052_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04053_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_04054_, _04053_, _04052_);
  and (_04055_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_04056_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_04057_, _04056_, _04055_);
  or (_04058_, _04057_, _04054_);
  and (_04059_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_04060_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_04061_, _04060_, _04059_);
  and (_04062_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_04063_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_04064_, _04063_, _04062_);
  or (_04065_, _04064_, _04061_);
  or (_04066_, _04065_, _04058_);
  and (_04067_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_04068_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_04069_, _04068_, _04067_);
  and (_04070_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_04071_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_04072_, _04071_, _04070_);
  or (_04073_, _04072_, _04069_);
  and (_04074_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_04075_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_04076_, _04075_, _04074_);
  and (_04077_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_04078_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_04079_, _04078_, _04077_);
  or (_04080_, _04079_, _04076_);
  or (_04081_, _04080_, _04073_);
  or (_04082_, _04081_, _04066_);
  and (_04083_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_04084_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_04085_, _04084_, _04083_);
  and (_04086_, _03868_, _42158_);
  and (_04087_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_04088_, _04087_, _04086_);
  or (_04089_, _04088_, _04085_);
  and (_04090_, _03879_, _03458_);
  and (_04091_, _03881_, _03516_);
  or (_04092_, _04091_, _04090_);
  and (_04093_, _03884_, _03717_);
  and (_04094_, _03886_, _03621_);
  or (_04095_, _04094_, _04093_);
  or (_04096_, _04095_, _04092_);
  or (_04097_, _04096_, _04089_);
  and (_04098_, _03786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_04099_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_04100_, _04099_, _04098_);
  or (_04101_, _04100_, _04097_);
  or (_04102_, _04101_, _04082_);
  or (_04103_, _03802_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_04104_, _04103_, _04102_);
  nor (_04105_, _03923_, _19126_);
  or (_04106_, _04105_, _03805_);
  or (_04107_, _04106_, _04104_);
  nand (_04108_, _03805_, _33837_);
  and (_04109_, _04108_, _42355_);
  and (_39508_, _04109_, _04107_);
  and (_04110_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_04111_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_04112_, _04111_, _04110_);
  and (_04113_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_04114_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_04115_, _04114_, _04113_);
  or (_04116_, _04115_, _04112_);
  and (_04117_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_04118_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_04119_, _04118_, _04117_);
  and (_04120_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_04121_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_04122_, _04121_, _04120_);
  or (_04123_, _04122_, _04119_);
  or (_04124_, _04123_, _04116_);
  and (_04125_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_04127_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_04128_, _04127_, _04125_);
  and (_04129_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_04130_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_04131_, _04130_, _04129_);
  or (_04132_, _04131_, _04128_);
  and (_04133_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_04134_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_04135_, _04134_, _04133_);
  and (_04136_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_04137_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_04138_, _04137_, _04136_);
  or (_04139_, _04138_, _04135_);
  or (_04140_, _04139_, _04132_);
  or (_04141_, _04140_, _04124_);
  and (_04142_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_04143_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_04144_, _04143_, _04142_);
  and (_04145_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_04146_, _03868_, _41972_);
  or (_04147_, _04146_, _04145_);
  or (_04148_, _04147_, _04144_);
  and (_04149_, _03879_, _03454_);
  and (_04150_, _03881_, _03496_);
  or (_04151_, _04150_, _04149_);
  and (_04152_, _03884_, _03738_);
  and (_04153_, _03886_, _03600_);
  or (_04154_, _04153_, _04152_);
  or (_04155_, _04154_, _04151_);
  or (_04156_, _04155_, _04148_);
  and (_04157_, _03786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_04158_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_04159_, _04158_, _04157_);
  or (_04160_, _04159_, _04156_);
  or (_04161_, _04160_, _04141_);
  or (_04162_, _03802_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_04163_, _04162_, _04161_);
  nor (_04164_, _03923_, _20158_);
  or (_04165_, _04164_, _03805_);
  or (_04166_, _04165_, _04163_);
  or (_04167_, _03987_, _34566_);
  and (_04168_, _04167_, _42355_);
  and (_39509_, _04168_, _04166_);
  or (_04169_, _03987_, _35229_);
  and (_04170_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_04171_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_04172_, _04171_, _04170_);
  and (_04173_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_04174_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_04175_, _04174_, _04173_);
  or (_04176_, _04175_, _04172_);
  and (_04177_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_04178_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_04179_, _04178_, _04177_);
  and (_04180_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_04181_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_04182_, _04181_, _04180_);
  or (_04183_, _04182_, _04179_);
  or (_04184_, _04183_, _04176_);
  and (_04185_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_04186_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_04187_, _04186_, _04185_);
  and (_04188_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_04189_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_04190_, _04189_, _04188_);
  or (_04191_, _04190_, _04187_);
  and (_04192_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_04193_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_04194_, _04193_, _04192_);
  and (_04195_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_04196_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_04197_, _04196_, _04195_);
  or (_04198_, _04197_, _04194_);
  or (_04199_, _04198_, _04191_);
  or (_04200_, _04199_, _04184_);
  and (_04201_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_04202_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_04203_, _04202_, _04201_);
  and (_04204_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_04205_, _03868_, _41889_);
  or (_04206_, _04205_, _04204_);
  or (_04207_, _04206_, _04203_);
  and (_04208_, _03881_, _03506_);
  and (_04209_, _03879_, _03469_);
  or (_04210_, _04209_, _04208_);
  and (_04211_, _03884_, _03731_);
  and (_04212_, _03886_, _03610_);
  or (_04213_, _04212_, _04211_);
  or (_04214_, _04213_, _04210_);
  or (_04215_, _04214_, _04207_);
  and (_04216_, _03786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_04217_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_04218_, _04217_, _04216_);
  or (_04219_, _04218_, _04215_);
  or (_04220_, _04219_, _04200_);
  or (_04221_, _03802_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_04222_, _04221_, _04220_);
  nor (_04223_, _03923_, _19324_);
  or (_04224_, _04223_, _03805_);
  or (_04225_, _04224_, _04222_);
  and (_04227_, _04225_, _42355_);
  and (_39510_, _04227_, _04169_);
  and (_04228_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04229_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_04230_, _04229_, _04228_);
  and (_04231_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_04232_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04233_, _04232_, _04231_);
  or (_04234_, _04233_, _04230_);
  and (_04235_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04236_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_04237_, _04236_, _04235_);
  and (_04238_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04239_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_04240_, _04239_, _04238_);
  or (_04241_, _04240_, _04237_);
  or (_04242_, _04241_, _04234_);
  and (_04243_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_04244_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_04245_, _04244_, _04243_);
  and (_04246_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_04247_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_04248_, _04247_, _04246_);
  or (_04249_, _04248_, _04245_);
  and (_04250_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_04251_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_04252_, _04251_, _04250_);
  and (_04253_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_04254_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_04255_, _04254_, _04253_);
  or (_04256_, _04255_, _04252_);
  or (_04257_, _04256_, _04249_);
  or (_04258_, _04257_, _04242_);
  and (_04259_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_04260_, _38003_);
  and (_04261_, _03868_, _04260_);
  or (_04262_, _04261_, _04259_);
  and (_04263_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_04264_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_04265_, _04264_, _04263_);
  or (_04266_, _04265_, _04262_);
  and (_04267_, _03881_, _03526_);
  and (_04268_, _03879_, _03465_);
  or (_04269_, _04268_, _04267_);
  and (_04270_, _03884_, _03711_);
  and (_04271_, _03886_, _03631_);
  or (_04272_, _04271_, _04270_);
  or (_04273_, _04272_, _04269_);
  or (_04274_, _04273_, _04266_);
  and (_04275_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_04276_, _03786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_04277_, _04276_, _04275_);
  or (_04278_, _04277_, _04274_);
  or (_04279_, _04278_, _04258_);
  or (_04280_, _03802_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_04281_, _04280_, _04279_);
  nor (_04282_, _03923_, _20310_);
  or (_04283_, _04282_, _03805_);
  or (_04284_, _04283_, _04281_);
  nand (_04285_, _03805_, _36025_);
  and (_04286_, _04285_, _42355_);
  and (_39511_, _04286_, _04284_);
  nand (_04287_, _03805_, _36752_);
  and (_04288_, _03810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_04289_, _03814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_04290_, _04289_, _04288_);
  and (_04291_, _03818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_04292_, _03821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_04293_, _04292_, _04291_);
  or (_04294_, _04293_, _04290_);
  and (_04295_, _03826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_04296_, _03828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_04297_, _04296_, _04295_);
  and (_04298_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04299_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_04300_, _04299_, _04298_);
  or (_04301_, _04300_, _04297_);
  or (_04302_, _04301_, _04294_);
  and (_04303_, _03841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_04304_, _03844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or (_04305_, _04304_, _04303_);
  and (_04306_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_04307_, _03849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_04308_, _04307_, _04306_);
  or (_04309_, _04308_, _04305_);
  and (_04310_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_04311_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04312_, _04311_, _04310_);
  and (_04313_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_04314_, _03859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_04315_, _04314_, _04313_);
  or (_04316_, _04315_, _04312_);
  or (_04317_, _04316_, _04309_);
  or (_04318_, _04317_, _04302_);
  and (_04319_, _03868_, _42069_);
  and (_04320_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_04321_, _04320_, _04319_);
  and (_04322_, _03804_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_04323_, _03875_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_04324_, _04323_, _04322_);
  or (_04326_, _04324_, _04321_);
  and (_04327_, _03879_, _03478_);
  and (_04328_, _03881_, _03512_);
  or (_04329_, _04328_, _04327_);
  and (_04330_, _03884_, _03721_);
  and (_04331_, _03886_, _03617_);
  or (_04332_, _04331_, _04330_);
  or (_04333_, _04332_, _04329_);
  or (_04334_, _04333_, _04326_);
  and (_04335_, _03794_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_04336_, _03786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_04337_, _04336_, _04335_);
  or (_04338_, _04337_, _04334_);
  or (_04339_, _04338_, _04318_);
  or (_04340_, _03802_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_04341_, _04340_, _04339_);
  nor (_04342_, _03923_, _19661_);
  or (_04343_, _04342_, _03805_);
  or (_04344_, _04343_, _04341_);
  and (_04345_, _04344_, _42355_);
  and (_39512_, _04345_, _04287_);
  and (_39582_, _42217_, _42355_);
  nor (_39585_, _42180_, rst);
  and (_39606_, _42370_, _42355_);
  nor (_39609_, _42037_, rst);
  nor (_39610_, _41939_, rst);
  not (_04346_, _00401_);
  nor (_04347_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_04348_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04349_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04348_);
  nor (_04350_, _04349_, _04347_);
  nor (_04351_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04352_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04348_);
  nor (_04353_, _04352_, _04351_);
  not (_04354_, _04353_);
  nor (_04355_, _04354_, _04350_);
  and (_04356_, _04353_, _04350_);
  nor (_04357_, _02214_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04358_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04348_);
  nor (_04359_, _04358_, _04357_);
  and (_04360_, _04359_, _04356_);
  nor (_04361_, _04359_, _04356_);
  nor (_04362_, _04361_, _04360_);
  not (_04363_, _04362_);
  nor (_04364_, _02234_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04365_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04348_);
  nor (_04366_, _04365_, _04364_);
  and (_04367_, _04366_, _04360_);
  nor (_04368_, _04366_, _04360_);
  nor (_04369_, _04368_, _04367_);
  and (_04370_, _04369_, _04363_);
  and (_04371_, _04370_, _04355_);
  and (_04372_, _04371_, _04346_);
  not (_04373_, _00319_);
  nor (_04374_, _04353_, _04350_);
  and (_04375_, _04374_, _04370_);
  and (_04376_, _04375_, _04373_);
  or (_04377_, _04376_, _04372_);
  not (_04378_, _00360_);
  and (_04379_, _04354_, _04350_);
  and (_04380_, _04379_, _04370_);
  and (_04381_, _04380_, _04378_);
  not (_04382_, _00042_);
  nor (_04383_, _04369_, _04362_);
  and (_04384_, _04383_, _04355_);
  and (_04385_, _04384_, _04382_);
  or (_04386_, _04385_, _04381_);
  or (_04387_, _04386_, _04377_);
  not (_04388_, _43226_);
  and (_04389_, _04383_, _04374_);
  and (_04390_, _04389_, _04388_);
  not (_04391_, _43267_);
  and (_04392_, _04383_, _04379_);
  and (_04393_, _04392_, _04391_);
  or (_04394_, _04393_, _04390_);
  not (_04395_, _00196_);
  not (_04396_, _04366_);
  and (_04397_, _04396_, _04362_);
  and (_04398_, _04397_, _04379_);
  and (_04399_, _04398_, _04395_);
  not (_04400_, _00124_);
  and (_04401_, _04397_, _04374_);
  and (_04402_, _04401_, _04400_);
  or (_04403_, _04402_, _04399_);
  not (_04404_, _00483_);
  and (_04405_, _04366_, _04362_);
  and (_04406_, _04405_, _04374_);
  and (_04407_, _04406_, _04404_);
  not (_04408_, _00237_);
  and (_04409_, _04397_, _04355_);
  and (_04410_, _04409_, _04408_);
  or (_04411_, _04410_, _04407_);
  or (_04412_, _04411_, _04403_);
  not (_04413_, _00083_);
  and (_04414_, _04368_, _04356_);
  and (_04415_, _04414_, _04413_);
  not (_04416_, _43185_);
  and (_04417_, _04367_, _04416_);
  not (_04418_, _00579_);
  and (_04420_, _04359_, _04355_);
  and (_04421_, _04420_, _04366_);
  and (_04422_, _04421_, _04418_);
  not (_04423_, _00278_);
  and (_04424_, _04396_, _04360_);
  and (_04425_, _04424_, _04423_);
  or (_04426_, _04425_, _04422_);
  or (_04427_, _04426_, _04417_);
  or (_04428_, _04427_, _04415_);
  not (_04429_, _00524_);
  and (_04430_, _04405_, _04379_);
  and (_04431_, _04430_, _04429_);
  not (_04432_, _00442_);
  and (_04433_, _04405_, _04356_);
  and (_04434_, _04433_, _04432_);
  or (_04435_, _04434_, _04431_);
  or (_04436_, _04435_, _04428_);
  or (_04437_, _04436_, _04412_);
  or (_04438_, _04437_, _04394_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04438_, _04387_);
  and (_04439_, _04371_, _04432_);
  and (_04440_, _04384_, _04413_);
  or (_04441_, _04440_, _04439_);
  and (_04442_, _04380_, _04346_);
  and (_04443_, _04375_, _04378_);
  or (_04444_, _04443_, _04442_);
  or (_04445_, _04444_, _04441_);
  and (_04446_, _04406_, _04429_);
  and (_04447_, _04409_, _04423_);
  or (_04448_, _04447_, _04446_);
  and (_04449_, _04430_, _04418_);
  and (_04450_, _04401_, _04395_);
  or (_04451_, _04450_, _04449_);
  or (_04452_, _04451_, _04448_);
  and (_04453_, _04414_, _04400_);
  and (_04454_, _04424_, _04373_);
  and (_04455_, _04421_, _04416_);
  and (_04456_, _04367_, _04388_);
  or (_04457_, _04456_, _04455_);
  or (_04458_, _04457_, _04454_);
  or (_04459_, _04458_, _04453_);
  and (_04460_, _04433_, _04404_);
  and (_04461_, _04398_, _04408_);
  or (_04462_, _04461_, _04460_);
  or (_04463_, _04462_, _04459_);
  or (_04464_, _04463_, _04452_);
  and (_04465_, _04392_, _04382_);
  and (_04466_, _04389_, _04391_);
  or (_04467_, _04466_, _04465_);
  or (_04468_, _04467_, _04464_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04468_, _04445_);
  and (_04469_, _04371_, _04404_);
  and (_04470_, _04375_, _04346_);
  or (_04471_, _04470_, _04469_);
  and (_04472_, _04380_, _04432_);
  and (_04473_, _04384_, _04400_);
  or (_04474_, _04473_, _04472_);
  or (_04475_, _04474_, _04471_);
  and (_04476_, _04392_, _04413_);
  and (_04477_, _04389_, _04382_);
  or (_04478_, _04477_, _04476_);
  and (_04479_, _04409_, _04373_);
  and (_04480_, _04398_, _04423_);
  or (_04481_, _04480_, _04479_);
  and (_04482_, _04401_, _04408_);
  and (_04483_, _04430_, _04416_);
  or (_04484_, _04483_, _04482_);
  or (_04485_, _04484_, _04481_);
  and (_04486_, _04414_, _04395_);
  and (_04487_, _04367_, _04391_);
  and (_04488_, _04424_, _04378_);
  and (_04489_, _04421_, _04388_);
  or (_04490_, _04489_, _04488_);
  or (_04491_, _04490_, _04487_);
  or (_04492_, _04491_, _04486_);
  and (_04493_, _04406_, _04418_);
  and (_04494_, _04433_, _04429_);
  or (_04495_, _04494_, _04493_);
  or (_04496_, _04495_, _04492_);
  or (_04497_, _04496_, _04485_);
  or (_04498_, _04497_, _04478_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04498_, _04475_);
  and (_04499_, _04380_, _04373_);
  and (_04500_, _04371_, _04378_);
  or (_04501_, _04500_, _04499_);
  and (_04502_, _04375_, _04423_);
  and (_04503_, _04384_, _04391_);
  or (_04504_, _04503_, _04502_);
  or (_04505_, _04504_, _04501_);
  and (_04506_, _04409_, _04395_);
  and (_04507_, _04401_, _04413_);
  or (_04508_, _04507_, _04506_);
  and (_04509_, _04433_, _04346_);
  and (_04510_, _04398_, _04400_);
  or (_04511_, _04510_, _04509_);
  or (_04512_, _04511_, _04508_);
  and (_04513_, _04414_, _04382_);
  and (_04514_, _04424_, _04408_);
  and (_04515_, _04367_, _04418_);
  and (_04516_, _04421_, _04429_);
  or (_04518_, _04516_, _04515_);
  or (_04519_, _04518_, _04514_);
  or (_04520_, _04519_, _04513_);
  and (_04521_, _04430_, _04404_);
  and (_04522_, _04406_, _04432_);
  or (_04523_, _04522_, _04521_);
  or (_04524_, _04523_, _04520_);
  or (_04525_, _04524_, _04512_);
  and (_04526_, _04389_, _04416_);
  and (_04527_, _04392_, _04388_);
  or (_04528_, _04527_, _04526_);
  or (_04529_, _04528_, _04525_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04529_, _04505_);
  not (_04530_, _00324_);
  and (_04531_, _04380_, _04530_);
  not (_04532_, _00365_);
  and (_04533_, _04371_, _04532_);
  or (_04534_, _04533_, _04531_);
  not (_04535_, _00283_);
  and (_04536_, _04375_, _04535_);
  not (_04537_, _00006_);
  and (_04538_, _04384_, _04537_);
  or (_04539_, _04538_, _04536_);
  or (_04540_, _04539_, _04534_);
  not (_04541_, _00488_);
  and (_04542_, _04430_, _04541_);
  not (_04543_, _00129_);
  and (_04544_, _04398_, _04543_);
  or (_04545_, _04544_, _04542_);
  not (_04546_, _00406_);
  and (_04547_, _04433_, _04546_);
  not (_04548_, _00201_);
  and (_04549_, _04409_, _04548_);
  or (_04550_, _04549_, _04547_);
  or (_04551_, _04550_, _04545_);
  not (_04552_, _00047_);
  and (_04553_, _04414_, _04552_);
  not (_04554_, _00587_);
  and (_04555_, _04367_, _04554_);
  not (_04556_, _00529_);
  and (_04557_, _04421_, _04556_);
  not (_04558_, _00242_);
  and (_04559_, _04424_, _04558_);
  or (_04560_, _04559_, _04557_);
  or (_04561_, _04560_, _04555_);
  or (_04562_, _04561_, _04553_);
  not (_04563_, _00447_);
  and (_04564_, _04406_, _04563_);
  not (_04565_, _00088_);
  and (_04566_, _04401_, _04565_);
  or (_04567_, _04566_, _04564_);
  or (_04568_, _04567_, _04562_);
  or (_04569_, _04568_, _04551_);
  not (_04570_, _43190_);
  and (_04571_, _04389_, _04570_);
  not (_04572_, _43231_);
  and (_04573_, _04392_, _04572_);
  or (_04574_, _04573_, _04571_);
  or (_04575_, _04574_, _04569_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _04575_, _04540_);
  not (_04576_, _00329_);
  and (_04577_, _04380_, _04576_);
  not (_04578_, _00370_);
  and (_04579_, _04371_, _04578_);
  or (_04580_, _04579_, _04577_);
  not (_04581_, _00288_);
  and (_04582_, _04375_, _04581_);
  not (_04583_, _00011_);
  and (_04584_, _04384_, _04583_);
  or (_04585_, _04584_, _04582_);
  or (_04586_, _04585_, _04580_);
  not (_04587_, _00206_);
  and (_04588_, _04409_, _04587_);
  not (_04589_, _00093_);
  and (_04590_, _04401_, _04589_);
  or (_04591_, _04590_, _04588_);
  not (_04592_, _00411_);
  and (_04593_, _04433_, _04592_);
  not (_04594_, _00139_);
  and (_04595_, _04398_, _04594_);
  or (_04596_, _04595_, _04593_);
  or (_04597_, _04596_, _04591_);
  not (_04598_, _00052_);
  and (_04599_, _04414_, _04598_);
  not (_04600_, _00594_);
  and (_04601_, _04367_, _04600_);
  not (_04602_, _00534_);
  and (_04603_, _04421_, _04602_);
  not (_04604_, _00247_);
  and (_04605_, _04424_, _04604_);
  or (_04606_, _04605_, _04603_);
  or (_04607_, _04606_, _04601_);
  or (_04608_, _04607_, _04599_);
  not (_04609_, _00493_);
  and (_04610_, _04430_, _04609_);
  not (_04611_, _00452_);
  and (_04612_, _04406_, _04611_);
  or (_04613_, _04612_, _04610_);
  or (_04614_, _04613_, _04608_);
  or (_04615_, _04614_, _04597_);
  not (_04617_, _43195_);
  and (_04618_, _04389_, _04617_);
  not (_04619_, _43236_);
  and (_04620_, _04392_, _04619_);
  or (_04621_, _04620_, _04618_);
  or (_04622_, _04621_, _04615_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _04622_, _04586_);
  not (_04623_, _00599_);
  and (_04624_, _04367_, _04623_);
  not (_04625_, _00016_);
  and (_04626_, _04384_, _04625_);
  not (_04627_, _43200_);
  and (_04628_, _04389_, _04627_);
  or (_04629_, _04628_, _04626_);
  not (_04630_, _43241_);
  and (_04631_, _04392_, _04630_);
  not (_04632_, _00211_);
  and (_04633_, _04409_, _04632_);
  not (_04634_, _00150_);
  and (_04635_, _04398_, _04634_);
  or (_04636_, _04635_, _04633_);
  not (_04637_, _00098_);
  and (_04638_, _04401_, _04637_);
  not (_04639_, _00057_);
  and (_04640_, _04414_, _04639_);
  or (_04641_, _04640_, _04638_);
  or (_04642_, _04641_, _04636_);
  or (_04643_, _04642_, _04631_);
  or (_04644_, _04643_, _04629_);
  not (_04645_, _00498_);
  and (_04646_, _04430_, _04645_);
  not (_04647_, _00539_);
  and (_04648_, _04421_, _04647_);
  or (_04649_, _04648_, _04646_);
  not (_04650_, _00416_);
  and (_04651_, _04433_, _04650_);
  not (_04652_, _00457_);
  and (_04653_, _04406_, _04652_);
  or (_04654_, _04653_, _04651_);
  or (_04655_, _04654_, _04649_);
  not (_04656_, _00375_);
  and (_04657_, _04371_, _04656_);
  not (_04658_, _00334_);
  and (_04659_, _04380_, _04658_);
  or (_04660_, _04659_, _04657_);
  not (_04661_, _00293_);
  and (_04662_, _04375_, _04661_);
  not (_04663_, _00252_);
  and (_04664_, _04424_, _04663_);
  or (_04665_, _04664_, _04662_);
  or (_04666_, _04665_, _04660_);
  or (_04667_, _04666_, _04655_);
  or (_04668_, _04667_, _04644_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _04668_, _04624_);
  not (_04669_, _00339_);
  and (_04670_, _04380_, _04669_);
  not (_04671_, _00380_);
  and (_04672_, _04371_, _04671_);
  or (_04673_, _04672_, _04670_);
  not (_04674_, _00298_);
  and (_04675_, _04375_, _04674_);
  not (_04676_, _00021_);
  and (_04677_, _04384_, _04676_);
  or (_04678_, _04677_, _04675_);
  or (_04679_, _04678_, _04673_);
  not (_04680_, _43205_);
  and (_04681_, _04389_, _04680_);
  not (_04682_, _43246_);
  and (_04683_, _04392_, _04682_);
  or (_04684_, _04683_, _04681_);
  not (_04685_, _00462_);
  and (_04686_, _04406_, _04685_);
  not (_04687_, _00421_);
  and (_04688_, _04433_, _04687_);
  or (_04689_, _04688_, _04686_);
  not (_04690_, _00216_);
  and (_04691_, _04409_, _04690_);
  not (_04692_, _00103_);
  and (_04693_, _04401_, _04692_);
  or (_04694_, _04693_, _04691_);
  or (_04695_, _04694_, _04689_);
  not (_04696_, _00062_);
  and (_04697_, _04414_, _04696_);
  not (_04698_, _00604_);
  and (_04699_, _04367_, _04698_);
  not (_04700_, _00545_);
  and (_04701_, _04421_, _04700_);
  not (_04702_, _00257_);
  and (_04703_, _04424_, _04702_);
  or (_04704_, _04703_, _04701_);
  or (_04705_, _04704_, _04699_);
  or (_04706_, _04705_, _04697_);
  not (_04707_, _00503_);
  and (_04708_, _04430_, _04707_);
  not (_04709_, _00161_);
  and (_04710_, _04398_, _04709_);
  or (_04711_, _04710_, _04708_);
  or (_04712_, _04711_, _04706_);
  or (_04713_, _04712_, _04695_);
  or (_04714_, _04713_, _04684_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _04714_, _04679_);
  not (_04715_, _00609_);
  and (_04716_, _04367_, _04715_);
  not (_04717_, _00026_);
  and (_04718_, _04384_, _04717_);
  not (_04719_, _43210_);
  and (_04720_, _04389_, _04719_);
  or (_04721_, _04720_, _04718_);
  not (_04722_, _43251_);
  and (_04723_, _04392_, _04722_);
  not (_04724_, _00221_);
  and (_04725_, _04409_, _04724_);
  not (_04726_, _00172_);
  and (_04727_, _04398_, _04726_);
  or (_04728_, _04727_, _04725_);
  not (_04729_, _00108_);
  and (_04730_, _04401_, _04729_);
  not (_04731_, _00067_);
  and (_04732_, _04414_, _04731_);
  or (_04733_, _04732_, _04730_);
  or (_04734_, _04733_, _04728_);
  or (_04735_, _04734_, _04723_);
  or (_04736_, _04735_, _04721_);
  not (_04737_, _00508_);
  and (_04738_, _04430_, _04737_);
  not (_04739_, _00553_);
  and (_04740_, _04421_, _04739_);
  or (_04741_, _04740_, _04738_);
  not (_04742_, _00426_);
  and (_04743_, _04433_, _04742_);
  not (_04744_, _00467_);
  and (_04745_, _04406_, _04744_);
  or (_04746_, _04745_, _04743_);
  or (_04747_, _04746_, _04741_);
  not (_04748_, _00385_);
  and (_04749_, _04371_, _04748_);
  not (_04750_, _00344_);
  and (_04751_, _04380_, _04750_);
  or (_04752_, _04751_, _04749_);
  not (_04753_, _00303_);
  and (_04754_, _04375_, _04753_);
  not (_04755_, _00262_);
  and (_04756_, _04424_, _04755_);
  or (_04757_, _04756_, _04754_);
  or (_04758_, _04757_, _04752_);
  or (_04759_, _04758_, _04747_);
  or (_04760_, _04759_, _04736_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _04760_, _04716_);
  not (_04761_, _00349_);
  and (_04762_, _04380_, _04761_);
  not (_04763_, _00390_);
  and (_04764_, _04371_, _04763_);
  or (_04765_, _04764_, _04762_);
  not (_04766_, _00308_);
  and (_04767_, _04375_, _04766_);
  not (_04768_, _00031_);
  and (_04769_, _04384_, _04768_);
  or (_04770_, _04769_, _04767_);
  or (_04771_, _04770_, _04765_);
  not (_04772_, _00513_);
  and (_04773_, _04430_, _04772_);
  not (_04774_, _00183_);
  and (_04775_, _04398_, _04774_);
  or (_04776_, _04775_, _04773_);
  not (_04777_, _00431_);
  and (_04778_, _04433_, _04777_);
  not (_04779_, _00226_);
  and (_04780_, _04409_, _04779_);
  or (_04781_, _04780_, _04778_);
  or (_04782_, _04781_, _04776_);
  not (_04783_, _00072_);
  and (_04784_, _04414_, _04783_);
  not (_04785_, _00267_);
  and (_04786_, _04424_, _04785_);
  not (_04787_, _00614_);
  and (_04788_, _04367_, _04787_);
  not (_04789_, _00561_);
  and (_04790_, _04421_, _04789_);
  or (_04791_, _04790_, _04788_);
  or (_04792_, _04791_, _04786_);
  or (_04793_, _04792_, _04784_);
  not (_04794_, _00472_);
  and (_04795_, _04406_, _04794_);
  not (_04796_, _00113_);
  and (_04797_, _04401_, _04796_);
  or (_04798_, _04797_, _04795_);
  or (_04799_, _04798_, _04793_);
  or (_04800_, _04799_, _04782_);
  not (_04801_, _43215_);
  and (_04802_, _04389_, _04801_);
  not (_04803_, _43256_);
  and (_04804_, _04392_, _04803_);
  or (_04805_, _04804_, _04802_);
  or (_04806_, _04805_, _04800_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _04806_, _04771_);
  not (_04807_, _00036_);
  and (_04808_, _04384_, _04807_);
  not (_04809_, _00395_);
  and (_04810_, _04371_, _04809_);
  or (_04811_, _04810_, _04808_);
  not (_04812_, _00354_);
  and (_04813_, _04380_, _04812_);
  not (_04814_, _00313_);
  and (_04815_, _04375_, _04814_);
  or (_04816_, _04815_, _04813_);
  or (_04817_, _04816_, _04811_);
  not (_04818_, _00118_);
  and (_04819_, _04401_, _04818_);
  not (_04820_, _00518_);
  and (_04821_, _04430_, _04820_);
  or (_04822_, _04821_, _04819_);
  not (_04823_, _00231_);
  and (_04824_, _04409_, _04823_);
  not (_04825_, _00436_);
  and (_04826_, _04433_, _04825_);
  or (_04827_, _04826_, _04824_);
  or (_04828_, _04827_, _04822_);
  not (_04829_, _00077_);
  and (_04830_, _04414_, _04829_);
  not (_04831_, _00272_);
  and (_04832_, _04424_, _04831_);
  not (_04833_, _00619_);
  and (_04834_, _04367_, _04833_);
  not (_04835_, _00569_);
  and (_04836_, _04421_, _04835_);
  or (_04837_, _04836_, _04834_);
  or (_04838_, _04837_, _04832_);
  or (_04839_, _04838_, _04830_);
  not (_04840_, _00190_);
  and (_04841_, _04398_, _04840_);
  not (_04842_, _00477_);
  and (_04843_, _04406_, _04842_);
  or (_04844_, _04843_, _04841_);
  or (_04845_, _04844_, _04839_);
  or (_04846_, _04845_, _04828_);
  not (_04847_, _43220_);
  and (_04848_, _04389_, _04847_);
  not (_04849_, _43261_);
  and (_04850_, _04392_, _04849_);
  or (_04851_, _04850_, _04848_);
  or (_04852_, _04851_, _04846_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _04852_, _04817_);
  and (_04853_, _04375_, _04546_);
  and (_04854_, _04384_, _04543_);
  or (_04855_, _04854_, _04853_);
  and (_04856_, _04380_, _04563_);
  and (_04857_, _04371_, _04541_);
  or (_04858_, _04857_, _04856_);
  or (_04859_, _04858_, _04855_);
  and (_04860_, _04389_, _04552_);
  and (_04861_, _04392_, _04565_);
  or (_04862_, _04861_, _04860_);
  and (_04863_, _04406_, _04554_);
  and (_04864_, _04409_, _04530_);
  or (_04865_, _04864_, _04863_);
  and (_04866_, _04433_, _04556_);
  and (_04867_, _04401_, _04558_);
  or (_04868_, _04867_, _04866_);
  or (_04869_, _04868_, _04865_);
  and (_04870_, _04414_, _04548_);
  and (_04871_, _04421_, _04572_);
  and (_04872_, _04424_, _04532_);
  and (_04873_, _04367_, _04537_);
  or (_04874_, _04873_, _04872_);
  or (_04875_, _04874_, _04871_);
  or (_04876_, _04875_, _04870_);
  and (_04877_, _04398_, _04535_);
  and (_04878_, _04430_, _04570_);
  or (_04879_, _04878_, _04877_);
  or (_04880_, _04879_, _04876_);
  or (_04881_, _04880_, _04869_);
  or (_04882_, _04881_, _04862_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04882_, _04859_);
  and (_04883_, _04371_, _04609_);
  and (_04884_, _04375_, _04592_);
  or (_04885_, _04884_, _04883_);
  and (_04886_, _04380_, _04611_);
  and (_04887_, _04384_, _04594_);
  or (_04888_, _04887_, _04886_);
  or (_04889_, _04888_, _04885_);
  and (_04890_, _04392_, _04589_);
  and (_04891_, _04389_, _04598_);
  or (_04892_, _04891_, _04890_);
  and (_04893_, _04409_, _04576_);
  and (_04894_, _04398_, _04581_);
  or (_04895_, _04894_, _04893_);
  and (_04896_, _04401_, _04604_);
  and (_04897_, _04430_, _04617_);
  or (_04898_, _04897_, _04896_);
  or (_04899_, _04898_, _04895_);
  and (_04900_, _04414_, _04587_);
  and (_04901_, _04367_, _04583_);
  and (_04902_, _04424_, _04578_);
  and (_04903_, _04421_, _04619_);
  or (_04904_, _04903_, _04902_);
  or (_04905_, _04904_, _04901_);
  or (_04906_, _04905_, _04900_);
  and (_04907_, _04406_, _04600_);
  and (_04908_, _04433_, _04602_);
  or (_04909_, _04908_, _04907_);
  or (_04910_, _04909_, _04906_);
  or (_04911_, _04910_, _04899_);
  or (_04912_, _04911_, _04892_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04912_, _04889_);
  and (_04913_, _04371_, _04645_);
  and (_04914_, _04375_, _04650_);
  or (_04915_, _04914_, _04913_);
  and (_04916_, _04380_, _04652_);
  and (_04917_, _04384_, _04634_);
  or (_04918_, _04917_, _04916_);
  or (_04919_, _04918_, _04915_);
  and (_04920_, _04392_, _04637_);
  and (_04921_, _04389_, _04639_);
  or (_04922_, _04921_, _04920_);
  and (_04923_, _04409_, _04658_);
  and (_04924_, _04398_, _04661_);
  or (_04925_, _04924_, _04923_);
  and (_04926_, _04401_, _04663_);
  and (_04927_, _04430_, _04627_);
  or (_04928_, _04927_, _04926_);
  or (_04929_, _04928_, _04925_);
  and (_04930_, _04414_, _04632_);
  and (_04931_, _04367_, _04625_);
  and (_04932_, _04424_, _04656_);
  and (_04933_, _04421_, _04630_);
  or (_04934_, _04933_, _04932_);
  or (_04935_, _04934_, _04931_);
  or (_04936_, _04935_, _04930_);
  and (_04937_, _04406_, _04623_);
  and (_04938_, _04433_, _04647_);
  or (_04939_, _04938_, _04937_);
  or (_04940_, _04939_, _04936_);
  or (_04941_, _04940_, _04929_);
  or (_04942_, _04941_, _04922_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04942_, _04919_);
  and (_04943_, _04375_, _04687_);
  and (_04944_, _04384_, _04709_);
  or (_04945_, _04944_, _04943_);
  and (_04946_, _04380_, _04685_);
  and (_04947_, _04371_, _04707_);
  or (_04948_, _04947_, _04946_);
  or (_04949_, _04948_, _04945_);
  and (_04950_, _04389_, _04696_);
  and (_04951_, _04392_, _04692_);
  or (_04952_, _04951_, _04950_);
  and (_04953_, _04406_, _04698_);
  and (_04954_, _04409_, _04669_);
  or (_04955_, _04954_, _04953_);
  and (_04956_, _04433_, _04700_);
  and (_04957_, _04401_, _04702_);
  or (_04958_, _04957_, _04956_);
  or (_04959_, _04958_, _04955_);
  and (_04960_, _04414_, _04690_);
  and (_04961_, _04421_, _04682_);
  and (_04962_, _04424_, _04671_);
  and (_04963_, _04367_, _04676_);
  or (_04964_, _04963_, _04962_);
  or (_04965_, _04964_, _04961_);
  or (_04966_, _04965_, _04960_);
  and (_04967_, _04398_, _04674_);
  and (_04968_, _04430_, _04680_);
  or (_04969_, _04968_, _04967_);
  or (_04970_, _04969_, _04966_);
  or (_04971_, _04970_, _04959_);
  or (_04972_, _04971_, _04952_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04972_, _04949_);
  and (_04973_, _04375_, _04742_);
  and (_04974_, _04384_, _04726_);
  or (_04975_, _04974_, _04973_);
  and (_04976_, _04380_, _04744_);
  and (_04977_, _04371_, _04737_);
  or (_04978_, _04977_, _04976_);
  or (_04979_, _04978_, _04975_);
  and (_04980_, _04389_, _04731_);
  and (_04981_, _04392_, _04729_);
  or (_04982_, _04981_, _04980_);
  and (_04983_, _04406_, _04715_);
  and (_04984_, _04409_, _04750_);
  or (_04985_, _04984_, _04983_);
  and (_04986_, _04433_, _04739_);
  and (_04987_, _04401_, _04755_);
  or (_04988_, _04987_, _04986_);
  or (_04989_, _04988_, _04985_);
  and (_04990_, _04414_, _04724_);
  and (_04991_, _04421_, _04722_);
  and (_04992_, _04424_, _04748_);
  and (_04993_, _04367_, _04717_);
  or (_04994_, _04993_, _04992_);
  or (_04995_, _04994_, _04991_);
  or (_04996_, _04995_, _04990_);
  and (_04997_, _04398_, _04753_);
  and (_04998_, _04430_, _04719_);
  or (_04999_, _04998_, _04997_);
  or (_05000_, _04999_, _04996_);
  or (_05001_, _05000_, _04989_);
  or (_05002_, _05001_, _04982_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _05002_, _04979_);
  and (_05003_, _04371_, _04772_);
  and (_05004_, _04375_, _04777_);
  or (_05005_, _05004_, _05003_);
  and (_05006_, _04380_, _04794_);
  and (_05007_, _04384_, _04774_);
  or (_05008_, _05007_, _05006_);
  or (_05009_, _05008_, _05005_);
  and (_05010_, _04392_, _04796_);
  and (_05011_, _04389_, _04783_);
  or (_05012_, _05011_, _05010_);
  and (_05013_, _04409_, _04761_);
  and (_05014_, _04398_, _04766_);
  or (_05015_, _05014_, _05013_);
  and (_05016_, _04401_, _04785_);
  and (_05017_, _04430_, _04801_);
  or (_05018_, _05017_, _05016_);
  or (_05019_, _05018_, _05015_);
  and (_05020_, _04414_, _04779_);
  and (_05021_, _04367_, _04768_);
  and (_05022_, _04424_, _04763_);
  and (_05023_, _04421_, _04803_);
  or (_05024_, _05023_, _05022_);
  or (_05025_, _05024_, _05021_);
  or (_05026_, _05025_, _05020_);
  and (_05027_, _04406_, _04787_);
  and (_05028_, _04433_, _04789_);
  or (_05029_, _05028_, _05027_);
  or (_05030_, _05029_, _05026_);
  or (_05031_, _05030_, _05019_);
  or (_05032_, _05031_, _05012_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _05032_, _05009_);
  and (_05033_, _04371_, _04820_);
  and (_05034_, _04375_, _04825_);
  or (_05035_, _05034_, _05033_);
  and (_05036_, _04380_, _04842_);
  and (_05037_, _04384_, _04840_);
  or (_05038_, _05037_, _05036_);
  or (_05039_, _05038_, _05035_);
  and (_05040_, _04392_, _04818_);
  and (_05041_, _04389_, _04829_);
  or (_05042_, _05041_, _05040_);
  and (_05043_, _04409_, _04812_);
  and (_05044_, _04398_, _04814_);
  or (_05045_, _05044_, _05043_);
  and (_05046_, _04401_, _04831_);
  and (_05047_, _04430_, _04847_);
  or (_05048_, _05047_, _05046_);
  or (_05049_, _05048_, _05045_);
  and (_05050_, _04414_, _04823_);
  and (_05051_, _04367_, _04807_);
  and (_05052_, _04424_, _04809_);
  and (_05053_, _04421_, _04849_);
  or (_05054_, _05053_, _05052_);
  or (_05055_, _05054_, _05051_);
  or (_05056_, _05055_, _05050_);
  and (_05057_, _04406_, _04833_);
  and (_05059_, _04433_, _04835_);
  or (_05061_, _05059_, _05057_);
  or (_05063_, _05061_, _05056_);
  or (_05065_, _05063_, _05049_);
  or (_05067_, _05065_, _05042_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _05067_, _05039_);
  and (_05070_, _04375_, _04530_);
  and (_05071_, _04380_, _04532_);
  or (_05072_, _05071_, _05070_);
  and (_05073_, _04371_, _04546_);
  and (_05074_, _04384_, _04552_);
  or (_05075_, _05074_, _05073_);
  or (_05076_, _05075_, _05072_);
  and (_05078_, _04389_, _04572_);
  and (_05079_, _04392_, _04537_);
  or (_05081_, _05079_, _05078_);
  and (_05082_, _04406_, _04541_);
  and (_05083_, _04409_, _04558_);
  or (_05085_, _05083_, _05082_);
  and (_05086_, _04430_, _04556_);
  and (_05087_, _04401_, _04543_);
  or (_05089_, _05087_, _05086_);
  or (_05090_, _05089_, _05085_);
  and (_05091_, _04414_, _04565_);
  and (_05093_, _04424_, _04535_);
  and (_05094_, _04421_, _04554_);
  and (_05095_, _04367_, _04570_);
  or (_05097_, _05095_, _05094_);
  or (_05098_, _05097_, _05093_);
  or (_05099_, _05098_, _05091_);
  and (_05101_, _04433_, _04563_);
  and (_05102_, _04398_, _04548_);
  or (_05103_, _05102_, _05101_);
  or (_05105_, _05103_, _05099_);
  or (_05106_, _05105_, _05090_);
  or (_05107_, _05106_, _05081_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05107_, _05076_);
  and (_05109_, _04371_, _04592_);
  and (_05110_, _04375_, _04576_);
  or (_05111_, _05110_, _05109_);
  and (_05112_, _04380_, _04578_);
  and (_05113_, _04384_, _04598_);
  or (_05114_, _05113_, _05112_);
  or (_05115_, _05114_, _05111_);
  and (_05116_, _04389_, _04619_);
  and (_05117_, _04392_, _04583_);
  or (_05118_, _05117_, _05116_);
  and (_05119_, _04401_, _04594_);
  and (_05120_, _04398_, _04587_);
  or (_05121_, _05120_, _05119_);
  and (_05122_, _04406_, _04609_);
  and (_05123_, _04409_, _04604_);
  or (_05124_, _05123_, _05122_);
  or (_05125_, _05124_, _05121_);
  and (_05126_, _04414_, _04589_);
  and (_05127_, _04367_, _04617_);
  and (_05128_, _04421_, _04600_);
  and (_05130_, _04424_, _04581_);
  or (_05131_, _05130_, _05128_);
  or (_05133_, _05131_, _05127_);
  or (_05134_, _05133_, _05126_);
  and (_05135_, _04430_, _04602_);
  and (_05137_, _04433_, _04611_);
  or (_05138_, _05137_, _05135_);
  or (_05139_, _05138_, _05134_);
  or (_05141_, _05139_, _05125_);
  or (_05142_, _05141_, _05118_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05142_, _05115_);
  and (_05144_, _04371_, _04650_);
  and (_05145_, _04380_, _04656_);
  or (_05146_, _05145_, _05144_);
  and (_05148_, _04375_, _04658_);
  and (_05149_, _04384_, _04639_);
  or (_05150_, _05149_, _05148_);
  or (_05152_, _05150_, _05146_);
  and (_05153_, _04389_, _04630_);
  and (_05154_, _04392_, _04625_);
  or (_05156_, _05154_, _05153_);
  and (_05157_, _04430_, _04647_);
  and (_05158_, _04409_, _04663_);
  or (_05160_, _05158_, _05157_);
  and (_05161_, _04433_, _04652_);
  and (_05162_, _04401_, _04634_);
  or (_05163_, _05162_, _05161_);
  or (_05164_, _05163_, _05160_);
  and (_05165_, _04414_, _04637_);
  and (_05166_, _04424_, _04661_);
  and (_05167_, _04421_, _04623_);
  and (_05168_, _04367_, _04627_);
  or (_05169_, _05168_, _05167_);
  or (_05170_, _05169_, _05166_);
  or (_05171_, _05170_, _05165_);
  and (_05172_, _04406_, _04645_);
  and (_05173_, _04398_, _04632_);
  or (_05174_, _05173_, _05172_);
  or (_05175_, _05174_, _05171_);
  or (_05176_, _05175_, _05164_);
  or (_05177_, _05176_, _05156_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05177_, _05152_);
  and (_05178_, _04375_, _04669_);
  and (_05179_, _04380_, _04671_);
  or (_05181_, _05179_, _05178_);
  and (_05182_, _04371_, _04687_);
  and (_05184_, _04384_, _04696_);
  or (_05185_, _05184_, _05182_);
  or (_05186_, _05185_, _05181_);
  and (_05188_, _04389_, _04682_);
  and (_05189_, _04392_, _04676_);
  or (_05190_, _05189_, _05188_);
  and (_05192_, _04398_, _04690_);
  and (_05193_, _04401_, _04709_);
  or (_05194_, _05193_, _05192_);
  and (_05196_, _04406_, _04707_);
  and (_05197_, _04409_, _04702_);
  or (_05198_, _05197_, _05196_);
  or (_05200_, _05198_, _05194_);
  and (_05201_, _04414_, _04692_);
  and (_05202_, _04367_, _04680_);
  and (_05204_, _04421_, _04698_);
  and (_05205_, _04424_, _04674_);
  or (_05206_, _05205_, _05204_);
  or (_05208_, _05206_, _05202_);
  or (_05209_, _05208_, _05201_);
  and (_05210_, _04430_, _04700_);
  and (_05212_, _04433_, _04685_);
  or (_05213_, _05212_, _05210_);
  or (_05214_, _05213_, _05209_);
  or (_05215_, _05214_, _05200_);
  or (_05216_, _05215_, _05190_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05216_, _05186_);
  and (_05217_, _04371_, _04742_);
  and (_05218_, _04375_, _04750_);
  or (_05219_, _05218_, _05217_);
  and (_05220_, _04380_, _04748_);
  and (_05221_, _04384_, _04731_);
  or (_05222_, _05221_, _05220_);
  or (_05223_, _05222_, _05219_);
  and (_05224_, _04389_, _04722_);
  and (_05225_, _04392_, _04717_);
  or (_05226_, _05225_, _05224_);
  and (_05227_, _04401_, _04726_);
  and (_05228_, _04398_, _04724_);
  or (_05229_, _05228_, _05227_);
  and (_05230_, _04406_, _04737_);
  and (_05231_, _04409_, _04755_);
  or (_05233_, _05231_, _05230_);
  or (_05234_, _05233_, _05229_);
  and (_05236_, _04414_, _04729_);
  and (_05237_, _04367_, _04719_);
  and (_05238_, _04421_, _04715_);
  and (_05240_, _04424_, _04753_);
  or (_05241_, _05240_, _05238_);
  or (_05242_, _05241_, _05237_);
  or (_05244_, _05242_, _05236_);
  and (_05245_, _04430_, _04739_);
  and (_05246_, _04433_, _04744_);
  or (_05248_, _05246_, _05245_);
  or (_05249_, _05248_, _05244_);
  or (_05250_, _05249_, _05234_);
  or (_05252_, _05250_, _05226_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05252_, _05223_);
  and (_05253_, _04371_, _04777_);
  and (_05255_, _04375_, _04761_);
  or (_05256_, _05255_, _05253_);
  and (_05257_, _04380_, _04763_);
  and (_05259_, _04384_, _04783_);
  or (_05260_, _05259_, _05257_);
  or (_05261_, _05260_, _05256_);
  and (_05263_, _04389_, _04803_);
  and (_05264_, _04392_, _04768_);
  or (_05265_, _05264_, _05263_);
  and (_05266_, _04401_, _04774_);
  and (_05267_, _04398_, _04779_);
  or (_05268_, _05267_, _05266_);
  and (_05269_, _04406_, _04772_);
  and (_05270_, _04409_, _04785_);
  or (_05271_, _05270_, _05269_);
  or (_05272_, _05271_, _05268_);
  and (_05273_, _04414_, _04796_);
  and (_05274_, _04367_, _04801_);
  and (_05275_, _04421_, _04787_);
  and (_05276_, _04424_, _04766_);
  or (_05277_, _05276_, _05275_);
  or (_05278_, _05277_, _05274_);
  or (_05279_, _05278_, _05273_);
  and (_05280_, _04430_, _04789_);
  and (_05281_, _04433_, _04794_);
  or (_05282_, _05281_, _05280_);
  or (_05283_, _05282_, _05279_);
  or (_05285_, _05283_, _05272_);
  or (_05286_, _05285_, _05265_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05286_, _05261_);
  and (_05288_, _04371_, _04825_);
  and (_05289_, _04375_, _04812_);
  or (_05291_, _05289_, _05288_);
  and (_05292_, _04380_, _04809_);
  and (_05293_, _04384_, _04829_);
  or (_05295_, _05293_, _05292_);
  or (_05296_, _05295_, _05291_);
  and (_05297_, _04389_, _04849_);
  and (_05299_, _04392_, _04807_);
  or (_05300_, _05299_, _05297_);
  and (_05301_, _04401_, _04840_);
  and (_05303_, _04398_, _04823_);
  or (_05304_, _05303_, _05301_);
  and (_05305_, _04406_, _04820_);
  and (_05307_, _04409_, _04831_);
  or (_05308_, _05307_, _05305_);
  or (_05309_, _05308_, _05304_);
  and (_05311_, _04414_, _04818_);
  and (_05312_, _04367_, _04847_);
  and (_05313_, _04421_, _04833_);
  and (_05315_, _04424_, _04814_);
  or (_05316_, _05315_, _05313_);
  or (_05317_, _05316_, _05312_);
  or (_05318_, _05317_, _05311_);
  and (_05319_, _04430_, _04835_);
  and (_05320_, _04433_, _04842_);
  or (_05321_, _05320_, _05319_);
  or (_05322_, _05321_, _05318_);
  or (_05323_, _05322_, _05309_);
  or (_05324_, _05323_, _05300_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05324_, _05296_);
  and (_05325_, _04371_, _04563_);
  and (_05326_, _04380_, _04546_);
  or (_05327_, _05326_, _05325_);
  and (_05328_, _04375_, _04532_);
  and (_05329_, _04384_, _04565_);
  or (_05330_, _05329_, _05328_);
  or (_05331_, _05330_, _05327_);
  and (_05332_, _04409_, _04535_);
  and (_05333_, _04401_, _04548_);
  or (_05334_, _05333_, _05332_);
  and (_05336_, _04433_, _04541_);
  and (_05337_, _04398_, _04558_);
  or (_05339_, _05337_, _05336_);
  or (_05340_, _05339_, _05334_);
  and (_05341_, _04414_, _04543_);
  and (_05343_, _04424_, _04530_);
  and (_05344_, _04421_, _04570_);
  and (_05345_, _04367_, _04572_);
  or (_05347_, _05345_, _05344_);
  or (_05348_, _05347_, _05343_);
  or (_05349_, _05348_, _05341_);
  and (_05351_, _04430_, _04554_);
  and (_05352_, _04406_, _04556_);
  or (_05353_, _05352_, _05351_);
  or (_05355_, _05353_, _05349_);
  or (_05356_, _05355_, _05340_);
  and (_05357_, _04392_, _04552_);
  and (_05359_, _04389_, _04537_);
  or (_05360_, _05359_, _05357_);
  or (_05361_, _05360_, _05356_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _05361_, _05331_);
  and (_05363_, _04371_, _04611_);
  and (_05364_, _04380_, _04592_);
  or (_05366_, _05364_, _05363_);
  and (_05367_, _04375_, _04578_);
  and (_05368_, _04384_, _04589_);
  or (_05369_, _05368_, _05367_);
  or (_05370_, _05369_, _05366_);
  and (_05371_, _04409_, _04581_);
  and (_05372_, _04401_, _04587_);
  or (_05373_, _05372_, _05371_);
  and (_05374_, _04433_, _04609_);
  and (_05375_, _04398_, _04604_);
  or (_05376_, _05375_, _05374_);
  or (_05377_, _05376_, _05373_);
  and (_05378_, _04414_, _04594_);
  and (_05379_, _04424_, _04576_);
  and (_05380_, _04421_, _04617_);
  and (_05381_, _04367_, _04619_);
  or (_05382_, _05381_, _05380_);
  or (_05383_, _05382_, _05379_);
  or (_05384_, _05383_, _05378_);
  and (_05385_, _04430_, _04600_);
  and (_05386_, _04406_, _04602_);
  or (_05388_, _05386_, _05385_);
  or (_05389_, _05388_, _05384_);
  or (_05391_, _05389_, _05377_);
  and (_05392_, _04392_, _04598_);
  and (_05393_, _04389_, _04583_);
  or (_05395_, _05393_, _05392_);
  or (_05396_, _05395_, _05391_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _05396_, _05370_);
  and (_05398_, _04371_, _04652_);
  and (_05399_, _04375_, _04656_);
  or (_05400_, _05399_, _05398_);
  and (_05402_, _04380_, _04650_);
  and (_05403_, _04384_, _04637_);
  or (_05404_, _05403_, _05402_);
  or (_05406_, _05404_, _05400_);
  and (_05407_, _04398_, _04663_);
  and (_05408_, _04401_, _04632_);
  or (_05410_, _05408_, _05407_);
  and (_05411_, _04406_, _04647_);
  and (_05412_, _04409_, _04661_);
  or (_05414_, _05412_, _05411_);
  or (_05415_, _05414_, _05410_);
  and (_05416_, _04414_, _04634_);
  and (_05418_, _04367_, _04630_);
  and (_05419_, _04424_, _04658_);
  and (_05420_, _04421_, _04627_);
  or (_05421_, _05420_, _05419_);
  or (_05422_, _05421_, _05418_);
  or (_05423_, _05422_, _05416_);
  and (_05424_, _04430_, _04623_);
  and (_05425_, _04433_, _04645_);
  or (_05426_, _05425_, _05424_);
  or (_05427_, _05426_, _05423_);
  or (_05428_, _05427_, _05415_);
  and (_05429_, _04392_, _04639_);
  and (_05430_, _04389_, _04625_);
  or (_05431_, _05430_, _05429_);
  or (_05432_, _05431_, _05428_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _05432_, _05406_);
  and (_05433_, _04371_, _04685_);
  and (_05434_, _04375_, _04671_);
  or (_05435_, _05434_, _05433_);
  and (_05436_, _04380_, _04687_);
  and (_05437_, _04384_, _04692_);
  or (_05439_, _05437_, _05436_);
  or (_05440_, _05439_, _05435_);
  and (_05442_, _04398_, _04702_);
  and (_05443_, _04401_, _04690_);
  or (_05444_, _05443_, _05442_);
  and (_05446_, _04406_, _04700_);
  and (_05447_, _04409_, _04674_);
  or (_05448_, _05447_, _05446_);
  or (_05450_, _05448_, _05444_);
  and (_05451_, _04414_, _04709_);
  and (_05452_, _04367_, _04682_);
  and (_05454_, _04424_, _04669_);
  and (_05455_, _04421_, _04680_);
  or (_05456_, _05455_, _05454_);
  or (_05458_, _05456_, _05452_);
  or (_05459_, _05458_, _05451_);
  and (_05460_, _04430_, _04698_);
  and (_05462_, _04433_, _04707_);
  or (_05463_, _05462_, _05460_);
  or (_05464_, _05463_, _05459_);
  or (_05466_, _05464_, _05450_);
  and (_05467_, _04392_, _04696_);
  and (_05468_, _04389_, _04676_);
  or (_05470_, _05468_, _05467_);
  or (_05471_, _05470_, _05466_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _05471_, _05440_);
  and (_05472_, _04371_, _04744_);
  and (_05473_, _04375_, _04748_);
  or (_05474_, _05473_, _05472_);
  and (_05475_, _04380_, _04742_);
  and (_05476_, _04384_, _04729_);
  or (_05477_, _05476_, _05475_);
  or (_05478_, _05477_, _05474_);
  and (_05479_, _04398_, _04755_);
  and (_05480_, _04401_, _04724_);
  or (_05481_, _05480_, _05479_);
  and (_05482_, _04406_, _04739_);
  and (_05483_, _04409_, _04753_);
  or (_05484_, _05483_, _05482_);
  or (_05485_, _05484_, _05481_);
  and (_05486_, _04414_, _04726_);
  and (_05487_, _04367_, _04722_);
  and (_05488_, _04424_, _04750_);
  and (_05489_, _04421_, _04719_);
  or (_05491_, _05489_, _05488_);
  or (_05492_, _05491_, _05487_);
  or (_05494_, _05492_, _05486_);
  and (_05495_, _04430_, _04715_);
  and (_05496_, _04433_, _04737_);
  or (_05498_, _05496_, _05495_);
  or (_05499_, _05498_, _05494_);
  or (_05500_, _05499_, _05485_);
  and (_05502_, _04392_, _04731_);
  and (_05503_, _04389_, _04717_);
  or (_05504_, _05503_, _05502_);
  or (_05506_, _05504_, _05500_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _05506_, _05478_);
  and (_05507_, _04380_, _04777_);
  and (_05509_, _04371_, _04794_);
  or (_05510_, _05509_, _05507_);
  and (_05511_, _04375_, _04763_);
  and (_05513_, _04384_, _04796_);
  or (_05514_, _05513_, _05511_);
  or (_05515_, _05514_, _05510_);
  and (_05517_, _04398_, _04785_);
  and (_05518_, _04401_, _04779_);
  or (_05519_, _05518_, _05517_);
  and (_05521_, _04430_, _04787_);
  and (_05522_, _04433_, _04772_);
  or (_05523_, _05522_, _05521_);
  or (_05524_, _05523_, _05519_);
  and (_05525_, _04414_, _04774_);
  and (_05526_, _04421_, _04801_);
  and (_05527_, _04424_, _04761_);
  and (_05528_, _04367_, _04803_);
  or (_05529_, _05528_, _05527_);
  or (_05530_, _05529_, _05526_);
  or (_05531_, _05530_, _05525_);
  and (_05532_, _04406_, _04789_);
  and (_05533_, _04409_, _04766_);
  or (_05534_, _05533_, _05532_);
  or (_05535_, _05534_, _05531_);
  or (_05536_, _05535_, _05524_);
  and (_05537_, _04392_, _04783_);
  and (_05538_, _04389_, _04768_);
  or (_05539_, _05538_, _05537_);
  or (_05540_, _05539_, _05536_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _05540_, _05515_);
  and (_05542_, _04371_, _04842_);
  and (_05543_, _04375_, _04809_);
  or (_05545_, _05543_, _05542_);
  and (_05546_, _04380_, _04825_);
  and (_05547_, _04384_, _04818_);
  or (_05549_, _05547_, _05546_);
  or (_05550_, _05549_, _05545_);
  and (_05551_, _04398_, _04831_);
  and (_05553_, _04401_, _04823_);
  or (_05554_, _05553_, _05551_);
  and (_05555_, _04406_, _04835_);
  and (_05557_, _04409_, _04814_);
  or (_05558_, _05557_, _05555_);
  or (_05559_, _05558_, _05554_);
  and (_05561_, _04414_, _04840_);
  and (_05562_, _04367_, _04849_);
  and (_05563_, _04424_, _04812_);
  and (_05565_, _04421_, _04847_);
  or (_05566_, _05565_, _05563_);
  or (_05567_, _05566_, _05562_);
  or (_05569_, _05567_, _05561_);
  and (_05570_, _04430_, _04833_);
  and (_05571_, _04433_, _04820_);
  or (_05573_, _05571_, _05570_);
  or (_05574_, _05573_, _05569_);
  or (_05575_, _05574_, _05559_);
  and (_05576_, _04392_, _04829_);
  and (_05577_, _04389_, _04807_);
  or (_05578_, _05577_, _05576_);
  or (_05579_, _05578_, _05575_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _05579_, _05550_);
  nand (_05580_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_05581_, \oc8051_golden_model_1.PC [3]);
  or (_05582_, \oc8051_golden_model_1.PC [2], _05581_);
  or (_05583_, _05582_, _05580_);
  or (_05584_, _05583_, _00436_);
  not (_05585_, \oc8051_golden_model_1.PC [1]);
  or (_05586_, _05585_, \oc8051_golden_model_1.PC [0]);
  or (_05587_, _05586_, _05582_);
  or (_05588_, _05587_, _00395_);
  and (_05589_, _05588_, _05584_);
  not (_05590_, \oc8051_golden_model_1.PC [2]);
  or (_05591_, _05590_, \oc8051_golden_model_1.PC [3]);
  or (_05592_, _05591_, _05580_);
  or (_05594_, _05592_, _00272_);
  or (_05595_, _05591_, _05586_);
  or (_05597_, _05595_, _00231_);
  and (_05598_, _05597_, _05594_);
  and (_05599_, _05598_, _05589_);
  nand (_05601_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05602_, _05601_, _05580_);
  or (_05603_, _05602_, _00619_);
  or (_05605_, _05601_, _05586_);
  or (_05606_, _05605_, _00569_);
  and (_05607_, _05606_, _05603_);
  or (_05609_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_05610_, _05609_, _05580_);
  or (_05611_, _05610_, _00077_);
  or (_05613_, _05609_, _05586_);
  or (_05614_, _05613_, _00036_);
  and (_05615_, _05614_, _05611_);
  and (_05617_, _05615_, _05607_);
  and (_05618_, _05617_, _05599_);
  not (_05619_, \oc8051_golden_model_1.PC [0]);
  or (_05621_, \oc8051_golden_model_1.PC [1], _05619_);
  or (_05622_, _05621_, _05601_);
  or (_05623_, _05622_, _00518_);
  or (_05625_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_05626_, _05625_, _05601_);
  or (_05627_, _05626_, _00477_);
  and (_05628_, _05627_, _05623_);
  or (_05629_, _05609_, _05625_);
  or (_05630_, _05629_, _43220_);
  or (_05631_, _05609_, _05621_);
  or (_05632_, _05631_, _43261_);
  and (_05633_, _05632_, _05630_);
  and (_05634_, _05633_, _05628_);
  or (_05635_, _05621_, _05582_);
  or (_05636_, _05635_, _00354_);
  or (_05637_, _05625_, _05582_);
  or (_05638_, _05637_, _00313_);
  and (_05639_, _05638_, _05636_);
  or (_05640_, _05621_, _05591_);
  or (_05641_, _05640_, _00190_);
  or (_05642_, _05625_, _05591_);
  or (_05643_, _05642_, _00118_);
  and (_05644_, _05643_, _05641_);
  and (_05645_, _05644_, _05639_);
  and (_05647_, _05645_, _05634_);
  and (_05648_, _05647_, _05618_);
  or (_05650_, _05583_, _00401_);
  or (_05651_, _05587_, _00360_);
  and (_05652_, _05651_, _05650_);
  or (_05654_, _05592_, _00237_);
  or (_05655_, _05595_, _00196_);
  and (_05656_, _05655_, _05654_);
  and (_05658_, _05656_, _05652_);
  or (_05659_, _05602_, _00579_);
  or (_05660_, _05605_, _00524_);
  and (_05662_, _05660_, _05659_);
  or (_05663_, _05610_, _00042_);
  or (_05664_, _05613_, _43267_);
  and (_05666_, _05664_, _05663_);
  and (_05667_, _05666_, _05662_);
  and (_05668_, _05667_, _05658_);
  or (_05670_, _05622_, _00483_);
  or (_05671_, _05626_, _00442_);
  and (_05672_, _05671_, _05670_);
  or (_05674_, _05629_, _43185_);
  or (_05675_, _05631_, _43226_);
  and (_05676_, _05675_, _05674_);
  and (_05678_, _05676_, _05672_);
  or (_05679_, _05635_, _00319_);
  or (_05680_, _05637_, _00278_);
  and (_05681_, _05680_, _05679_);
  or (_05682_, _05640_, _00124_);
  or (_05683_, _05642_, _00083_);
  and (_05684_, _05683_, _05682_);
  and (_05685_, _05684_, _05681_);
  and (_05686_, _05685_, _05678_);
  and (_05687_, _05686_, _05668_);
  and (_05688_, _05687_, _05648_);
  or (_05689_, _05583_, _00426_);
  or (_05690_, _05587_, _00385_);
  and (_05691_, _05690_, _05689_);
  or (_05692_, _05592_, _00262_);
  or (_05693_, _05595_, _00221_);
  and (_05694_, _05693_, _05692_);
  and (_05695_, _05694_, _05691_);
  or (_05696_, _05602_, _00609_);
  or (_05697_, _05605_, _00553_);
  and (_05698_, _05697_, _05696_);
  or (_05700_, _05610_, _00067_);
  or (_05701_, _05613_, _00026_);
  and (_05703_, _05701_, _05700_);
  and (_05704_, _05703_, _05698_);
  and (_05705_, _05704_, _05695_);
  or (_05707_, _05622_, _00508_);
  or (_05708_, _05626_, _00467_);
  and (_05709_, _05708_, _05707_);
  or (_05711_, _05629_, _43210_);
  or (_05712_, _05631_, _43251_);
  and (_05713_, _05712_, _05711_);
  and (_05715_, _05713_, _05709_);
  or (_05716_, _05635_, _00344_);
  or (_05717_, _05637_, _00303_);
  and (_05719_, _05717_, _05716_);
  or (_05720_, _05640_, _00172_);
  or (_05721_, _05642_, _00108_);
  and (_05723_, _05721_, _05720_);
  and (_05724_, _05723_, _05719_);
  and (_05725_, _05724_, _05715_);
  nand (_05727_, _05725_, _05705_);
  or (_05728_, _05583_, _00431_);
  or (_05729_, _05587_, _00390_);
  and (_05731_, _05729_, _05728_);
  or (_05732_, _05592_, _00267_);
  or (_05733_, _05595_, _00226_);
  and (_05734_, _05733_, _05732_);
  and (_05735_, _05734_, _05731_);
  or (_05736_, _05602_, _00614_);
  or (_05737_, _05605_, _00561_);
  and (_05738_, _05737_, _05736_);
  or (_05739_, _05610_, _00072_);
  or (_05740_, _05613_, _00031_);
  and (_05741_, _05740_, _05739_);
  and (_05742_, _05741_, _05738_);
  and (_05743_, _05742_, _05735_);
  or (_05744_, _05622_, _00513_);
  or (_05745_, _05626_, _00472_);
  and (_05746_, _05745_, _05744_);
  or (_05747_, _05629_, _43215_);
  or (_05748_, _05631_, _43256_);
  and (_05749_, _05748_, _05747_);
  and (_05750_, _05749_, _05746_);
  or (_05751_, _05635_, _00349_);
  or (_05753_, _05637_, _00308_);
  and (_05754_, _05753_, _05751_);
  or (_05756_, _05640_, _00183_);
  or (_05757_, _05642_, _00113_);
  and (_05758_, _05757_, _05756_);
  and (_05760_, _05758_, _05754_);
  and (_05761_, _05760_, _05750_);
  nand (_05762_, _05761_, _05743_);
  or (_05764_, _05762_, _05727_);
  not (_05765_, _05764_);
  and (_05766_, _05765_, _05688_);
  or (_05768_, _05583_, _00406_);
  or (_05769_, _05587_, _00365_);
  and (_05770_, _05769_, _05768_);
  or (_05772_, _05592_, _00242_);
  or (_05773_, _05595_, _00201_);
  and (_05774_, _05773_, _05772_);
  and (_05776_, _05774_, _05770_);
  or (_05777_, _05602_, _00587_);
  or (_05778_, _05605_, _00529_);
  and (_05780_, _05778_, _05777_);
  or (_05781_, _05610_, _00047_);
  or (_05782_, _05613_, _00006_);
  and (_05784_, _05782_, _05781_);
  and (_05785_, _05784_, _05780_);
  and (_05786_, _05785_, _05776_);
  or (_05787_, _05622_, _00488_);
  or (_05788_, _05626_, _00447_);
  and (_05789_, _05788_, _05787_);
  or (_05790_, _05629_, _43190_);
  or (_05791_, _05631_, _43231_);
  and (_05792_, _05791_, _05790_);
  and (_05793_, _05792_, _05789_);
  or (_05794_, _05635_, _00324_);
  or (_05795_, _05637_, _00283_);
  and (_05796_, _05795_, _05794_);
  or (_05797_, _05640_, _00129_);
  or (_05798_, _05642_, _00088_);
  and (_05799_, _05798_, _05797_);
  and (_05800_, _05799_, _05796_);
  and (_05801_, _05800_, _05793_);
  and (_05802_, _05801_, _05786_);
  or (_05803_, _05583_, _00416_);
  or (_05804_, _05587_, _00375_);
  and (_05806_, _05804_, _05803_);
  or (_05807_, _05592_, _00252_);
  or (_05809_, _05595_, _00211_);
  and (_05810_, _05809_, _05807_);
  and (_05811_, _05810_, _05806_);
  or (_05813_, _05602_, _00599_);
  or (_05814_, _05605_, _00539_);
  and (_05815_, _05814_, _05813_);
  or (_05817_, _05610_, _00057_);
  or (_05818_, _05613_, _00016_);
  and (_05819_, _05818_, _05817_);
  and (_05821_, _05819_, _05815_);
  and (_05822_, _05821_, _05811_);
  or (_05823_, _05622_, _00498_);
  or (_05825_, _05626_, _00457_);
  and (_05826_, _05825_, _05823_);
  or (_05827_, _05629_, _43200_);
  or (_05829_, _05631_, _43241_);
  and (_05830_, _05829_, _05827_);
  and (_05831_, _05830_, _05826_);
  or (_05833_, _05635_, _00334_);
  or (_05834_, _05637_, _00293_);
  and (_05835_, _05834_, _05833_);
  or (_05837_, _05640_, _00150_);
  or (_05838_, _05642_, _00098_);
  and (_05839_, _05838_, _05837_);
  and (_05840_, _05839_, _05835_);
  and (_05841_, _05840_, _05831_);
  nand (_05842_, _05841_, _05822_);
  or (_05843_, _05583_, _00421_);
  or (_05844_, _05587_, _00380_);
  and (_05845_, _05844_, _05843_);
  or (_05846_, _05592_, _00257_);
  or (_05847_, _05595_, _00216_);
  and (_05848_, _05847_, _05846_);
  and (_05849_, _05848_, _05845_);
  or (_05850_, _05602_, _00604_);
  or (_05851_, _05605_, _00545_);
  and (_05852_, _05851_, _05850_);
  or (_05853_, _05610_, _00062_);
  or (_05854_, _05613_, _00021_);
  and (_05855_, _05854_, _05853_);
  and (_05856_, _05855_, _05852_);
  and (_05857_, _05856_, _05849_);
  or (_05859_, _05622_, _00503_);
  or (_05860_, _05626_, _00462_);
  and (_05862_, _05860_, _05859_);
  or (_05863_, _05629_, _43205_);
  or (_05864_, _05631_, _43246_);
  and (_05866_, _05864_, _05863_);
  and (_05867_, _05866_, _05862_);
  or (_05868_, _05635_, _00339_);
  or (_05870_, _05637_, _00298_);
  and (_05871_, _05870_, _05868_);
  or (_05872_, _05640_, _00161_);
  or (_05874_, _05642_, _00103_);
  and (_05875_, _05874_, _05872_);
  and (_05876_, _05875_, _05871_);
  and (_05878_, _05876_, _05867_);
  nand (_05879_, _05878_, _05857_);
  not (_05880_, _05879_);
  nor (_05882_, _05880_, _05842_);
  and (_05883_, _05882_, _05802_);
  and (_05884_, _05883_, _05766_);
  not (_05886_, _05884_);
  and (_05887_, _05879_, _05842_);
  nand (_05888_, _05887_, _05802_);
  not (_05890_, _05888_);
  and (_05891_, _05890_, _05766_);
  and (_05892_, _05725_, _05705_);
  or (_05893_, _05762_, _05892_);
  not (_05894_, _05893_);
  and (_05895_, _05894_, _05688_);
  or (_05896_, _05583_, _00411_);
  or (_05897_, _05587_, _00370_);
  and (_05898_, _05897_, _05896_);
  or (_05899_, _05592_, _00247_);
  or (_05900_, _05595_, _00206_);
  and (_05901_, _05900_, _05899_);
  and (_05902_, _05901_, _05898_);
  or (_05903_, _05602_, _00594_);
  or (_05904_, _05605_, _00534_);
  and (_05905_, _05904_, _05903_);
  or (_05906_, _05610_, _00052_);
  or (_05907_, _05613_, _00011_);
  and (_05908_, _05907_, _05906_);
  and (_05909_, _05908_, _05905_);
  and (_05910_, _05909_, _05902_);
  or (_05911_, _05622_, _00493_);
  or (_05912_, _05626_, _00452_);
  and (_05913_, _05912_, _05911_);
  or (_05914_, _05629_, _43195_);
  or (_05915_, _05631_, _43236_);
  and (_05916_, _05915_, _05914_);
  and (_05917_, _05916_, _05913_);
  or (_05918_, _05635_, _00329_);
  or (_05919_, _05637_, _00288_);
  and (_05920_, _05919_, _05918_);
  or (_05921_, _05640_, _00139_);
  or (_05922_, _05642_, _00093_);
  and (_05923_, _05922_, _05921_);
  and (_05924_, _05923_, _05920_);
  and (_05925_, _05924_, _05917_);
  nand (_05926_, _05925_, _05910_);
  not (_05927_, _05926_);
  and (_05928_, _05927_, _05802_);
  or (_05929_, _05879_, _05842_);
  not (_05930_, _05929_);
  and (_05931_, _05930_, _05928_);
  and (_05932_, _05931_, _05895_);
  not (_05933_, _05932_);
  or (_05934_, _05927_, _05802_);
  or (_05935_, _05934_, _05929_);
  nand (_05936_, _05647_, _05618_);
  or (_05937_, _05687_, _05936_);
  nor (_05938_, _05937_, _05893_);
  not (_05939_, _05938_);
  or (_05940_, _05939_, _05935_);
  or (_05941_, _05926_, _05802_);
  or (_05942_, _05941_, _05929_);
  and (_05943_, _05761_, _05743_);
  or (_05944_, _05943_, _05892_);
  or (_05945_, _05944_, _05937_);
  or (_05946_, _05945_, _05942_);
  or (_05947_, _05687_, _05648_);
  or (_05948_, _05947_, _05893_);
  or (_05949_, _05948_, _05942_);
  and (_05950_, _05949_, _05946_);
  or (_05951_, _05943_, _05727_);
  or (_05952_, _05951_, _05937_);
  or (_05953_, _05952_, _05942_);
  or (_05954_, _05764_, _05947_);
  or (_05955_, _05954_, _05942_);
  and (_05956_, _05955_, _05953_);
  or (_05957_, _05947_, _05944_);
  or (_05958_, _05957_, _05942_);
  or (_05959_, _05951_, _05947_);
  or (_05960_, _05959_, _05942_);
  and (_05961_, _05960_, _05958_);
  and (_05962_, _05961_, _05956_);
  and (_05963_, _05962_, _05950_);
  or (_05964_, _05963_, _05619_);
  nand (_05965_, _05963_, _05619_);
  nand (_05966_, _05965_, _05964_);
  nand (_05967_, _05966_, _05940_);
  not (_05968_, _05941_);
  and (_05969_, _05880_, _05842_);
  and (_05970_, _05969_, _05968_);
  nor (_05971_, _05764_, _05937_);
  and (_05972_, _05971_, _05970_);
  not (_05973_, _05942_);
  and (_05974_, _05973_, _05938_);
  nor (_05975_, _05974_, _05972_);
  not (_05976_, _05940_);
  and (_05977_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_05978_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_05979_, _05978_, _05977_);
  nand (_05980_, _05979_, _05976_);
  and (_05981_, _05980_, _05975_);
  nand (_05982_, _05981_, _05967_);
  not (_05983_, _05971_);
  nor (_05984_, _05983_, _05935_);
  not (_05985_, _05984_);
  or (_05986_, _05975_, \oc8051_golden_model_1.PC [0]);
  and (_05987_, _05986_, _05985_);
  nand (_05988_, _05987_, _05982_);
  and (_05989_, _05766_, _05973_);
  not (_05990_, _05989_);
  and (_05991_, _05973_, _05895_);
  not (_05992_, _05951_);
  and (_05993_, _05992_, _05688_);
  and (_05994_, _05993_, _05973_);
  nor (_05995_, _05994_, _05991_);
  and (_05996_, _05995_, _05990_);
  and (_05997_, _05971_, _05973_);
  not (_05998_, _05997_);
  and (_05999_, _05687_, _05936_);
  and (_06000_, _05999_, _05992_);
  and (_06001_, _06000_, _05973_);
  not (_06002_, _05944_);
  and (_06003_, _05999_, _06002_);
  and (_06004_, _06003_, _05973_);
  nor (_06005_, _06004_, _06001_);
  and (_06006_, _06005_, _05998_);
  and (_06007_, _05999_, _05765_);
  and (_06008_, _06007_, _05973_);
  not (_06009_, _06008_);
  and (_06010_, _06002_, _05688_);
  and (_06011_, _06010_, _05973_);
  and (_06012_, _05999_, _05894_);
  and (_06013_, _06012_, _05973_);
  nor (_06014_, _06013_, _06011_);
  and (_06015_, _06014_, _06009_);
  and (_06016_, _06015_, _06006_);
  and (_06017_, _06016_, _05996_);
  not (_06018_, \oc8051_golden_model_1.ACC [0]);
  and (_06019_, _06018_, \oc8051_golden_model_1.PC [0]);
  and (_06020_, \oc8051_golden_model_1.ACC [0], _05619_);
  or (_06021_, _06020_, _05985_);
  or (_06022_, _06021_, _06019_);
  and (_06023_, _06022_, _06017_);
  nand (_06024_, _06023_, _05988_);
  or (_06025_, _06017_, \oc8051_golden_model_1.PC [0]);
  nand (_06026_, _06025_, _06024_);
  and (_06027_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_06028_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_06029_, _06028_, _06027_);
  and (_06030_, _06029_, _05977_);
  nor (_06031_, _06029_, _05977_);
  nor (_06032_, _06031_, _06030_);
  nand (_06033_, _06032_, _05976_);
  and (_06034_, _05621_, _05586_);
  not (_06035_, _06034_);
  and (_06036_, _06035_, _05940_);
  nand (_06037_, _06036_, _05963_);
  nand (_06038_, _06037_, _06033_);
  nand (_06039_, _06038_, _05975_);
  and (_06040_, _05975_, _05963_);
  or (_06041_, _06040_, \oc8051_golden_model_1.PC [1]);
  nand (_06042_, _06041_, _06039_);
  nand (_06043_, _06042_, _05985_);
  not (_06044_, \oc8051_golden_model_1.ACC [1]);
  nor (_06045_, _06034_, _06044_);
  and (_06046_, _06034_, _06044_);
  nor (_06047_, _06046_, _06045_);
  and (_06048_, _06047_, _06020_);
  nor (_06049_, _06047_, _06020_);
  nor (_06050_, _06049_, _06048_);
  and (_06051_, _06050_, _05984_);
  not (_06052_, _06051_);
  and (_06053_, _06052_, _06017_);
  nand (_06054_, _06053_, _06043_);
  or (_06055_, _06017_, _05585_);
  nand (_06056_, _06055_, _06054_);
  or (_06057_, _06056_, _06026_);
  and (_06058_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_06059_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_06060_, _06059_, _06058_);
  and (_06061_, _06040_, _06017_);
  or (_06062_, _06061_, _06060_);
  nor (_06063_, _06030_, _06027_);
  and (_06064_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06065_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06066_, _06065_, _06064_);
  not (_06067_, _06066_);
  nor (_06068_, _06067_, _06063_);
  and (_06069_, _06067_, _06063_);
  nor (_06070_, _06069_, _06068_);
  or (_06071_, _06070_, _05940_);
  nor (_06072_, _05580_, _05590_);
  and (_06073_, _05580_, _05590_);
  nor (_06074_, _06073_, _06072_);
  not (_06075_, _06074_);
  and (_06076_, _06075_, _05940_);
  nand (_06077_, _06076_, _05963_);
  nand (_06078_, _06077_, _06071_);
  and (_06079_, _05985_, _05975_);
  and (_06080_, _06079_, _06078_);
  nor (_06081_, _06048_, _06045_);
  and (_06082_, _06074_, \oc8051_golden_model_1.ACC [2]);
  nor (_06083_, _06074_, \oc8051_golden_model_1.ACC [2]);
  nor (_06084_, _06083_, _06082_);
  not (_06085_, _06084_);
  nor (_06086_, _06085_, _06081_);
  and (_06087_, _06085_, _06081_);
  nor (_06088_, _06087_, _06086_);
  nor (_06089_, _06088_, _05985_);
  or (_06090_, _06089_, _06080_);
  nand (_06091_, _06090_, _06017_);
  and (_06092_, _06091_, _06062_);
  nor (_06093_, _05601_, _05585_);
  nor (_06094_, _06058_, \oc8051_golden_model_1.PC [3]);
  nor (_06095_, _06094_, _06093_);
  or (_06096_, _06095_, _06061_);
  nor (_06097_, _06086_, _06082_);
  not (_06098_, _05592_);
  nor (_06099_, _06072_, _05581_);
  nor (_06100_, _06099_, _06098_);
  nor (_06101_, _06100_, \oc8051_golden_model_1.ACC [3]);
  and (_06102_, _06100_, \oc8051_golden_model_1.ACC [3]);
  nor (_06103_, _06102_, _06101_);
  nor (_06104_, _06103_, _06097_);
  and (_06105_, _06103_, _06097_);
  nor (_06106_, _06105_, _06104_);
  nor (_06107_, _06106_, _05985_);
  nor (_06108_, _06068_, _06064_);
  and (_06109_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_06110_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_06111_, _06110_, _06109_);
  not (_06112_, _06111_);
  nor (_06113_, _06112_, _06108_);
  and (_06114_, _06112_, _06108_);
  nor (_06115_, _06114_, _06113_);
  or (_06116_, _06115_, _05940_);
  and (_06117_, _05940_, _06100_);
  nand (_06118_, _06117_, _05963_);
  nand (_06119_, _06118_, _06116_);
  and (_06120_, _06119_, _06079_);
  or (_06121_, _06120_, _06107_);
  nand (_06122_, _06121_, _06017_);
  nand (_06123_, _06122_, _06096_);
  or (_06124_, _06123_, _06092_);
  or (_06125_, _06124_, _06057_);
  or (_06126_, _06125_, _00401_);
  nand (_06127_, _06091_, _06062_);
  and (_06128_, _06122_, _06096_);
  or (_06129_, _06128_, _06127_);
  or (_06130_, _06129_, _06057_);
  or (_06131_, _06130_, _00237_);
  and (_06132_, _06131_, _06126_);
  and (_06133_, _06055_, _06054_);
  or (_06134_, _06133_, _06026_);
  or (_06135_, _06134_, _06129_);
  or (_06136_, _06135_, _00124_);
  and (_06137_, _06025_, _06024_);
  or (_06138_, _06133_, _06137_);
  or (_06139_, _06128_, _06092_);
  or (_06140_, _06139_, _06138_);
  or (_06141_, _06140_, _43185_);
  and (_06142_, _06141_, _06136_);
  and (_06143_, _06142_, _06132_);
  or (_06144_, _06123_, _06127_);
  or (_06145_, _06144_, _06057_);
  or (_06146_, _06145_, _00579_);
  or (_06147_, _06139_, _06057_);
  or (_06148_, _06147_, _00042_);
  and (_06149_, _06148_, _06146_);
  or (_06150_, _06056_, _06137_);
  or (_06151_, _06150_, _06144_);
  or (_06152_, _06151_, _00524_);
  or (_06153_, _06134_, _06124_);
  or (_06154_, _06153_, _00319_);
  and (_06155_, _06154_, _06152_);
  and (_06156_, _06155_, _06149_);
  and (_06157_, _06156_, _06143_);
  or (_06158_, _06150_, _06129_);
  or (_06159_, _06158_, _00196_);
  or (_06160_, _06138_, _06129_);
  or (_06161_, _06160_, _00083_);
  and (_06162_, _06161_, _06159_);
  or (_06163_, _06144_, _06138_);
  or (_06164_, _06163_, _00442_);
  or (_06165_, _06139_, _06134_);
  or (_06166_, _06165_, _43226_);
  and (_06167_, _06166_, _06164_);
  and (_06168_, _06167_, _06162_);
  or (_06169_, _06150_, _06124_);
  or (_06170_, _06169_, _00360_);
  or (_06171_, _06150_, _06139_);
  or (_06172_, _06171_, _43267_);
  and (_06173_, _06172_, _06170_);
  or (_06174_, _06144_, _06134_);
  or (_06175_, _06174_, _00483_);
  or (_06176_, _06138_, _06124_);
  or (_06177_, _06176_, _00278_);
  and (_06178_, _06177_, _06175_);
  and (_06179_, _06178_, _06173_);
  and (_06180_, _06179_, _06168_);
  nand (_06181_, _06180_, _06157_);
  or (_06182_, _06176_, _00298_);
  or (_06183_, _06135_, _00161_);
  and (_06184_, _06183_, _06182_);
  or (_06185_, _06145_, _00604_);
  or (_06186_, _06130_, _00257_);
  and (_06187_, _06186_, _06185_);
  and (_06188_, _06187_, _06184_);
  or (_06189_, _06153_, _00339_);
  or (_06190_, _06160_, _00103_);
  and (_06191_, _06190_, _06189_);
  or (_06192_, _06140_, _43205_);
  or (_06193_, _06165_, _43246_);
  and (_06194_, _06193_, _06192_);
  and (_06195_, _06194_, _06191_);
  and (_06196_, _06195_, _06188_);
  or (_06197_, _06174_, _00503_);
  or (_06198_, _06125_, _00421_);
  and (_06199_, _06198_, _06197_);
  or (_06200_, _06158_, _00216_);
  or (_06201_, _06171_, _00021_);
  and (_06202_, _06201_, _06200_);
  and (_06203_, _06202_, _06199_);
  or (_06204_, _06163_, _00462_);
  or (_06205_, _06169_, _00380_);
  and (_06206_, _06205_, _06204_);
  or (_06207_, _06151_, _00545_);
  or (_06208_, _06147_, _00062_);
  and (_06209_, _06208_, _06207_);
  and (_06210_, _06209_, _06206_);
  and (_06211_, _06210_, _06203_);
  and (_06212_, _06211_, _06196_);
  or (_06213_, _06212_, _06181_);
  nor (_06214_, _06213_, _05933_);
  and (_06215_, _06003_, _05970_);
  not (_06216_, _06215_);
  nor (_06217_, _06216_, _06181_);
  or (_06218_, _06158_, _00201_);
  or (_06219_, _06135_, _00129_);
  and (_06220_, _06219_, _06218_);
  or (_06221_, _06147_, _00047_);
  or (_06222_, _06171_, _00006_);
  and (_06223_, _06222_, _06221_);
  and (_06224_, _06223_, _06220_);
  or (_06225_, _06163_, _00447_);
  or (_06226_, _06153_, _00324_);
  and (_06227_, _06226_, _06225_);
  or (_06228_, _06125_, _00406_);
  or (_06229_, _06176_, _00283_);
  and (_06230_, _06229_, _06228_);
  and (_06231_, _06230_, _06227_);
  and (_06232_, _06231_, _06224_);
  or (_06233_, _06140_, _43190_);
  or (_06234_, _06165_, _43231_);
  and (_06235_, _06234_, _06233_);
  or (_06236_, _06130_, _00242_);
  or (_06237_, _06160_, _00088_);
  and (_06238_, _06237_, _06236_);
  and (_06239_, _06238_, _06235_);
  or (_06240_, _06145_, _00587_);
  or (_06241_, _06151_, _00529_);
  and (_06242_, _06241_, _06240_);
  or (_06243_, _06174_, _00488_);
  or (_06244_, _06169_, _00365_);
  and (_06245_, _06244_, _06243_);
  and (_06246_, _06245_, _06242_);
  and (_06247_, _06246_, _06239_);
  nand (_06248_, _06247_, _06232_);
  and (_06249_, _06248_, _06217_);
  not (_06250_, _06248_);
  not (_06251_, _05972_);
  and (_06252_, _05926_, _05802_);
  and (_06253_, _06252_, _05969_);
  and (_06254_, _06253_, _05971_);
  not (_06255_, _05934_);
  and (_06256_, _05969_, _06255_);
  and (_06257_, _06256_, _05971_);
  nor (_06258_, _06257_, _06254_);
  and (_06259_, _05971_, _05879_);
  not (_06260_, _06259_);
  and (_06261_, _06260_, _06258_);
  and (_06262_, _06261_, _06251_);
  nor (_06263_, _06262_, _06181_);
  and (_06264_, _06263_, _06250_);
  and (_06265_, _06252_, _05930_);
  and (_06266_, _06265_, _05938_);
  not (_06267_, _06266_);
  nor (_06268_, _06267_, _06213_);
  not (_06269_, _05945_);
  and (_06270_, _06265_, _06269_);
  not (_06271_, _06270_);
  nor (_06272_, _06271_, _06213_);
  nor (_06273_, _06271_, _06181_);
  not (_06274_, _06273_);
  not (_06275_, _05954_);
  and (_06276_, _06275_, _05931_);
  and (_06277_, _06265_, _06275_);
  not (_06278_, _06277_);
  nor (_06279_, _06278_, _06213_);
  not (_06280_, _05948_);
  and (_06281_, _06265_, _06280_);
  not (_06282_, _06281_);
  or (_06283_, _06282_, _06213_);
  nor (_06284_, _06282_, _06181_);
  and (_06285_, _05970_, _06280_);
  not (_06286_, _06285_);
  nor (_06287_, _06286_, _06181_);
  and (_06288_, _06287_, _06248_);
  not (_06289_, _05958_);
  and (_06290_, _06265_, _05993_);
  not (_06291_, _06290_);
  and (_06292_, _05993_, _05970_);
  not (_06293_, _06292_);
  not (_06294_, _06181_);
  nor (_06295_, _06174_, _00518_);
  nor (_06296_, _06125_, _00436_);
  nor (_06297_, _06296_, _06295_);
  nor (_06298_, _06160_, _00118_);
  nor (_06299_, _06140_, _43220_);
  nor (_06300_, _06299_, _06298_);
  and (_06301_, _06300_, _06297_);
  nor (_06302_, _06169_, _00395_);
  nor (_06303_, _06153_, _00354_);
  nor (_06304_, _06303_, _06302_);
  nor (_06305_, _06145_, _00619_);
  nor (_06306_, _06163_, _00477_);
  nor (_06307_, _06306_, _06305_);
  and (_06308_, _06307_, _06304_);
  and (_06309_, _06308_, _06301_);
  nor (_06310_, _06130_, _00272_);
  nor (_06311_, _06158_, _00231_);
  nor (_06312_, _06311_, _06310_);
  nor (_06313_, _06135_, _00190_);
  nor (_06314_, _06147_, _00077_);
  nor (_06315_, _06314_, _06313_);
  and (_06316_, _06315_, _06312_);
  nor (_06317_, _06171_, _00036_);
  nor (_06318_, _06165_, _43261_);
  nor (_06319_, _06318_, _06317_);
  nor (_06320_, _06151_, _00569_);
  nor (_06321_, _06176_, _00313_);
  nor (_06322_, _06321_, _06320_);
  and (_06323_, _06322_, _06319_);
  and (_06324_, _06323_, _06316_);
  and (_06325_, _06324_, _06309_);
  and (_06326_, _06325_, _06294_);
  and (_06327_, _06212_, _06181_);
  or (_06328_, _06327_, _06326_);
  and (_06329_, _06265_, _06003_);
  and (_06330_, _06265_, _05971_);
  nor (_06331_, _06330_, _06329_);
  not (_06332_, _06331_);
  and (_06333_, _06332_, _06328_);
  nor (_06334_, _05888_, _05952_);
  not (_06335_, _06334_);
  not (_06336_, _05952_);
  and (_06337_, _05882_, _06336_);
  and (_06338_, _05887_, _06255_);
  and (_06339_, _05887_, _05968_);
  or (_06340_, _06339_, _06338_);
  and (_06341_, _06340_, _06336_);
  nor (_06342_, _06341_, _06337_);
  and (_06343_, _06342_, _06335_);
  not (_06344_, _06343_);
  and (_06345_, _05970_, _06275_);
  not (_06346_, _06345_);
  and (_06347_, _05970_, _06269_);
  nor (_06348_, _06347_, _06276_);
  nand (_06349_, _06348_, _06346_);
  nor (_06350_, _06349_, _06344_);
  or (_06351_, _06350_, _06212_);
  and (_06352_, _06328_, _06281_);
  not (_06353_, \oc8051_golden_model_1.SP [3]);
  and (_06354_, _06280_, _05931_);
  and (_06355_, _06354_, _06353_);
  not (_06356_, _06212_);
  not (_06357_, _05959_);
  and (_06358_, _05970_, _06357_);
  or (_06359_, _06358_, _06285_);
  nand (_06360_, _06359_, _06356_);
  nor (_06361_, _06354_, _06281_);
  not (_06362_, \oc8051_golden_model_1.PSW [3]);
  or (_06363_, _06359_, _06362_);
  and (_06364_, _06363_, _06361_);
  or (_06365_, _06364_, _06345_);
  and (_06366_, _06365_, _06360_);
  or (_06367_, _06366_, _06355_);
  and (_06368_, _06269_, _05931_);
  nor (_06369_, _06368_, _06270_);
  and (_06370_, _06336_, _05931_);
  and (_06371_, _06265_, _06336_);
  nor (_06372_, _06371_, _06370_);
  and (_06373_, _06372_, _06369_);
  and (_06374_, _06373_, _06278_);
  and (_06375_, _06374_, _06367_);
  or (_06376_, _06375_, _06352_);
  and (_06377_, _06376_, _06351_);
  not (_06378_, _06328_);
  nor (_06379_, _06374_, _06378_);
  and (_06380_, _05970_, _05938_);
  nand (_06381_, _06348_, _06343_);
  and (_06382_, _06381_, _06212_);
  or (_06383_, _06382_, _06380_);
  or (_06384_, _06383_, _06379_);
  or (_06385_, _06384_, _06377_);
  not (_06386_, _06380_);
  nor (_06387_, _06386_, _06212_);
  nor (_06388_, _06387_, _06266_);
  nand (_06389_, _06388_, _06385_);
  and (_06390_, _06328_, _06266_);
  nor (_06391_, _06390_, _05972_);
  nand (_06392_, _06391_, _06389_);
  and (_06393_, _06265_, _05766_);
  nor (_06394_, _06393_, _05932_);
  and (_06395_, _05938_, _05931_);
  not (_06396_, _06395_);
  not (_06397_, _05935_);
  and (_06398_, _06000_, _06397_);
  nor (_06399_, _06398_, _06215_);
  and (_06400_, _06399_, _06396_);
  and (_06401_, _05887_, _06252_);
  and (_06402_, _05882_, _06252_);
  or (_06403_, _06402_, _06401_);
  and (_06404_, _06403_, _06269_);
  not (_06405_, _06404_);
  and (_06406_, _06405_, _06400_);
  and (_06407_, _05882_, _06255_);
  nand (_06408_, _06407_, _06269_);
  and (_06409_, _05887_, _05928_);
  nand (_06410_, _06409_, _06269_);
  and (_06411_, _06410_, _06408_);
  and (_06412_, _06411_, _06286_);
  and (_06413_, _06338_, _06269_);
  and (_06414_, _05882_, _05927_);
  and (_06415_, _06414_, _06269_);
  nor (_06416_, _06415_, _06413_);
  and (_06417_, _06416_, _06412_);
  and (_06418_, _05969_, _05928_);
  and (_06419_, _06418_, _06269_);
  nor (_06420_, _06419_, _06347_);
  and (_06421_, _06253_, _06269_);
  and (_06422_, _06256_, _06269_);
  or (_06423_, _06422_, _06421_);
  not (_06424_, _06423_);
  and (_06425_, _06424_, _06420_);
  and (_06426_, _06012_, _06397_);
  and (_06427_, _06339_, _06269_);
  nor (_06428_, _06427_, _06426_);
  and (_06429_, _06428_, _06425_);
  and (_06430_, _06429_, _06417_);
  and (_06431_, _06430_, _06406_);
  and (_06432_, _06265_, _05895_);
  not (_06433_, _06432_);
  and (_06434_, _05993_, _05931_);
  not (_06435_, _06434_);
  and (_06436_, _06010_, _05931_);
  and (_06437_, _06007_, _06397_);
  nor (_06438_, _06437_, _06436_);
  and (_06439_, _06438_, _06435_);
  and (_06440_, _06439_, _06433_);
  and (_06441_, _06440_, _06431_);
  and (_06442_, _06441_, _06394_);
  nor (_06443_, _06442_, _05619_);
  and (_06444_, _06442_, _05619_);
  nor (_06445_, _06444_, _06443_);
  not (_06446_, _06445_);
  nor (_06447_, _06444_, _05585_);
  and (_06448_, _06444_, _05585_);
  nor (_06449_, _06448_, _06447_);
  and (_06450_, _06449_, _06446_);
  not (_06451_, _06060_);
  nor (_06452_, _06442_, _06451_);
  and (_06453_, _06394_, _06074_);
  and (_06454_, _06453_, _06441_);
  nor (_06455_, _06454_, _06452_);
  not (_06456_, _06095_);
  nor (_06457_, _06442_, _06456_);
  not (_06458_, _06100_);
  and (_06459_, _06442_, _06458_);
  nor (_06460_, _06459_, _06457_);
  nor (_06461_, _06460_, _06455_);
  and (_06462_, _06461_, _06450_);
  and (_06463_, _06462_, _04698_);
  not (_06464_, _06463_);
  nor (_06465_, _06449_, _06445_);
  and (_06466_, _06461_, _06465_);
  and (_06467_, _06466_, _04707_);
  and (_06468_, _06449_, _06445_);
  and (_06469_, _06468_, _06461_);
  and (_06470_, _06469_, _04700_);
  nor (_06471_, _06470_, _06467_);
  not (_06472_, _06455_);
  nor (_06473_, _06460_, _06472_);
  and (_06474_, _06450_, _06473_);
  and (_06475_, _06474_, _04687_);
  nor (_06476_, _06449_, _06446_);
  and (_06477_, _06476_, _06461_);
  and (_06478_, _06477_, _04685_);
  nor (_06479_, _06478_, _06475_);
  and (_06480_, _06479_, _06471_);
  and (_06481_, _06468_, _06473_);
  and (_06482_, _06481_, _04671_);
  and (_06483_, _06465_, _06473_);
  and (_06484_, _06483_, _04669_);
  nor (_06485_, _06484_, _06482_);
  and (_06486_, _06460_, _06472_);
  and (_06487_, _06486_, _06450_);
  and (_06488_, _06487_, _04702_);
  and (_06489_, _06476_, _06473_);
  and (_06490_, _06489_, _04674_);
  nor (_06491_, _06490_, _06488_);
  and (_06492_, _06491_, _06485_);
  and (_06493_, _06492_, _06480_);
  and (_06494_, _06486_, _06465_);
  and (_06495_, _06494_, _04709_);
  and (_06496_, _06468_, _06486_);
  and (_06497_, _06496_, _04690_);
  nor (_06498_, _06497_, _06495_);
  and (_06499_, _06460_, _06455_);
  and (_06500_, _06499_, _06450_);
  and (_06501_, _06500_, _04696_);
  and (_06502_, _06476_, _06486_);
  and (_06503_, _06502_, _04692_);
  nor (_06504_, _06503_, _06501_);
  and (_06505_, _06504_, _06498_);
  and (_06506_, _06499_, _06476_);
  and (_06507_, _06506_, _04680_);
  not (_06508_, _06507_);
  and (_06509_, _06499_, _06468_);
  and (_06510_, _06509_, _04676_);
  and (_06511_, _06499_, _06465_);
  and (_06512_, _06511_, _04682_);
  nor (_06513_, _06512_, _06510_);
  and (_06514_, _06513_, _06508_);
  and (_06515_, _06514_, _06505_);
  and (_06516_, _06515_, _06493_);
  and (_06517_, _06516_, _06464_);
  nor (_06518_, _06517_, _06251_);
  nor (_06519_, _06518_, _06332_);
  and (_06520_, _06519_, _06392_);
  or (_06521_, _06520_, _06333_);
  and (_06522_, _06010_, _05970_);
  not (_06523_, _06522_);
  and (_06524_, _06265_, _06000_);
  nor (_06525_, _06524_, _06398_);
  and (_06526_, _06000_, _05970_);
  not (_06527_, _06526_);
  and (_06528_, _06527_, _06525_);
  and (_06529_, _06528_, _06523_);
  and (_06530_, _06012_, _05970_);
  not (_06531_, _06530_);
  and (_06532_, _06265_, _06012_);
  nor (_06533_, _06532_, _06426_);
  and (_06534_, _06533_, _06531_);
  and (_06535_, _06265_, _06007_);
  nor (_06536_, _06535_, _06437_);
  and (_06537_, _06007_, _05970_);
  not (_06538_, _06537_);
  and (_06539_, _06538_, _06536_);
  and (_06540_, _06539_, _06534_);
  and (_06541_, _06540_, _06529_);
  nand (_06542_, _06541_, _06521_);
  and (_06543_, _06265_, _06010_);
  nor (_06544_, _06541_, _06356_);
  nor (_06545_, _06544_, _06543_);
  and (_06546_, _06545_, _06542_);
  and (_06547_, _06543_, \oc8051_golden_model_1.SP [3]);
  or (_06548_, _06547_, _06436_);
  nor (_06549_, _06548_, _06546_);
  and (_06550_, _06436_, _06328_);
  or (_06551_, _06550_, _06549_);
  and (_06552_, _06551_, _06293_);
  and (_06553_, _06292_, _06212_);
  or (_06554_, _06553_, _06552_);
  nand (_06555_, _06554_, _06291_);
  and (_06556_, _06290_, _06353_);
  nor (_06557_, _06556_, _06434_);
  and (_06558_, _06557_, _06555_);
  and (_06559_, _05970_, _05895_);
  nor (_06560_, _06328_, _06435_);
  or (_06561_, _06560_, _06559_);
  nor (_06562_, _06561_, _06558_);
  and (_06563_, _06559_, _06212_);
  or (_06564_, _06563_, _06562_);
  nand (_06565_, _06564_, _05933_);
  and (_06566_, _05766_, _05970_);
  and (_06567_, _06328_, _05932_);
  nor (_06568_, _06567_, _06566_);
  nand (_06569_, _06568_, _06565_);
  not (_06570_, _06566_);
  nor (_06571_, _06570_, _06212_);
  not (_06572_, _06571_);
  and (_06573_, _06572_, _06569_);
  nor (_06574_, _06145_, _00614_);
  nor (_06575_, _06153_, _00349_);
  nor (_06576_, _06575_, _06574_);
  nor (_06577_, _06169_, _00390_);
  nor (_06578_, _06147_, _00072_);
  nor (_06579_, _06578_, _06577_);
  and (_06580_, _06579_, _06576_);
  nor (_06581_, _06130_, _00267_);
  nor (_06582_, _06160_, _00113_);
  nor (_06583_, _06582_, _06581_);
  nor (_06584_, _06174_, _00513_);
  nor (_06585_, _06163_, _00472_);
  nor (_06586_, _06585_, _06584_);
  and (_06587_, _06586_, _06583_);
  and (_06588_, _06587_, _06580_);
  nor (_06589_, _06135_, _00183_);
  nor (_06590_, _06171_, _00031_);
  nor (_06591_, _06590_, _06589_);
  nor (_06592_, _06140_, _43215_);
  nor (_06593_, _06165_, _43256_);
  nor (_06594_, _06593_, _06592_);
  and (_06595_, _06594_, _06591_);
  nor (_06596_, _06151_, _00561_);
  nor (_06597_, _06158_, _00226_);
  nor (_06598_, _06597_, _06596_);
  nor (_06599_, _06125_, _00431_);
  nor (_06600_, _06176_, _00308_);
  nor (_06601_, _06600_, _06599_);
  and (_06602_, _06601_, _06598_);
  and (_06603_, _06602_, _06595_);
  and (_06604_, _06603_, _06588_);
  nor (_06605_, _06604_, _06181_);
  nor (_06606_, _06266_, _05932_);
  and (_06607_, _06606_, _06435_);
  and (_06608_, _06607_, _06331_);
  nor (_06609_, _06436_, _06281_);
  and (_06610_, _06609_, _06374_);
  and (_06611_, _06610_, _06608_);
  not (_06612_, _06611_);
  and (_06613_, _06612_, _06605_);
  not (_06614_, _06613_);
  nor (_06615_, _06147_, _00057_);
  nor (_06616_, _06171_, _00016_);
  nor (_06617_, _06616_, _06615_);
  nor (_06618_, _06135_, _00150_);
  nor (_06619_, _06165_, _43241_);
  nor (_06620_, _06619_, _06618_);
  and (_06621_, _06620_, _06617_);
  nor (_06622_, _06163_, _00457_);
  nor (_06623_, _06169_, _00375_);
  nor (_06624_, _06623_, _06622_);
  nor (_06625_, _06145_, _00599_);
  nor (_06626_, _06174_, _00498_);
  nor (_06627_, _06626_, _06625_);
  and (_06628_, _06627_, _06624_);
  and (_06629_, _06628_, _06621_);
  nor (_06630_, _06153_, _00334_);
  nor (_06632_, _06160_, _00098_);
  nor (_06633_, _06632_, _06630_);
  nor (_06634_, _06125_, _00416_);
  nor (_06635_, _06140_, _43200_);
  nor (_06636_, _06635_, _06634_);
  and (_06637_, _06636_, _06633_);
  nor (_06638_, _06176_, _00293_);
  nor (_06639_, _06158_, _00211_);
  nor (_06640_, _06639_, _06638_);
  nor (_06641_, _06151_, _00539_);
  nor (_06642_, _06130_, _00252_);
  nor (_06643_, _06642_, _06641_);
  and (_06644_, _06643_, _06640_);
  and (_06645_, _06644_, _06637_);
  and (_06646_, _06645_, _06629_);
  not (_06647_, _06646_);
  nor (_06648_, _06380_, _06359_);
  nand (_06649_, _06648_, _06343_);
  or (_06650_, _06649_, _06349_);
  nor (_06651_, _06566_, _06559_);
  and (_06652_, _06651_, _06293_);
  nand (_06653_, _06652_, _06541_);
  or (_06654_, _06653_, _06650_);
  and (_06655_, _06654_, _06647_);
  not (_06656_, _06655_);
  and (_06657_, _06462_, _04623_);
  not (_06658_, _06657_);
  and (_06659_, _06500_, _04639_);
  and (_06660_, _06502_, _04637_);
  nor (_06661_, _06660_, _06659_);
  and (_06662_, _06496_, _04632_);
  and (_06663_, _06494_, _04634_);
  nor (_06664_, _06663_, _06662_);
  and (_06665_, _06664_, _06661_);
  and (_06666_, _06506_, _04627_);
  not (_06667_, _06666_);
  and (_06668_, _06511_, _04630_);
  and (_06669_, _06509_, _04625_);
  nor (_06670_, _06669_, _06668_);
  and (_06671_, _06670_, _06667_);
  and (_06672_, _06671_, _06665_);
  and (_06673_, _06466_, _04645_);
  and (_06674_, _06469_, _04647_);
  nor (_06675_, _06674_, _06673_);
  and (_06676_, _06474_, _04650_);
  and (_06677_, _06477_, _04652_);
  nor (_06678_, _06677_, _06676_);
  and (_06679_, _06678_, _06675_);
  and (_06680_, _06483_, _04658_);
  and (_06681_, _06481_, _04656_);
  nor (_06682_, _06681_, _06680_);
  and (_06683_, _06489_, _04661_);
  and (_06684_, _06487_, _04663_);
  nor (_06685_, _06684_, _06683_);
  and (_06686_, _06685_, _06682_);
  and (_06687_, _06686_, _06679_);
  and (_06688_, _06687_, _06672_);
  and (_06689_, _06688_, _06658_);
  nor (_06690_, _06689_, _06251_);
  or (_06691_, _05993_, _06010_);
  or (_06692_, _06007_, _06000_);
  or (_06693_, _06692_, _06691_);
  and (_06694_, _06693_, _05926_);
  or (_06695_, _06012_, _05895_);
  nor (_06696_, _05937_, _05892_);
  or (_06697_, _06696_, _05766_);
  or (_06698_, _06697_, _06695_);
  or (_06699_, _06698_, _06694_);
  and (_06700_, _06699_, _05887_);
  not (_06701_, _06700_);
  and (_06702_, _05887_, _05926_);
  not (_06703_, _06702_);
  and (_06704_, _05959_, _05948_);
  nor (_06705_, _06704_, _06703_);
  not (_06706_, _06705_);
  and (_06707_, _06290_, \oc8051_golden_model_1.SP [2]);
  and (_06708_, _06543_, \oc8051_golden_model_1.SP [2]);
  nor (_06709_, _06708_, _06707_);
  and (_06710_, _06709_, _06706_);
  and (_06711_, _06702_, _06275_);
  and (_06712_, _06702_, _05971_);
  nor (_06713_, _06712_, _06711_);
  and (_06714_, _05887_, _05927_);
  and (_06715_, _06714_, _05993_);
  and (_06716_, _06714_, _06007_);
  nor (_06717_, _06716_, _06715_);
  and (_06718_, _06717_, _06713_);
  and (_06719_, _06714_, _06275_);
  and (_06720_, _06714_, _06280_);
  nor (_06721_, _06720_, _06719_);
  not (_06722_, _06714_);
  nor (_06723_, _06000_, _05971_);
  nor (_06724_, _06723_, _06722_);
  not (_06725_, _06724_);
  and (_06726_, _06725_, _06721_);
  and (_06727_, _06354_, \oc8051_golden_model_1.SP [2]);
  nor (_06728_, _06010_, _06357_);
  nor (_06729_, _06728_, _06722_);
  nor (_06730_, _06729_, _06727_);
  and (_06731_, _06730_, _06726_);
  and (_06732_, _06731_, _06718_);
  and (_06733_, _06732_, _06710_);
  and (_06734_, _06733_, _06701_);
  not (_06735_, _06734_);
  nor (_06736_, _06735_, _06690_);
  and (_06737_, _06736_, _06656_);
  and (_06738_, _06737_, _06614_);
  not (_06739_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_06740_, _06566_, _06248_);
  not (_06741_, _06740_);
  and (_06742_, _06380_, _06248_);
  nor (_06743_, _06372_, _06213_);
  and (_06744_, _06347_, _06248_);
  nand (_06745_, _06345_, _06248_);
  and (_06746_, _06359_, _06248_);
  nor (_06747_, _05883_, _06253_);
  and (_06748_, _06747_, _05888_);
  nor (_06749_, _06748_, _05948_);
  not (_06750_, _06749_);
  nor (_06751_, _06409_, _05970_);
  and (_06752_, _06751_, _06747_);
  nor (_06753_, _06752_, _05959_);
  not (_06754_, _06753_);
  and (_06755_, _06401_, _06357_);
  not (_06756_, _06755_);
  not (_06757_, _05957_);
  and (_06758_, _06253_, _06757_);
  nor (_06759_, _06758_, _06285_);
  and (_06760_, _06759_, _06756_);
  and (_06761_, _06760_, _06754_);
  and (_06762_, _06761_, _06750_);
  or (_06763_, _06762_, _06746_);
  nand (_06764_, _06763_, _06282_);
  nand (_06765_, _06283_, _06764_);
  not (_06766_, \oc8051_golden_model_1.SP [0]);
  and (_06767_, _06354_, _06766_);
  nor (_06768_, _06767_, _06345_);
  and (_06769_, _06253_, _06275_);
  nor (_06770_, _05883_, _05890_);
  nor (_06771_, _06770_, _05954_);
  nor (_06772_, _06771_, _06769_);
  and (_06773_, _06772_, _06768_);
  nand (_06774_, _06773_, _06765_);
  nand (_06775_, _06774_, _06745_);
  and (_06776_, _06775_, _06278_);
  or (_06777_, _06279_, _06776_);
  not (_06778_, _06276_);
  nor (_06779_, _06778_, _06248_);
  not (_06780_, _06401_);
  and (_06781_, _06751_, _06780_);
  and (_06782_, _06781_, _06747_);
  nor (_06783_, _06782_, _05945_);
  nor (_06784_, _06783_, _06779_);
  and (_06785_, _06784_, _06777_);
  or (_06786_, _06785_, _06744_);
  nand (_06787_, _06786_, _06369_);
  nor (_06788_, _06369_, _06213_);
  nor (_06789_, _06788_, _06344_);
  nand (_06790_, _06789_, _06787_);
  nor (_06791_, _06343_, _06248_);
  and (_06792_, _06253_, _06336_);
  not (_06793_, _06792_);
  and (_06794_, _06793_, _06372_);
  not (_06795_, _06794_);
  nor (_06796_, _06795_, _06791_);
  and (_06797_, _06796_, _06790_);
  or (_06798_, _06797_, _06743_);
  nor (_06799_, _06781_, _05939_);
  not (_06800_, _06799_);
  and (_06801_, _05882_, _05928_);
  and (_06802_, _06801_, _05938_);
  not (_06803_, _06802_);
  and (_06804_, _06402_, _05938_);
  and (_06805_, _06253_, _05938_);
  nor (_06806_, _06805_, _06804_);
  and (_06807_, _06806_, _06803_);
  and (_06808_, _06807_, _06800_);
  and (_06809_, _06808_, _06798_);
  or (_06810_, _06809_, _06742_);
  and (_06811_, _06810_, _06267_);
  or (_06812_, _06811_, _06268_);
  and (_06813_, _06801_, _05971_);
  nor (_06814_, _06402_, _06409_);
  nor (_06815_, _06253_, _06401_);
  nand (_06816_, _06815_, _06814_);
  and (_06817_, _06816_, _05971_);
  nor (_06818_, _06817_, _06813_);
  and (_06819_, _06818_, _06812_);
  and (_06820_, _06483_, _04530_);
  and (_06821_, _06496_, _04548_);
  nor (_06822_, _06821_, _06820_);
  and (_06823_, _06511_, _04572_);
  and (_06824_, _06494_, _04543_);
  nor (_06825_, _06824_, _06823_);
  and (_06826_, _06825_, _06822_);
  and (_06827_, _06487_, _04558_);
  and (_06828_, _06506_, _04570_);
  nor (_06829_, _06828_, _06827_);
  and (_06830_, _06481_, _04532_);
  and (_06831_, _06502_, _04565_);
  nor (_06832_, _06831_, _06830_);
  and (_06833_, _06832_, _06829_);
  and (_06834_, _06833_, _06826_);
  and (_06835_, _06462_, _04554_);
  and (_06836_, _06474_, _04546_);
  nor (_06837_, _06836_, _06835_);
  and (_06838_, _06469_, _04556_);
  and (_06839_, _06477_, _04563_);
  nor (_06840_, _06839_, _06838_);
  and (_06841_, _06840_, _06837_);
  and (_06842_, _06489_, _04535_);
  and (_06843_, _06509_, _04537_);
  nor (_06844_, _06843_, _06842_);
  and (_06845_, _06466_, _04541_);
  and (_06846_, _06500_, _04552_);
  nor (_06847_, _06846_, _06845_);
  and (_06848_, _06847_, _06844_);
  and (_06849_, _06848_, _06841_);
  and (_06850_, _06849_, _06834_);
  and (_06851_, _06850_, _05972_);
  nor (_06852_, _06851_, _06330_);
  and (_06853_, _06852_, _06819_);
  not (_06854_, _06330_);
  nor (_06855_, _06854_, _06213_);
  or (_06856_, _06855_, _06853_);
  and (_06857_, _06253_, _06003_);
  nor (_06858_, _06857_, _06329_);
  and (_06859_, _06858_, _06856_);
  not (_06860_, _06329_);
  nor (_06861_, _06860_, _06213_);
  or (_06862_, _06861_, _06859_);
  and (_06863_, _06401_, _06000_);
  and (_06864_, _06409_, _06000_);
  nor (_06865_, _06864_, _06863_);
  and (_06866_, _06801_, _06000_);
  not (_06867_, _06866_);
  and (_06868_, _06253_, _06000_);
  and (_06869_, _06402_, _06000_);
  nor (_06870_, _06869_, _06868_);
  and (_06871_, _06870_, _06867_);
  and (_06872_, _06871_, _06865_);
  and (_06873_, _06872_, _06862_);
  nor (_06874_, _06528_, _06248_);
  not (_06875_, _06012_);
  nor (_06876_, _06748_, _06875_);
  nor (_06877_, _06876_, _06874_);
  and (_06878_, _06877_, _06873_);
  nor (_06879_, _06540_, _06248_);
  and (_06880_, _05890_, _06007_);
  and (_06881_, _06801_, _06007_);
  and (_06882_, _06402_, _06007_);
  and (_06883_, _06253_, _06007_);
  or (_06884_, _06883_, _06882_);
  or (_06885_, _06884_, _06881_);
  nor (_06886_, _06885_, _06880_);
  and (_06887_, _06402_, _06010_);
  not (_06888_, _06887_);
  not (_06889_, _06010_);
  nor (_06890_, _06781_, _06889_);
  and (_06891_, _06801_, _06010_);
  and (_06892_, _06253_, _06010_);
  or (_06893_, _06892_, _06891_);
  nor (_06894_, _06893_, _06890_);
  and (_06895_, _06894_, _06888_);
  and (_06896_, _06895_, _06886_);
  not (_06897_, _06896_);
  nor (_06898_, _06897_, _06879_);
  and (_06899_, _06898_, _06878_);
  and (_06900_, _06522_, _06248_);
  nor (_06901_, _06900_, _06899_);
  and (_06902_, _06543_, _06766_);
  nor (_06903_, _06902_, _06901_);
  not (_06904_, _05993_);
  nor (_06905_, _06782_, _06904_);
  and (_06906_, _06436_, _06213_);
  nor (_06907_, _06906_, _06905_);
  and (_06908_, _06907_, _06903_);
  and (_06909_, _06292_, _06248_);
  nor (_06910_, _06909_, _06908_);
  and (_06911_, _06290_, _06766_);
  nor (_06912_, _06911_, _06910_);
  not (_06913_, _05895_);
  nor (_06914_, _06782_, _06913_);
  and (_06915_, _06434_, _06213_);
  nor (_06916_, _06915_, _06914_);
  and (_06917_, _06916_, _06912_);
  and (_06918_, _06559_, _06248_);
  or (_06919_, _06918_, _06917_);
  and (_06920_, _06919_, _05933_);
  or (_06921_, _06920_, _06214_);
  not (_06922_, _05891_);
  and (_06923_, _06253_, _05766_);
  not (_06924_, _06923_);
  nor (_06925_, _05884_, _06566_);
  and (_06926_, _06925_, _06924_);
  and (_06927_, _06926_, _06922_);
  nand (_06928_, _06927_, _06921_);
  nand (_06929_, _06928_, _06741_);
  or (_06930_, _06929_, _06739_);
  nor (_06931_, _06125_, _00426_);
  nor (_06932_, _06165_, _43251_);
  nor (_06933_, _06932_, _06931_);
  nor (_06934_, _06145_, _00609_);
  nor (_06935_, _06135_, _00172_);
  nor (_06936_, _06935_, _06934_);
  and (_06937_, _06936_, _06933_);
  nor (_06938_, _06169_, _00385_);
  nor (_06939_, _06153_, _00344_);
  nor (_06940_, _06939_, _06938_);
  nor (_06941_, _06151_, _00553_);
  nor (_06942_, _06147_, _00067_);
  nor (_06943_, _06942_, _06941_);
  and (_06944_, _06943_, _06940_);
  and (_06945_, _06944_, _06937_);
  nor (_06946_, _06130_, _00262_);
  nor (_06947_, _06158_, _00221_);
  nor (_06948_, _06947_, _06946_);
  nor (_06949_, _06160_, _00108_);
  nor (_06950_, _06140_, _43210_);
  nor (_06951_, _06950_, _06949_);
  and (_06952_, _06951_, _06948_);
  nor (_06953_, _06176_, _00303_);
  nor (_06954_, _06171_, _00026_);
  nor (_06955_, _06954_, _06953_);
  nor (_06956_, _06174_, _00508_);
  nor (_06957_, _06163_, _00467_);
  nor (_06958_, _06957_, _06956_);
  and (_06959_, _06958_, _06955_);
  and (_06960_, _06959_, _06952_);
  and (_06961_, _06960_, _06945_);
  nor (_06962_, _06961_, _06181_);
  and (_06963_, _06962_, _06612_);
  not (_06964_, _06963_);
  nor (_06965_, _06130_, _00247_);
  nor (_06966_, _06147_, _00052_);
  nor (_06967_, _06966_, _06965_);
  nor (_06968_, _06151_, _00534_);
  nor (_06969_, _06153_, _00329_);
  nor (_06970_, _06969_, _06968_);
  and (_06971_, _06970_, _06967_);
  nor (_06972_, _06158_, _00206_);
  nor (_06973_, _06135_, _00139_);
  nor (_06974_, _06973_, _06972_);
  nor (_06975_, _06160_, _00093_);
  nor (_06976_, _06140_, _43195_);
  nor (_06977_, _06976_, _06975_);
  and (_06978_, _06977_, _06974_);
  and (_06979_, _06978_, _06971_);
  nor (_06980_, _06163_, _00452_);
  nor (_06981_, _06125_, _00411_);
  nor (_06982_, _06981_, _06980_);
  nor (_06983_, _06145_, _00594_);
  nor (_06984_, _06174_, _00493_);
  nor (_06985_, _06984_, _06983_);
  and (_06986_, _06985_, _06982_);
  nor (_06987_, _06171_, _00011_);
  nor (_06988_, _06165_, _43236_);
  nor (_06989_, _06988_, _06987_);
  nor (_06990_, _06169_, _00370_);
  nor (_06991_, _06176_, _00288_);
  nor (_06992_, _06991_, _06990_);
  and (_06993_, _06992_, _06989_);
  and (_06994_, _06993_, _06986_);
  and (_06995_, _06994_, _06979_);
  not (_06996_, _06995_);
  and (_06997_, _06996_, _06654_);
  not (_06998_, _06997_);
  and (_06999_, _06462_, _04600_);
  not (_07000_, _06999_);
  and (_07001_, _06494_, _04594_);
  and (_07002_, _06496_, _04587_);
  nor (_07003_, _07002_, _07001_);
  and (_07004_, _06500_, _04598_);
  and (_07005_, _06502_, _04589_);
  nor (_07006_, _07005_, _07004_);
  and (_07007_, _07006_, _07003_);
  and (_07008_, _06506_, _04617_);
  not (_07009_, _07008_);
  and (_07010_, _06509_, _04583_);
  and (_07011_, _06511_, _04619_);
  nor (_07012_, _07011_, _07010_);
  and (_07013_, _07012_, _07009_);
  and (_07014_, _07013_, _07007_);
  and (_07015_, _06469_, _04602_);
  and (_07016_, _06466_, _04609_);
  nor (_07017_, _07016_, _07015_);
  and (_07018_, _06477_, _04611_);
  and (_07019_, _06474_, _04592_);
  nor (_07020_, _07019_, _07018_);
  and (_07021_, _07020_, _07017_);
  and (_07022_, _06481_, _04578_);
  and (_07023_, _06483_, _04576_);
  nor (_07024_, _07023_, _07022_);
  and (_07025_, _06489_, _04581_);
  and (_07026_, _06487_, _04604_);
  nor (_07027_, _07026_, _07025_);
  and (_07028_, _07027_, _07024_);
  and (_07029_, _07028_, _07021_);
  and (_07030_, _07029_, _07014_);
  and (_07031_, _07030_, _07000_);
  nor (_07032_, _07031_, _06251_);
  and (_07033_, _06354_, \oc8051_golden_model_1.SP [1]);
  nand (_07034_, _05882_, _05926_);
  nor (_07035_, _07034_, _06904_);
  nor (_07036_, _07035_, _07033_);
  and (_07037_, _06543_, \oc8051_golden_model_1.SP [1]);
  or (_07038_, _06696_, _06275_);
  and (_07039_, _07038_, _06702_);
  nor (_07040_, _07039_, _07037_);
  and (_07041_, _07040_, _07036_);
  not (_07042_, _05766_);
  nor (_07043_, _07034_, _07042_);
  nor (_07044_, _07034_, _05948_);
  nor (_07045_, _07044_, _07043_);
  nor (_07046_, _07034_, _05954_);
  or (_07047_, _07046_, _06712_);
  nor (_07048_, _07047_, _06705_);
  and (_07049_, _07048_, _07045_);
  and (_07050_, _07049_, _07041_);
  nor (_07051_, _06696_, _06357_);
  nand (_07052_, _05727_, _05688_);
  and (_07053_, _07052_, _06723_);
  and (_07054_, _07053_, _07051_);
  or (_07055_, _07054_, _07034_);
  or (_07056_, _05766_, _06012_);
  nor (_07057_, _07056_, _06693_);
  or (_07058_, _07057_, _06703_);
  not (_07059_, _06007_);
  nor (_07060_, _07034_, _07059_);
  not (_07061_, _07060_);
  nand (_07062_, _06702_, _05895_);
  and (_07063_, _07062_, _07061_);
  and (_07064_, _06290_, \oc8051_golden_model_1.SP [1]);
  and (_07065_, _06402_, _06012_);
  and (_07066_, _06407_, _06012_);
  or (_07067_, _07066_, _07065_);
  nor (_07068_, _07067_, _07064_);
  and (_07069_, _07068_, _07063_);
  and (_07070_, _07069_, _07058_);
  and (_07071_, _07070_, _07055_);
  and (_07072_, _07071_, _07050_);
  not (_07073_, _07072_);
  nor (_07074_, _07073_, _07032_);
  and (_07075_, _07074_, _06998_);
  and (_07076_, _07075_, _06964_);
  not (_07077_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_07078_, _06928_, _06741_);
  or (_07079_, _07078_, _07077_);
  and (_07080_, _07079_, _07076_);
  nand (_07081_, _07080_, _06930_);
  not (_07082_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_07083_, _07078_, _07082_);
  not (_07084_, _07076_);
  not (_07085_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_07086_, _06929_, _07085_);
  and (_07087_, _07086_, _07084_);
  nand (_07088_, _07087_, _07083_);
  nand (_07089_, _07088_, _07081_);
  nand (_07090_, _07089_, _06738_);
  not (_07091_, _06738_);
  not (_07092_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_07093_, _07078_, _07092_);
  not (_07094_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_07095_, _06929_, _07094_);
  and (_07096_, _07095_, _07084_);
  nand (_07097_, _07096_, _07093_);
  not (_07098_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_07099_, _06929_, _07098_);
  not (_07100_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_07101_, _07078_, _07100_);
  and (_07102_, _07101_, _07076_);
  nand (_07103_, _07102_, _07099_);
  nand (_07104_, _07103_, _07097_);
  nand (_07105_, _07104_, _07091_);
  nand (_07106_, _07105_, _07090_);
  nand (_07107_, _07106_, _06573_);
  not (_07108_, _06573_);
  not (_07109_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_07110_, _07078_, _07109_);
  not (_07111_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_07112_, _06929_, _07111_);
  and (_07113_, _07112_, _07084_);
  nand (_07114_, _07113_, _07110_);
  nand (_07115_, _07078_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand (_07116_, _06929_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_07117_, _07116_, _07076_);
  nand (_07118_, _07117_, _07115_);
  nand (_07119_, _07118_, _07114_);
  nand (_07120_, _07119_, _06738_);
  not (_07121_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_07122_, _07078_, _07121_);
  not (_07123_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_07124_, _06929_, _07123_);
  and (_07125_, _07124_, _07084_);
  nand (_07126_, _07125_, _07122_);
  nand (_07127_, _07078_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand (_07128_, _06929_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_07129_, _07128_, _07076_);
  nand (_07130_, _07129_, _07127_);
  nand (_07131_, _07130_, _07126_);
  nand (_07132_, _07131_, _07091_);
  nand (_07133_, _07132_, _07120_);
  nand (_07134_, _07133_, _07108_);
  and (_07135_, _07134_, _07107_);
  and (_07136_, _07135_, _06289_);
  nor (_07137_, _06418_, _05973_);
  nor (_07138_, _06253_, _06801_);
  and (_07139_, _07138_, _07137_);
  nor (_07140_, _07139_, _05957_);
  not (_07141_, _07140_);
  nor (_07142_, _07141_, _07136_);
  and (_07143_, _06338_, _06357_);
  not (_07144_, _07143_);
  nor (_07145_, _07144_, _06181_);
  and (_07146_, _07145_, _06250_);
  nor (_07147_, _07146_, _07142_);
  and (_07148_, _06401_, _06280_);
  nor (_07149_, _06814_, _05948_);
  nor (_07150_, _07149_, _07148_);
  and (_07151_, _06801_, _06280_);
  and (_07152_, _06339_, _06357_);
  and (_07153_, _07152_, \oc8051_golden_model_1.SP [0]);
  nor (_07154_, _07153_, _07151_);
  and (_07155_, _07154_, _07150_);
  and (_07156_, _07155_, _07147_);
  nand (_07157_, _07134_, _07107_);
  nor (_07158_, _06253_, _06256_);
  nor (_07159_, _07158_, _05948_);
  and (_07160_, _07159_, _07157_);
  nor (_07161_, _07160_, _06287_);
  and (_07162_, _07161_, _07156_);
  nor (_07163_, _07162_, _06288_);
  nor (_07164_, _07163_, _06284_);
  not (_07165_, _07164_);
  and (_07166_, _07165_, _06283_);
  nor (_07167_, _05949_, _06766_);
  nor (_07168_, _07167_, _07166_);
  not (_07169_, _06354_);
  nor (_07170_, _07169_, _06181_);
  and (_07171_, _07170_, _06250_);
  nor (_07172_, _07171_, _06771_);
  and (_07173_, _07172_, _07168_);
  nor (_07174_, _07158_, _05954_);
  and (_07175_, _07174_, _07157_);
  not (_07176_, _07175_);
  and (_07177_, _07176_, _07173_);
  nor (_07178_, _06278_, _06181_);
  nor (_07179_, _06346_, _06181_);
  and (_07180_, _07179_, _06250_);
  nor (_07181_, _07180_, _07178_);
  and (_07182_, _07181_, _07177_);
  nor (_07183_, _07182_, _06279_);
  nor (_07184_, _07183_, _06276_);
  and (_07185_, _06276_, _06766_);
  or (_07186_, _07185_, _07184_);
  and (_07187_, _07186_, _06274_);
  nor (_07188_, _07187_, _06272_);
  nor (_07189_, _05946_, _06766_);
  not (_07190_, _07189_);
  and (_07191_, _06337_, _05802_);
  nor (_07192_, _07191_, _06334_);
  and (_07193_, _07192_, _07190_);
  not (_07194_, _07193_);
  nor (_07195_, _07194_, _07188_);
  nor (_07196_, _06267_, _06181_);
  nor (_07197_, _07158_, _05952_);
  and (_07198_, _07197_, _07157_);
  nor (_07199_, _07198_, _07196_);
  and (_07200_, _07199_, _07195_);
  nor (_07201_, _07200_, _06268_);
  nor (_07202_, _07201_, _05974_);
  and (_07203_, _05974_, _06766_);
  nor (_07204_, _07203_, _07202_);
  not (_07205_, _06003_);
  nor (_07206_, _06770_, _07205_);
  or (_07207_, _07206_, _07204_);
  nor (_07208_, _07207_, _06264_);
  nor (_07209_, _07158_, _07205_);
  and (_07210_, _07209_, _07157_);
  nor (_07211_, _07210_, _06217_);
  and (_07212_, _07211_, _07208_);
  nor (_07213_, _07212_, _06249_);
  nor (_07214_, _07213_, _06004_);
  and (_07215_, _06004_, _06766_);
  nor (_07216_, _07215_, _07214_);
  not (_07217_, _06532_);
  nor (_07218_, _07217_, _06181_);
  not (_07219_, _06426_);
  and (_07220_, _06525_, _07219_);
  nor (_07221_, _07220_, _06181_);
  nor (_07222_, _07221_, _07218_);
  nor (_07223_, _07222_, _06248_);
  nor (_07224_, _07223_, _06013_);
  not (_07225_, _07224_);
  nor (_07226_, _07225_, _07216_);
  and (_07227_, _06013_, _06766_);
  nor (_07228_, _07227_, _07226_);
  not (_07229_, _06437_);
  nor (_07230_, _07229_, _06181_);
  not (_07231_, _06535_);
  nor (_07232_, _07231_, _06181_);
  nor (_07233_, _07232_, _07230_);
  nor (_07234_, _07233_, _06248_);
  nor (_07235_, _07234_, _07228_);
  and (_07236_, _06011_, \oc8051_golden_model_1.SP [0]);
  nor (_07237_, _06770_, _06913_);
  nor (_07238_, _07237_, _07236_);
  and (_07239_, _07238_, _07235_);
  not (_07240_, _06559_);
  nor (_07241_, _07240_, _06181_);
  and (_07242_, _06253_, _05895_);
  and (_07243_, _06256_, _05895_);
  nor (_07244_, _07243_, _07242_);
  not (_07245_, _07244_);
  and (_07246_, _07245_, _07157_);
  nor (_07247_, _07246_, _07241_);
  and (_07248_, _07247_, _07239_);
  and (_07249_, _07241_, _06248_);
  nor (_07250_, _07249_, _07248_);
  nor (_07251_, _06181_, _05933_);
  nor (_07252_, _06432_, _05991_);
  nor (_07253_, _07252_, _06766_);
  nor (_07254_, _07253_, _07251_);
  not (_07255_, _07254_);
  nor (_07256_, _07255_, _07250_);
  nor (_07257_, _07256_, _06214_);
  nor (_07258_, _07257_, _05891_);
  and (_07259_, _07258_, _05886_);
  and (_07260_, _06256_, _05766_);
  or (_07261_, _07260_, _06923_);
  and (_07262_, _07261_, _07157_);
  not (_07263_, _07262_);
  and (_07264_, _07263_, _07259_);
  nor (_07265_, _06570_, _06181_);
  and (_07266_, _07265_, _06250_);
  not (_07267_, _07266_);
  and (_07268_, _07267_, _07264_);
  and (_07269_, _06714_, _05766_);
  and (_07270_, _06962_, _05932_);
  not (_07271_, \oc8051_golden_model_1.SP [1]);
  and (_07272_, _07271_, \oc8051_golden_model_1.SP [0]);
  and (_07273_, \oc8051_golden_model_1.SP [1], _06766_);
  nor (_07274_, _07273_, _07272_);
  not (_07275_, _07274_);
  and (_07276_, _07275_, _06011_);
  and (_07277_, _06996_, _06217_);
  and (_07278_, _06962_, _06266_);
  and (_07279_, _07275_, _06276_);
  and (_07280_, _06996_, _06287_);
  nor (_07281_, _07158_, _05957_);
  not (_07282_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_07283_, _06929_, _07282_);
  not (_07284_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_07285_, _07078_, _07284_);
  and (_07286_, _07285_, _07076_);
  nand (_07287_, _07286_, _07283_);
  not (_07288_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_07289_, _07078_, _07288_);
  not (_07290_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_07291_, _06929_, _07290_);
  and (_07292_, _07291_, _07084_);
  nand (_07293_, _07292_, _07289_);
  nand (_07294_, _07293_, _07287_);
  nand (_07295_, _07294_, _06738_);
  not (_07296_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_07297_, _07078_, _07296_);
  not (_07298_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_07299_, _06929_, _07298_);
  and (_07300_, _07299_, _07084_);
  nand (_07301_, _07300_, _07297_);
  not (_07302_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_07303_, _06929_, _07302_);
  not (_07304_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_07305_, _07078_, _07304_);
  and (_07306_, _07305_, _07076_);
  nand (_07307_, _07306_, _07303_);
  nand (_07308_, _07307_, _07301_);
  nand (_07309_, _07308_, _07091_);
  nand (_07310_, _07309_, _07295_);
  nand (_07311_, _07310_, _06573_);
  nand (_07312_, _06929_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_07313_, _07078_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_07314_, _07313_, _07084_);
  nand (_07315_, _07314_, _07312_);
  nand (_07316_, _07078_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_07317_, _06929_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_07318_, _07317_, _07076_);
  nand (_07319_, _07318_, _07316_);
  nand (_07320_, _07319_, _07315_);
  nand (_07321_, _07320_, _06738_);
  nand (_07322_, _06929_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_07323_, _07078_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_07324_, _07323_, _07084_);
  nand (_07325_, _07324_, _07322_);
  nand (_07326_, _07078_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_07327_, _06929_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_07328_, _07327_, _07076_);
  nand (_07329_, _07328_, _07326_);
  nand (_07330_, _07329_, _07325_);
  nand (_07331_, _07330_, _07091_);
  nand (_07332_, _07331_, _07321_);
  nand (_07333_, _07332_, _07108_);
  nand (_07334_, _07333_, _07311_);
  and (_07335_, _07334_, _06289_);
  or (_07336_, _07335_, _07281_);
  and (_07337_, _07145_, _06995_);
  nor (_07338_, _07337_, _07336_);
  and (_07339_, _07274_, _07152_);
  not (_07340_, _07339_);
  and (_07341_, _06414_, _06280_);
  nor (_07342_, _07341_, _06720_);
  and (_07343_, _07342_, _07340_);
  and (_07344_, _07343_, _07338_);
  and (_07345_, _07334_, _07159_);
  nor (_07346_, _07345_, _06287_);
  and (_07347_, _07346_, _07344_);
  nor (_07348_, _07347_, _07280_);
  and (_07349_, _06961_, _06284_);
  or (_07350_, _07349_, _07348_);
  nor (_07351_, _07275_, _05949_);
  or (_07352_, _07351_, _07350_);
  and (_07353_, _07170_, _06995_);
  and (_07354_, _06414_, _06275_);
  nor (_07355_, _07354_, _06719_);
  not (_07356_, _07355_);
  nor (_07357_, _07356_, _07353_);
  not (_07358_, _07357_);
  nor (_07359_, _07358_, _07352_);
  and (_07360_, _07334_, _07174_);
  nor (_07361_, _07360_, _07179_);
  and (_07362_, _07361_, _07359_);
  and (_07363_, _07179_, _06996_);
  nor (_07364_, _07363_, _07362_);
  and (_07365_, _06961_, _07178_);
  nor (_07366_, _07365_, _07364_);
  and (_07367_, _07366_, _06778_);
  nor (_07368_, _07367_, _07279_);
  and (_07369_, _06961_, _06273_);
  or (_07370_, _07369_, _07368_);
  nor (_07371_, _07275_, _05946_);
  not (_07372_, _07371_);
  and (_07373_, _06414_, _06336_);
  and (_07374_, _06714_, _06336_);
  nor (_07375_, _07374_, _07373_);
  and (_07376_, _07375_, _07372_);
  not (_07377_, _07376_);
  nor (_07378_, _07377_, _07370_);
  and (_07379_, _07334_, _07197_);
  nor (_07380_, _07379_, _07196_);
  and (_07381_, _07380_, _07378_);
  nor (_07382_, _07381_, _07278_);
  nor (_07383_, _07382_, _05974_);
  and (_07384_, _07275_, _05974_);
  nor (_07385_, _07384_, _07383_);
  and (_07386_, _06263_, _06995_);
  and (_07387_, _06003_, _05927_);
  and (_07388_, _07387_, _05879_);
  nor (_07389_, _07388_, _07386_);
  not (_07390_, _07389_);
  nor (_07391_, _07390_, _07385_);
  and (_07392_, _07334_, _07209_);
  nor (_07393_, _07392_, _06217_);
  and (_07394_, _07393_, _07391_);
  nor (_07395_, _07394_, _07277_);
  nor (_07396_, _07395_, _06004_);
  and (_07397_, _07275_, _06004_);
  nor (_07398_, _07397_, _07396_);
  nor (_07399_, _07222_, _06996_);
  nor (_07400_, _07399_, _06013_);
  not (_07401_, _07400_);
  nor (_07402_, _07401_, _07398_);
  and (_07403_, _07275_, _06013_);
  nor (_07404_, _07403_, _07402_);
  nor (_07405_, _06536_, _06181_);
  and (_07406_, _07405_, _06995_);
  or (_07407_, _07406_, _06011_);
  nor (_07408_, _07407_, _07404_);
  nor (_07409_, _07408_, _07276_);
  and (_07410_, _06414_, _05895_);
  not (_07411_, _07410_);
  nand (_07412_, _06714_, _05895_);
  and (_07413_, _07412_, _07411_);
  not (_07414_, _07413_);
  nor (_07415_, _07414_, _07409_);
  and (_07416_, _07334_, _07245_);
  nor (_07417_, _07416_, _07241_);
  and (_07418_, _07417_, _07415_);
  and (_07419_, _07241_, _06996_);
  nor (_07420_, _07419_, _07418_);
  nor (_07421_, _07275_, _07252_);
  nor (_07422_, _07421_, _07251_);
  not (_07423_, _07422_);
  nor (_07424_, _07423_, _07420_);
  nor (_07425_, _07424_, _07270_);
  and (_07426_, _06414_, _05766_);
  or (_07427_, _07426_, _07425_);
  nor (_07428_, _07427_, _07269_);
  and (_07429_, _07334_, _07261_);
  nor (_07430_, _07429_, _07265_);
  and (_07431_, _07430_, _07428_);
  and (_07432_, _07265_, _06996_);
  nor (_07433_, _07432_, _07431_);
  not (_07434_, _00000_);
  and (_07435_, _06337_, _06252_);
  nor (_07436_, _07435_, _07209_);
  nor (_07437_, _07373_, _07159_);
  and (_07438_, _07437_, _07436_);
  not (_07439_, _07261_);
  and (_07440_, _07439_, _07244_);
  nor (_07441_, _07197_, _07174_);
  and (_07442_, _07441_, _07440_);
  and (_07443_, _07442_, _07438_);
  not (_07444_, _06414_);
  not (_07445_, _06409_);
  and (_07446_, _07034_, _07445_);
  and (_07447_, _07446_, _07444_);
  nor (_07448_, _07447_, _07205_);
  and (_07449_, _07444_, _07158_);
  nor (_07450_, _07449_, _05957_);
  not (_07451_, _05970_);
  nand (_07452_, _07137_, _07451_);
  and (_07453_, _07452_, _06757_);
  nor (_07454_, _07453_, _07450_);
  not (_07455_, _07454_);
  nor (_07456_, _07455_, _07448_);
  and (_07457_, _07456_, _07443_);
  not (_07458_, _05946_);
  nor (_07459_, _05974_, _07458_);
  not (_07460_, _05949_);
  nor (_07461_, _06004_, _07460_);
  and (_07462_, _07461_, _07459_);
  and (_07463_, _06702_, _06280_);
  nor (_07464_, _07341_, _07463_);
  and (_07465_, _05887_, _05895_);
  or (_07466_, _06339_, _06702_);
  and (_07467_, _07466_, _06003_);
  nor (_07468_, _07467_, _07465_);
  and (_07469_, _07468_, _07464_);
  and (_07470_, _07469_, _07462_);
  not (_07471_, _07045_);
  nor (_07472_, _06407_, _06409_);
  and (_07473_, _07472_, _06780_);
  nor (_07474_, _07473_, _05952_);
  nor (_07475_, _07474_, _07471_);
  and (_07476_, _07475_, _07470_);
  nor (_07477_, _07046_, _07152_);
  nor (_07478_, _07426_, _06719_);
  and (_07479_, _07478_, _07477_);
  and (_07480_, _07252_, _06014_);
  and (_07481_, _07480_, _07479_);
  and (_07482_, _05887_, _05766_);
  nor (_07483_, _07354_, _07482_);
  nor (_07484_, _07410_, _06276_);
  and (_07485_, _07484_, _07483_);
  nor (_07486_, _07034_, _06913_);
  nor (_07487_, _07486_, _06720_);
  nor (_07488_, _06711_, _06341_);
  and (_07489_, _07488_, _07487_);
  and (_07490_, _07489_, _07485_);
  and (_07491_, _07490_, _07481_);
  and (_07492_, _07491_, _07476_);
  and (_07493_, _07492_, _07457_);
  not (_07494_, _07493_);
  nor (_07495_, _07494_, _07221_);
  nor (_07496_, _06273_, _06287_);
  nor (_07497_, _07265_, _07170_);
  and (_07498_, _07497_, _07496_);
  and (_07499_, _07498_, _07495_);
  not (_07500_, _07405_);
  nor (_07501_, _07241_, _07218_);
  and (_07502_, _07501_, _07500_);
  nor (_07503_, _07179_, _07196_);
  nor (_07504_, _06284_, _07178_);
  and (_07505_, _07504_, _07503_);
  nor (_07506_, _06181_, _06251_);
  nor (_07507_, _07506_, _07251_);
  not (_07508_, _07466_);
  and (_07509_, _07508_, _07446_);
  nor (_07510_, _07509_, _05983_);
  not (_07511_, _07510_);
  and (_07512_, _06414_, _05971_);
  nor (_07513_, _07512_, _07143_);
  and (_07514_, _07513_, _06258_);
  and (_07515_, _07514_, _07511_);
  nor (_07516_, _07515_, _06181_);
  nor (_07517_, _07516_, _06217_);
  and (_07518_, _07517_, _07507_);
  and (_07519_, _07518_, _07505_);
  and (_07520_, _07519_, _07502_);
  and (_07521_, _07520_, _07499_);
  nor (_07522_, _07521_, _07434_);
  not (_07523_, _07522_);
  nor (_07524_, _07523_, _07433_);
  and (_07525_, _07524_, _07268_);
  not (_07526_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_07527_, _06929_, _07526_);
  not (_07528_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_07529_, _07078_, _07528_);
  and (_07530_, _07529_, _07076_);
  nand (_07531_, _07530_, _07527_);
  not (_07532_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_07533_, _07078_, _07532_);
  not (_07534_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_07535_, _06929_, _07534_);
  and (_07536_, _07535_, _07084_);
  nand (_07537_, _07536_, _07533_);
  nand (_07538_, _07537_, _07531_);
  nand (_07539_, _07538_, _06738_);
  not (_07540_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_07541_, _07078_, _07540_);
  not (_07542_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_07543_, _06929_, _07542_);
  and (_07544_, _07543_, _07084_);
  nand (_07545_, _07544_, _07541_);
  not (_07546_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_07547_, _06929_, _07546_);
  not (_07548_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_07549_, _07078_, _07548_);
  and (_07550_, _07549_, _07076_);
  nand (_07551_, _07550_, _07547_);
  nand (_07552_, _07551_, _07545_);
  nand (_07553_, _07552_, _07091_);
  nand (_07554_, _07553_, _07539_);
  nand (_07555_, _07554_, _06573_);
  nand (_07556_, _06929_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_07557_, _07078_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_07558_, _07557_, _07084_);
  nand (_07559_, _07558_, _07556_);
  nand (_07560_, _07078_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_07561_, _06929_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_07562_, _07561_, _07076_);
  nand (_07563_, _07562_, _07560_);
  nand (_07564_, _07563_, _07559_);
  nand (_07565_, _07564_, _06738_);
  nand (_07566_, _06929_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_07567_, _07078_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_07568_, _07567_, _07084_);
  nand (_07569_, _07568_, _07566_);
  nand (_07570_, _07078_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_07571_, _06929_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_07572_, _07571_, _07076_);
  nand (_07573_, _07572_, _07570_);
  nand (_07574_, _07573_, _07569_);
  nand (_07575_, _07574_, _07091_);
  nand (_07576_, _07575_, _07565_);
  nand (_07577_, _07576_, _07108_);
  nand (_07578_, _07577_, _07555_);
  and (_07579_, _07578_, _07261_);
  and (_07580_, _07578_, _07209_);
  and (_07581_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_07582_, _07581_, \oc8051_golden_model_1.SP [2]);
  nor (_07583_, _07582_, \oc8051_golden_model_1.SP [3]);
  and (_07584_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_07585_, _07584_, \oc8051_golden_model_1.SP [3]);
  and (_07586_, _07585_, \oc8051_golden_model_1.SP [0]);
  nor (_07587_, _07586_, _07583_);
  and (_07588_, _07587_, _05974_);
  not (_07589_, _06325_);
  and (_07590_, _07589_, _07196_);
  and (_07591_, _07587_, _07458_);
  and (_07592_, _06325_, _06284_);
  and (_07593_, _07578_, _07159_);
  and (_07594_, _07587_, _07152_);
  and (_07595_, _07578_, _06289_);
  and (_07596_, _05958_, _06362_);
  nor (_07597_, _07596_, _07145_);
  not (_07598_, _07597_);
  nor (_07599_, _07598_, _07595_);
  and (_07600_, _07145_, _06356_);
  nor (_07601_, _07600_, _07599_);
  nor (_07602_, _07601_, _07152_);
  or (_07603_, _07602_, _07159_);
  nor (_07604_, _07603_, _07594_);
  or (_07605_, _07604_, _06287_);
  nor (_07606_, _07605_, _07593_);
  and (_07607_, _06287_, _06356_);
  or (_07608_, _07607_, _06284_);
  nor (_07609_, _07608_, _07606_);
  nor (_07610_, _07609_, _07592_);
  nor (_07611_, _07610_, _07460_);
  nor (_07612_, _07587_, _05949_);
  nor (_07613_, _07612_, _07170_);
  not (_07614_, _07613_);
  nor (_07615_, _07614_, _07611_);
  and (_07616_, _07170_, _06356_);
  nor (_07617_, _07616_, _07174_);
  not (_07618_, _07617_);
  nor (_07619_, _07618_, _07615_);
  and (_07620_, _07578_, _07174_);
  nor (_07621_, _07620_, _07179_);
  not (_07622_, _07621_);
  nor (_07623_, _07622_, _07619_);
  and (_07624_, _07179_, _06356_);
  or (_07625_, _07624_, _07178_);
  nor (_07626_, _07625_, _07623_);
  and (_07627_, _06325_, _07178_);
  nor (_07628_, _07627_, _07626_);
  and (_07629_, _07628_, _06778_);
  and (_07630_, _07587_, _06276_);
  nor (_07631_, _07630_, _07629_);
  nor (_07632_, _07631_, _06273_);
  nor (_07633_, _06274_, _06328_);
  or (_07634_, _07633_, _07632_);
  and (_07635_, _07634_, _05946_);
  or (_07636_, _07635_, _07197_);
  nor (_07637_, _07636_, _07591_);
  and (_07638_, _07578_, _07197_);
  nor (_07639_, _07638_, _07196_);
  not (_07640_, _07639_);
  nor (_07641_, _07640_, _07637_);
  nor (_07642_, _07641_, _07590_);
  nor (_07643_, _07642_, _05974_);
  nor (_07644_, _07643_, _07588_);
  nor (_07645_, _07644_, _06263_);
  and (_07646_, _06263_, _06356_);
  nor (_07647_, _07646_, _07209_);
  not (_07648_, _07647_);
  nor (_07649_, _07648_, _07645_);
  or (_07650_, _07649_, _06217_);
  nor (_07651_, _07650_, _07580_);
  nor (_07652_, _06216_, _06213_);
  nor (_07653_, _07652_, _07651_);
  nor (_07654_, _07653_, _06004_);
  and (_07655_, _07587_, _06004_);
  not (_07656_, _07655_);
  and (_07657_, _07656_, _07222_);
  not (_07658_, _07657_);
  nor (_07659_, _07658_, _07654_);
  nor (_07660_, _07222_, _06356_);
  nor (_07661_, _07660_, _06013_);
  not (_07662_, _07661_);
  nor (_07663_, _07662_, _07659_);
  and (_07664_, _07587_, _06013_);
  or (_07665_, _07664_, _07405_);
  nor (_07666_, _07665_, _07663_);
  and (_07667_, _07405_, _06212_);
  or (_07668_, _07667_, _06011_);
  nor (_07669_, _07668_, _07666_);
  and (_07670_, _07587_, _06011_);
  nor (_07671_, _07670_, _07245_);
  not (_07672_, _07671_);
  nor (_07673_, _07672_, _07669_);
  and (_07674_, _07578_, _07245_);
  nor (_07675_, _07674_, _07241_);
  not (_07676_, _07675_);
  nor (_07677_, _07676_, _07673_);
  not (_07678_, _07252_);
  and (_07679_, _07241_, _06356_);
  nor (_07680_, _07679_, _07678_);
  not (_07681_, _07680_);
  nor (_07682_, _07681_, _07677_);
  nor (_07683_, _07587_, _07252_);
  nor (_07684_, _07683_, _07251_);
  not (_07685_, _07684_);
  nor (_07686_, _07685_, _07682_);
  and (_07687_, _07251_, _07589_);
  nor (_07688_, _07687_, _07261_);
  not (_07689_, _07688_);
  nor (_07690_, _07689_, _07686_);
  or (_07691_, _07690_, _07265_);
  nor (_07692_, _07691_, _07579_);
  and (_07693_, _07265_, _06356_);
  nor (_07694_, _07693_, _07692_);
  and (_07695_, _06605_, _05932_);
  nor (_07696_, _07581_, \oc8051_golden_model_1.SP [2]);
  nor (_07697_, _07696_, _07582_);
  and (_07698_, _07697_, _06011_);
  and (_07699_, _06647_, _06217_);
  and (_07700_, _06605_, _06266_);
  and (_07701_, _07697_, _06276_);
  and (_07702_, _06605_, _06281_);
  and (_07703_, _06647_, _06287_);
  not (_07704_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_07705_, _06929_, _07704_);
  not (_07706_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_07707_, _07078_, _07706_);
  and (_07708_, _07707_, _07076_);
  nand (_07709_, _07708_, _07705_);
  not (_07710_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_07711_, _07078_, _07710_);
  not (_07712_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_07713_, _06929_, _07712_);
  and (_07714_, _07713_, _07084_);
  nand (_07715_, _07714_, _07711_);
  nand (_07716_, _07715_, _07709_);
  nand (_07717_, _07716_, _06738_);
  not (_07718_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_07719_, _07078_, _07718_);
  not (_07720_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_07721_, _06929_, _07720_);
  and (_07722_, _07721_, _07084_);
  nand (_07723_, _07722_, _07719_);
  not (_07724_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_07725_, _06929_, _07724_);
  not (_07726_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_07727_, _07078_, _07726_);
  and (_07728_, _07727_, _07076_);
  nand (_07729_, _07728_, _07725_);
  nand (_07730_, _07729_, _07723_);
  nand (_07731_, _07730_, _07091_);
  nand (_07732_, _07731_, _07717_);
  nand (_07733_, _07732_, _06573_);
  not (_07734_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_07735_, _07078_, _07734_);
  not (_07736_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_07737_, _06929_, _07736_);
  and (_07738_, _07737_, _07084_);
  nand (_07739_, _07738_, _07735_);
  nand (_07740_, _07078_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_07741_, _06929_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_07742_, _07741_, _07076_);
  nand (_07743_, _07742_, _07740_);
  nand (_07744_, _07743_, _07739_);
  nand (_07745_, _07744_, _06738_);
  not (_07746_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_07747_, _07078_, _07746_);
  not (_07748_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_07749_, _06929_, _07748_);
  and (_07750_, _07749_, _07084_);
  nand (_07751_, _07750_, _07747_);
  nand (_07752_, _07078_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_07753_, _06929_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_07754_, _07753_, _07076_);
  nand (_07755_, _07754_, _07752_);
  nand (_07756_, _07755_, _07751_);
  nand (_07757_, _07756_, _07091_);
  nand (_07758_, _07757_, _07745_);
  nand (_07759_, _07758_, _07108_);
  nand (_07760_, _07759_, _07733_);
  or (_07761_, _07760_, _05942_);
  and (_07762_, _07761_, _07453_);
  and (_07763_, _07145_, _06646_);
  nor (_07764_, _07763_, _07762_);
  not (_07765_, _07697_);
  and (_07766_, _07765_, _07152_);
  not (_07767_, _07766_);
  nor (_07768_, _07044_, _07341_);
  and (_07769_, _07768_, _07767_);
  and (_07770_, _07769_, _07764_);
  and (_07771_, _07760_, _07159_);
  nor (_07772_, _07771_, _06287_);
  and (_07773_, _07772_, _07770_);
  nor (_07774_, _07773_, _07703_);
  nor (_07775_, _07774_, _06284_);
  nor (_07776_, _07775_, _07702_);
  nor (_07777_, _07697_, _05949_);
  nor (_07778_, _07777_, _07776_);
  and (_07779_, _07170_, _06646_);
  and (_07780_, _05882_, _06275_);
  nor (_07781_, _07780_, _07779_);
  and (_07782_, _07781_, _07778_);
  and (_07783_, _07760_, _07174_);
  nor (_07784_, _07783_, _07179_);
  and (_07785_, _07784_, _07782_);
  and (_07786_, _07179_, _06647_);
  nor (_07787_, _07786_, _07785_);
  and (_07788_, _06604_, _07178_);
  nor (_07789_, _07788_, _07787_);
  and (_07790_, _07789_, _06778_);
  nor (_07791_, _07790_, _07701_);
  and (_07792_, _06273_, _06604_);
  or (_07793_, _07792_, _07791_);
  nor (_07794_, _07697_, _05946_);
  nor (_07795_, _07794_, _06337_);
  not (_07796_, _07795_);
  nor (_07797_, _07796_, _07793_);
  and (_07798_, _07760_, _07197_);
  nor (_07799_, _07798_, _07196_);
  and (_07800_, _07799_, _07797_);
  nor (_07801_, _07800_, _07700_);
  nor (_07802_, _07801_, _05974_);
  and (_07803_, _07697_, _05974_);
  nor (_07804_, _07803_, _07802_);
  and (_07805_, _06263_, _06646_);
  and (_07806_, _05882_, _06003_);
  nor (_07807_, _07806_, _07805_);
  not (_07808_, _07807_);
  nor (_07809_, _07808_, _07804_);
  and (_07810_, _07760_, _07209_);
  nor (_07811_, _07810_, _06217_);
  and (_07812_, _07811_, _07809_);
  nor (_07813_, _07812_, _07699_);
  nor (_07814_, _07813_, _06004_);
  and (_07815_, _07697_, _06004_);
  nor (_07816_, _07815_, _07814_);
  nor (_07817_, _07222_, _06647_);
  nor (_07818_, _07817_, _06013_);
  not (_07819_, _07818_);
  nor (_07820_, _07819_, _07816_);
  and (_07821_, _07697_, _06013_);
  nor (_07822_, _07821_, _07820_);
  and (_07823_, _07405_, _06646_);
  or (_07824_, _07823_, _06011_);
  nor (_07825_, _07824_, _07822_);
  nor (_07826_, _07825_, _07698_);
  and (_07827_, _05882_, _05895_);
  nor (_07828_, _07827_, _07826_);
  and (_07829_, _07760_, _07245_);
  nor (_07830_, _07829_, _07241_);
  and (_07831_, _07830_, _07828_);
  and (_07832_, _07241_, _06647_);
  nor (_07833_, _07832_, _07831_);
  nor (_07834_, _07697_, _07252_);
  nor (_07835_, _07834_, _07251_);
  not (_07836_, _07835_);
  nor (_07837_, _07836_, _07833_);
  nor (_07838_, _07837_, _07695_);
  nor (_07839_, _07426_, _07043_);
  not (_07840_, _07839_);
  nor (_07841_, _07840_, _07838_);
  and (_07842_, _07760_, _07261_);
  nor (_07843_, _07842_, _07265_);
  and (_07844_, _07843_, _07841_);
  and (_07845_, _07265_, _06647_);
  nor (_07846_, _07845_, _07844_);
  nor (_07847_, _07846_, _07523_);
  not (_07848_, _07847_);
  nor (_07849_, _07848_, _07694_);
  and (_07850_, _07849_, _07525_);
  or (_07851_, _07850_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_07852_, _07584_, _06766_);
  nor (_07853_, _07697_, _07273_);
  nor (_07854_, _07853_, _07852_);
  and (_07855_, _07585_, _06766_);
  nor (_07856_, _07852_, _07587_);
  nor (_07857_, _07856_, _07855_);
  not (_07858_, _07152_);
  and (_07859_, _07252_, _07858_);
  and (_07860_, _07859_, _06014_);
  and (_07861_, _07860_, _07462_);
  nor (_07862_, _07861_, _07434_);
  and (_07863_, _07862_, _07857_);
  and (_07864_, _07863_, _07854_);
  and (_07865_, _07864_, _07272_);
  not (_07866_, _07865_);
  and (_07867_, _07866_, _07851_);
  not (_07868_, _07850_);
  and (_07869_, _06995_, _06250_);
  and (_07870_, _06646_, _06212_);
  and (_07871_, _07870_, _07869_);
  and (_07872_, _06325_, _06181_);
  not (_07873_, _06604_);
  and (_07874_, _06961_, _07873_);
  and (_07875_, _07874_, _07872_);
  and (_07876_, _07875_, _07871_);
  and (_07877_, _07876_, \oc8051_golden_model_1.P2 [7]);
  not (_07878_, _07877_);
  and (_07879_, _06646_, _06356_);
  and (_07880_, _07879_, _07869_);
  and (_07881_, _07875_, _07880_);
  and (_07882_, _07881_, \oc8051_golden_model_1.IE [7]);
  nor (_07883_, _06961_, _06604_);
  and (_07884_, _07883_, _07872_);
  and (_07885_, _07884_, _07871_);
  and (_07886_, _07885_, \oc8051_golden_model_1.P3 [7]);
  nor (_07887_, _07886_, _07882_);
  and (_07888_, _07887_, _07878_);
  not (_07889_, _06961_);
  and (_07890_, _07889_, _06604_);
  and (_07891_, _07890_, _07872_);
  and (_07892_, _06995_, _06248_);
  and (_07893_, _07892_, _07879_);
  and (_07894_, _07893_, _07891_);
  and (_07895_, _07894_, \oc8051_golden_model_1.SBUF [7]);
  and (_07896_, _06961_, _06604_);
  and (_07897_, _07896_, _07872_);
  nor (_07898_, _06646_, _06212_);
  and (_07899_, _07892_, _07898_);
  and (_07900_, _07899_, _07897_);
  and (_07901_, _07900_, \oc8051_golden_model_1.TH1 [7]);
  nor (_07902_, _07901_, _07895_);
  and (_07903_, _07902_, _07888_);
  and (_07904_, _07893_, _07897_);
  and (_07905_, _07904_, \oc8051_golden_model_1.TMOD [7]);
  not (_07906_, _07905_);
  and (_07907_, _07898_, _07869_);
  and (_07908_, _07907_, _07897_);
  and (_07909_, _07908_, \oc8051_golden_model_1.TH0 [7]);
  nor (_07910_, _06995_, _06248_);
  and (_07911_, _07910_, _07879_);
  and (_07912_, _07911_, _07897_);
  and (_07913_, _07912_, \oc8051_golden_model_1.TL0 [7]);
  nor (_07914_, _07913_, _07909_);
  and (_07915_, _07914_, _07906_);
  and (_07916_, _07880_, _07897_);
  and (_07917_, _07916_, \oc8051_golden_model_1.TCON [7]);
  and (_07918_, _07892_, _07870_);
  and (_07919_, _07918_, _07897_);
  and (_07920_, _07919_, \oc8051_golden_model_1.SP [7]);
  nor (_07921_, _07920_, _07917_);
  and (_07922_, _07921_, _07915_);
  and (_07923_, _07922_, _07903_);
  nor (_07924_, _06325_, _06294_);
  and (_07925_, _07924_, _07890_);
  and (_07926_, _07925_, _07871_);
  and (_07927_, _07926_, \oc8051_golden_model_1.PSW [7]);
  not (_07928_, _07927_);
  and (_07929_, _07924_, _07874_);
  and (_07930_, _07929_, _07871_);
  and (_07931_, _07930_, \oc8051_golden_model_1.ACC [7]);
  and (_07932_, _07883_, _07924_);
  and (_07933_, _07932_, _07871_);
  and (_07934_, _07933_, \oc8051_golden_model_1.B [7]);
  nor (_07935_, _07934_, _07931_);
  and (_07936_, _07935_, _07928_);
  and (_07937_, _07884_, _07880_);
  and (_07938_, _07937_, \oc8051_golden_model_1.IP [7]);
  and (_07939_, _07897_, _06212_);
  nor (_07940_, _06995_, _06250_);
  and (_07941_, _07940_, _06647_);
  and (_07942_, _07941_, _07939_);
  and (_07943_, _07942_, \oc8051_golden_model_1.PCON [7]);
  nor (_07944_, _07943_, _07938_);
  and (_07945_, _07944_, _07936_);
  and (_07946_, _07897_, _07871_);
  and (_07947_, _07946_, \oc8051_golden_model_1.P0 [7]);
  not (_07948_, _07947_);
  and (_07949_, _07910_, _06646_);
  and (_07950_, _07949_, _07939_);
  and (_07951_, _07950_, \oc8051_golden_model_1.DPL [7]);
  and (_07952_, _07940_, _07870_);
  and (_07953_, _07952_, _07897_);
  and (_07954_, _07953_, \oc8051_golden_model_1.DPH [7]);
  nor (_07955_, _07954_, _07951_);
  and (_07956_, _07955_, _07948_);
  and (_07957_, _07940_, _07879_);
  and (_07958_, _07957_, _07897_);
  and (_07959_, _07958_, \oc8051_golden_model_1.TL1 [7]);
  not (_07960_, _07959_);
  and (_07961_, _07891_, _07871_);
  and (_07962_, _07961_, \oc8051_golden_model_1.P1 [7]);
  and (_07963_, _07880_, _07891_);
  and (_07964_, _07963_, \oc8051_golden_model_1.SCON [7]);
  nor (_07965_, _07964_, _07962_);
  and (_07966_, _07965_, _07960_);
  and (_07967_, _07966_, _07956_);
  and (_07968_, _07967_, _07945_);
  and (_07969_, _07968_, _07923_);
  not (_07970_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_07971_, _06929_, _07970_);
  not (_07972_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_07973_, _07078_, _07972_);
  and (_07974_, _07973_, _07076_);
  nand (_07975_, _07974_, _07971_);
  not (_07976_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_07977_, _07078_, _07976_);
  not (_07978_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_07979_, _06929_, _07978_);
  and (_07980_, _07979_, _07084_);
  nand (_07981_, _07980_, _07977_);
  nand (_07982_, _07981_, _07975_);
  nand (_07983_, _07982_, _06738_);
  not (_07984_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_07985_, _07078_, _07984_);
  not (_07986_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_07987_, _06929_, _07986_);
  and (_07988_, _07987_, _07084_);
  nand (_07989_, _07988_, _07985_);
  not (_07990_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_07991_, _06929_, _07990_);
  not (_07992_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_07993_, _07078_, _07992_);
  and (_07994_, _07993_, _07076_);
  nand (_07995_, _07994_, _07991_);
  nand (_07996_, _07995_, _07989_);
  nand (_07997_, _07996_, _07091_);
  nand (_07998_, _07997_, _07983_);
  nand (_07999_, _07998_, _06573_);
  nand (_08000_, _06929_, \oc8051_golden_model_1.IRAM[11] [7]);
  not (_08001_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_08002_, _06929_, _08001_);
  and (_08003_, _08002_, _07084_);
  nand (_08004_, _08003_, _08000_);
  nand (_08005_, _07078_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_08006_, _06929_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_08007_, _08006_, _07076_);
  nand (_08008_, _08007_, _08005_);
  nand (_08009_, _08008_, _08004_);
  nand (_08010_, _08009_, _06738_);
  nand (_08011_, _06929_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_08012_, _07078_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_08013_, _08012_, _07084_);
  nand (_08014_, _08013_, _08011_);
  nand (_08015_, _07078_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_08016_, _06929_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_08017_, _08016_, _07076_);
  nand (_08018_, _08017_, _08015_);
  nand (_08019_, _08018_, _08014_);
  nand (_08020_, _08019_, _07091_);
  nand (_08021_, _08020_, _08010_);
  nand (_08022_, _08021_, _07108_);
  nand (_08023_, _08022_, _07999_);
  or (_08024_, _08023_, _06181_);
  and (_08025_, _08024_, _07969_);
  not (_08026_, _08025_);
  and (_08027_, _07876_, \oc8051_golden_model_1.P2 [6]);
  not (_08028_, _08027_);
  and (_08029_, _07894_, \oc8051_golden_model_1.SBUF [6]);
  not (_08030_, _08029_);
  and (_08031_, _07881_, \oc8051_golden_model_1.IE [6]);
  and (_08032_, _07885_, \oc8051_golden_model_1.P3 [6]);
  nor (_08033_, _08032_, _08031_);
  and (_08034_, _08033_, _08030_);
  and (_08035_, _08034_, _08028_);
  and (_08036_, _07946_, \oc8051_golden_model_1.P0 [6]);
  not (_08037_, _08036_);
  and (_08038_, _07950_, \oc8051_golden_model_1.DPL [6]);
  and (_08039_, _07953_, \oc8051_golden_model_1.DPH [6]);
  nor (_08040_, _08039_, _08038_);
  and (_08041_, _08040_, _08037_);
  and (_08042_, _07958_, \oc8051_golden_model_1.TL1 [6]);
  and (_08043_, _07900_, \oc8051_golden_model_1.TH1 [6]);
  nor (_08044_, _08043_, _08042_);
  and (_08045_, _07963_, \oc8051_golden_model_1.SCON [6]);
  and (_08046_, _07961_, \oc8051_golden_model_1.P1 [6]);
  nor (_08047_, _08046_, _08045_);
  and (_08048_, _08047_, _08044_);
  and (_08049_, _08048_, _08041_);
  and (_08050_, _08049_, _08035_);
  and (_08051_, _07937_, \oc8051_golden_model_1.IP [6]);
  not (_08052_, _08051_);
  and (_08053_, _07933_, \oc8051_golden_model_1.B [6]);
  and (_08054_, _07930_, \oc8051_golden_model_1.ACC [6]);
  nor (_08055_, _08054_, _08053_);
  and (_08056_, _08055_, _08052_);
  and (_08057_, _07942_, \oc8051_golden_model_1.PCON [6]);
  and (_08058_, _07926_, \oc8051_golden_model_1.PSW [6]);
  nor (_08059_, _08058_, _08057_);
  and (_08060_, _08059_, _08056_);
  and (_08061_, _07916_, \oc8051_golden_model_1.TCON [6]);
  not (_08062_, _08061_);
  and (_08063_, _07912_, \oc8051_golden_model_1.TL0 [6]);
  and (_08064_, _07908_, \oc8051_golden_model_1.TH0 [6]);
  nor (_08065_, _08064_, _08063_);
  and (_08066_, _08065_, _08062_);
  and (_08067_, _07904_, \oc8051_golden_model_1.TMOD [6]);
  and (_08068_, _07919_, \oc8051_golden_model_1.SP [6]);
  nor (_08069_, _08068_, _08067_);
  and (_08070_, _08069_, _08066_);
  and (_08071_, _08070_, _08060_);
  and (_08072_, _08071_, _08050_);
  not (_08073_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_08074_, _06929_, _08073_);
  not (_08075_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_08076_, _07078_, _08075_);
  and (_08077_, _08076_, _07076_);
  nand (_08078_, _08077_, _08074_);
  not (_08079_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_08080_, _07078_, _08079_);
  not (_08081_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_08082_, _06929_, _08081_);
  and (_08083_, _08082_, _07084_);
  nand (_08084_, _08083_, _08080_);
  nand (_08085_, _08084_, _08078_);
  nand (_08086_, _08085_, _06738_);
  not (_08087_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_08088_, _07078_, _08087_);
  not (_08089_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_08090_, _06929_, _08089_);
  and (_08091_, _08090_, _07084_);
  nand (_08092_, _08091_, _08088_);
  not (_08093_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_08094_, _06929_, _08093_);
  not (_08095_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_08096_, _07078_, _08095_);
  and (_08097_, _08096_, _07076_);
  nand (_08098_, _08097_, _08094_);
  nand (_08099_, _08098_, _08092_);
  nand (_08100_, _08099_, _07091_);
  nand (_08101_, _08100_, _08086_);
  nand (_08102_, _08101_, _06573_);
  nand (_08103_, _06929_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_08104_, _07078_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_08105_, _08104_, _07084_);
  nand (_08106_, _08105_, _08103_);
  nand (_08107_, _07078_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_08108_, _06929_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_08109_, _08108_, _07076_);
  nand (_08110_, _08109_, _08107_);
  nand (_08111_, _08110_, _08106_);
  nand (_08112_, _08111_, _06738_);
  nand (_08113_, _06929_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_08114_, _07078_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_08115_, _08114_, _07084_);
  nand (_08116_, _08115_, _08113_);
  nand (_08117_, _07078_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_08118_, _06929_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_08119_, _08118_, _07076_);
  nand (_08120_, _08119_, _08117_);
  nand (_08121_, _08120_, _08116_);
  nand (_08122_, _08121_, _07091_);
  nand (_08123_, _08122_, _08112_);
  nand (_08124_, _08123_, _07108_);
  nand (_08125_, _08124_, _08102_);
  or (_08126_, _08125_, _06181_);
  and (_08127_, _08126_, _08072_);
  not (_08128_, _08127_);
  and (_08129_, _07876_, \oc8051_golden_model_1.P2 [5]);
  not (_08130_, _08129_);
  and (_08131_, _07881_, \oc8051_golden_model_1.IE [5]);
  and (_08132_, _07885_, \oc8051_golden_model_1.P3 [5]);
  nor (_08133_, _08132_, _08131_);
  and (_08134_, _08133_, _08130_);
  and (_08135_, _07894_, \oc8051_golden_model_1.SBUF [5]);
  and (_08136_, _07900_, \oc8051_golden_model_1.TH1 [5]);
  nor (_08137_, _08136_, _08135_);
  and (_08138_, _08137_, _08134_);
  and (_08139_, _07916_, \oc8051_golden_model_1.TCON [5]);
  not (_08140_, _08139_);
  and (_08141_, _07908_, \oc8051_golden_model_1.TH0 [5]);
  and (_08142_, _07912_, \oc8051_golden_model_1.TL0 [5]);
  nor (_08143_, _08142_, _08141_);
  and (_08144_, _08143_, _08140_);
  and (_08145_, _07904_, \oc8051_golden_model_1.TMOD [5]);
  and (_08146_, _07919_, \oc8051_golden_model_1.SP [5]);
  nor (_08147_, _08146_, _08145_);
  and (_08148_, _08147_, _08144_);
  and (_08149_, _08148_, _08138_);
  and (_08150_, _07926_, \oc8051_golden_model_1.PSW [5]);
  not (_08151_, _08150_);
  and (_08152_, _07930_, \oc8051_golden_model_1.ACC [5]);
  and (_08153_, _07933_, \oc8051_golden_model_1.B [5]);
  nor (_08154_, _08153_, _08152_);
  and (_08155_, _08154_, _08151_);
  and (_08156_, _07937_, \oc8051_golden_model_1.IP [5]);
  and (_08157_, _07942_, \oc8051_golden_model_1.PCON [5]);
  nor (_08158_, _08157_, _08156_);
  and (_08159_, _08158_, _08155_);
  and (_08160_, _07946_, \oc8051_golden_model_1.P0 [5]);
  not (_08161_, _08160_);
  and (_08162_, _07950_, \oc8051_golden_model_1.DPL [5]);
  and (_08163_, _07953_, \oc8051_golden_model_1.DPH [5]);
  nor (_08164_, _08163_, _08162_);
  and (_08165_, _08164_, _08161_);
  and (_08166_, _07958_, \oc8051_golden_model_1.TL1 [5]);
  not (_08167_, _08166_);
  and (_08168_, _07961_, \oc8051_golden_model_1.P1 [5]);
  and (_08169_, _07963_, \oc8051_golden_model_1.SCON [5]);
  nor (_08170_, _08169_, _08168_);
  and (_08171_, _08170_, _08167_);
  and (_08172_, _08171_, _08165_);
  and (_08173_, _08172_, _08159_);
  and (_08174_, _08173_, _08149_);
  not (_08175_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_08176_, _06929_, _08175_);
  not (_08177_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_08178_, _07078_, _08177_);
  and (_08179_, _08178_, _07076_);
  nand (_08180_, _08179_, _08176_);
  not (_08181_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_08182_, _07078_, _08181_);
  not (_08183_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_08184_, _06929_, _08183_);
  and (_08185_, _08184_, _07084_);
  nand (_08186_, _08185_, _08182_);
  nand (_08187_, _08186_, _08180_);
  nand (_08188_, _08187_, _06738_);
  not (_08189_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_08190_, _07078_, _08189_);
  not (_08191_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_08192_, _06929_, _08191_);
  and (_08193_, _08192_, _07084_);
  nand (_08194_, _08193_, _08190_);
  not (_08195_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_08196_, _06929_, _08195_);
  not (_08197_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_08198_, _07078_, _08197_);
  and (_08199_, _08198_, _07076_);
  nand (_08200_, _08199_, _08196_);
  nand (_08201_, _08200_, _08194_);
  nand (_08202_, _08201_, _07091_);
  nand (_08203_, _08202_, _08188_);
  nand (_08204_, _08203_, _06573_);
  nand (_08205_, _06929_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_08206_, _07078_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_08207_, _08206_, _07084_);
  nand (_08208_, _08207_, _08205_);
  nand (_08209_, _07078_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_08210_, _06929_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_08211_, _08210_, _07076_);
  nand (_08212_, _08211_, _08209_);
  nand (_08213_, _08212_, _08208_);
  nand (_08214_, _08213_, _06738_);
  not (_08215_, \oc8051_golden_model_1.IRAM[15] [5]);
  or (_08216_, _07078_, _08215_);
  nand (_08217_, _07078_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_08218_, _08217_, _07084_);
  nand (_08219_, _08218_, _08216_);
  nand (_08220_, _07078_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_08221_, _06929_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_08222_, _08221_, _07076_);
  nand (_08223_, _08222_, _08220_);
  nand (_08224_, _08223_, _08219_);
  nand (_08225_, _08224_, _07091_);
  nand (_08226_, _08225_, _08214_);
  nand (_08227_, _08226_, _07108_);
  nand (_08228_, _08227_, _08204_);
  or (_08229_, _08228_, _06181_);
  and (_08230_, _08229_, _08174_);
  not (_08231_, _08230_);
  and (_08232_, _07926_, \oc8051_golden_model_1.PSW [3]);
  and (_08233_, _07930_, \oc8051_golden_model_1.ACC [3]);
  nor (_08234_, _08233_, _08232_);
  and (_08235_, _07894_, \oc8051_golden_model_1.SBUF [3]);
  and (_08236_, _07933_, \oc8051_golden_model_1.B [3]);
  nor (_08237_, _08236_, _08235_);
  and (_08238_, _08237_, _08234_);
  and (_08239_, _07881_, \oc8051_golden_model_1.IE [3]);
  and (_08240_, _07885_, \oc8051_golden_model_1.P3 [3]);
  nor (_08241_, _08240_, _08239_);
  and (_08242_, _07876_, \oc8051_golden_model_1.P2 [3]);
  and (_08243_, _07937_, \oc8051_golden_model_1.IP [3]);
  nor (_08244_, _08243_, _08242_);
  and (_08245_, _08244_, _08241_);
  and (_08246_, _07904_, \oc8051_golden_model_1.TMOD [3]);
  and (_08247_, _07958_, \oc8051_golden_model_1.TL1 [3]);
  nor (_08248_, _08247_, _08246_);
  and (_08249_, _07912_, \oc8051_golden_model_1.TL0 [3]);
  and (_08250_, _07963_, \oc8051_golden_model_1.SCON [3]);
  nor (_08251_, _08250_, _08249_);
  and (_08252_, _08251_, _08248_);
  and (_08253_, _08252_, _08245_);
  and (_08254_, _08253_, _08238_);
  and (_08255_, _07892_, _06646_);
  and (_08256_, _07939_, _08255_);
  and (_08257_, _08256_, \oc8051_golden_model_1.SP [3]);
  not (_08258_, _08257_);
  and (_08259_, _07942_, \oc8051_golden_model_1.PCON [3]);
  and (_08260_, _07940_, _06646_);
  and (_08261_, _08260_, _07939_);
  and (_08262_, _08261_, \oc8051_golden_model_1.DPH [3]);
  nor (_08263_, _08262_, _08259_);
  and (_08264_, _08263_, _08258_);
  and (_08265_, _07908_, \oc8051_golden_model_1.TH0 [3]);
  and (_08266_, _07900_, \oc8051_golden_model_1.TH1 [3]);
  nor (_08267_, _08266_, _08265_);
  and (_08268_, _07916_, \oc8051_golden_model_1.TCON [3]);
  and (_08269_, _07961_, \oc8051_golden_model_1.P1 [3]);
  nor (_08270_, _08269_, _08268_);
  and (_08271_, _08270_, _08267_);
  and (_08272_, _07946_, \oc8051_golden_model_1.P0 [3]);
  and (_08273_, _07950_, \oc8051_golden_model_1.DPL [3]);
  nor (_08274_, _08273_, _08272_);
  and (_08275_, _08274_, _08271_);
  and (_08276_, _08275_, _08264_);
  and (_08277_, _08276_, _08254_);
  or (_08278_, _07578_, _06181_);
  and (_08279_, _08278_, _08277_);
  not (_08280_, _08279_);
  and (_08281_, _07926_, \oc8051_golden_model_1.PSW [1]);
  and (_08282_, _07933_, \oc8051_golden_model_1.B [1]);
  nor (_08283_, _08282_, _08281_);
  and (_08284_, _07894_, \oc8051_golden_model_1.SBUF [1]);
  and (_08285_, _07881_, \oc8051_golden_model_1.IE [1]);
  nor (_08286_, _08285_, _08284_);
  and (_08287_, _08286_, _08283_);
  and (_08288_, _07912_, \oc8051_golden_model_1.TL0 [1]);
  and (_08289_, _07930_, \oc8051_golden_model_1.ACC [1]);
  nor (_08290_, _08289_, _08288_);
  and (_08291_, _07908_, \oc8051_golden_model_1.TH0 [1]);
  and (_08292_, _07885_, \oc8051_golden_model_1.P3 [1]);
  nor (_08293_, _08292_, _08291_);
  and (_08294_, _08293_, _08290_);
  and (_08295_, _07961_, \oc8051_golden_model_1.P1 [1]);
  and (_08296_, _07876_, \oc8051_golden_model_1.P2 [1]);
  nor (_08297_, _08296_, _08295_);
  and (_08298_, _07963_, \oc8051_golden_model_1.SCON [1]);
  and (_08299_, _07937_, \oc8051_golden_model_1.IP [1]);
  nor (_08300_, _08299_, _08298_);
  and (_08301_, _08300_, _08297_);
  and (_08302_, _08301_, _08294_);
  and (_08303_, _08302_, _08287_);
  and (_08304_, _07946_, \oc8051_golden_model_1.P0 [1]);
  not (_08305_, _08304_);
  and (_08306_, _07950_, \oc8051_golden_model_1.DPL [1]);
  and (_08307_, _08256_, \oc8051_golden_model_1.SP [1]);
  nor (_08308_, _08307_, _08306_);
  and (_08309_, _08308_, _08305_);
  and (_08310_, _07958_, \oc8051_golden_model_1.TL1 [1]);
  and (_08311_, _07900_, \oc8051_golden_model_1.TH1 [1]);
  nor (_08312_, _08311_, _08310_);
  and (_08313_, _07916_, \oc8051_golden_model_1.TCON [1]);
  and (_08314_, _07904_, \oc8051_golden_model_1.TMOD [1]);
  nor (_08315_, _08314_, _08313_);
  and (_08316_, _08315_, _08312_);
  and (_08317_, _07942_, \oc8051_golden_model_1.PCON [1]);
  and (_08318_, _08261_, \oc8051_golden_model_1.DPH [1]);
  nor (_08319_, _08318_, _08317_);
  and (_08320_, _08319_, _08316_);
  and (_08321_, _08320_, _08309_);
  and (_08322_, _08321_, _08303_);
  or (_08323_, _07334_, _06181_);
  and (_08324_, _08323_, _08322_);
  not (_08325_, _08324_);
  and (_08326_, _07876_, \oc8051_golden_model_1.P2 [0]);
  not (_08327_, _08326_);
  and (_08328_, _07881_, \oc8051_golden_model_1.IE [0]);
  and (_08329_, _07885_, \oc8051_golden_model_1.P3 [0]);
  nor (_08330_, _08329_, _08328_);
  and (_08331_, _07894_, \oc8051_golden_model_1.SBUF [0]);
  not (_08332_, _08331_);
  and (_08333_, _08332_, _08330_);
  and (_08334_, _08333_, _08327_);
  and (_08335_, _07946_, \oc8051_golden_model_1.P0 [0]);
  not (_08336_, _08335_);
  and (_08337_, _07950_, \oc8051_golden_model_1.DPL [0]);
  and (_08338_, _07953_, \oc8051_golden_model_1.DPH [0]);
  nor (_08339_, _08338_, _08337_);
  and (_08340_, _08339_, _08336_);
  and (_08341_, _07961_, \oc8051_golden_model_1.P1 [0]);
  and (_08342_, _07963_, \oc8051_golden_model_1.SCON [0]);
  nor (_08343_, _08342_, _08341_);
  and (_08344_, _07900_, \oc8051_golden_model_1.TH1 [0]);
  and (_08345_, _07958_, \oc8051_golden_model_1.TL1 [0]);
  nor (_08346_, _08345_, _08344_);
  and (_08347_, _08346_, _08343_);
  and (_08348_, _08347_, _08340_);
  and (_08349_, _08348_, _08334_);
  and (_08350_, _07926_, \oc8051_golden_model_1.PSW [0]);
  not (_08351_, _08350_);
  and (_08352_, _07933_, \oc8051_golden_model_1.B [0]);
  and (_08353_, _07930_, \oc8051_golden_model_1.ACC [0]);
  nor (_08354_, _08353_, _08352_);
  and (_08355_, _08354_, _08351_);
  and (_08356_, _07937_, \oc8051_golden_model_1.IP [0]);
  and (_08357_, _07942_, \oc8051_golden_model_1.PCON [0]);
  nor (_08358_, _08357_, _08356_);
  and (_08359_, _08358_, _08355_);
  and (_08360_, _07904_, \oc8051_golden_model_1.TMOD [0]);
  not (_08361_, _08360_);
  and (_08362_, _07912_, \oc8051_golden_model_1.TL0 [0]);
  and (_08363_, _07908_, \oc8051_golden_model_1.TH0 [0]);
  nor (_08364_, _08363_, _08362_);
  and (_08365_, _08364_, _08361_);
  and (_08366_, _07916_, \oc8051_golden_model_1.TCON [0]);
  and (_08367_, _07919_, \oc8051_golden_model_1.SP [0]);
  nor (_08368_, _08367_, _08366_);
  and (_08369_, _08368_, _08365_);
  and (_08370_, _08369_, _08359_);
  and (_08371_, _08370_, _08349_);
  not (_08372_, _08371_);
  and (_08373_, _07135_, _06294_);
  or (_08374_, _08373_, _08372_);
  and (_08375_, _08374_, _08325_);
  and (_08376_, _07894_, \oc8051_golden_model_1.SBUF [2]);
  not (_08377_, _08376_);
  and (_08378_, _07885_, \oc8051_golden_model_1.P3 [2]);
  and (_08379_, _07881_, \oc8051_golden_model_1.IE [2]);
  nor (_08380_, _08379_, _08378_);
  and (_08381_, _08380_, _08377_);
  and (_08382_, _07876_, \oc8051_golden_model_1.P2 [2]);
  and (_08383_, _07900_, \oc8051_golden_model_1.TH1 [2]);
  nor (_08384_, _08383_, _08382_);
  and (_08385_, _08384_, _08381_);
  and (_08386_, _07904_, \oc8051_golden_model_1.TMOD [2]);
  not (_08387_, _08386_);
  and (_08388_, _07912_, \oc8051_golden_model_1.TL0 [2]);
  and (_08389_, _07908_, \oc8051_golden_model_1.TH0 [2]);
  nor (_08390_, _08389_, _08388_);
  and (_08391_, _08390_, _08387_);
  and (_08392_, _07916_, \oc8051_golden_model_1.TCON [2]);
  and (_08393_, _07946_, \oc8051_golden_model_1.P0 [2]);
  nor (_08394_, _08393_, _08392_);
  and (_08395_, _08394_, _08391_);
  and (_08396_, _08395_, _08385_);
  and (_08397_, _07926_, \oc8051_golden_model_1.PSW [2]);
  not (_08398_, _08397_);
  and (_08399_, _07930_, \oc8051_golden_model_1.ACC [2]);
  and (_08400_, _07933_, \oc8051_golden_model_1.B [2]);
  nor (_08401_, _08400_, _08399_);
  and (_08402_, _08401_, _08398_);
  and (_08403_, _07937_, \oc8051_golden_model_1.IP [2]);
  and (_08404_, _07942_, \oc8051_golden_model_1.PCON [2]);
  nor (_08405_, _08404_, _08403_);
  and (_08406_, _08405_, _08402_);
  and (_08407_, _07919_, \oc8051_golden_model_1.SP [2]);
  not (_08408_, _08407_);
  and (_08409_, _07950_, \oc8051_golden_model_1.DPL [2]);
  and (_08410_, _07953_, \oc8051_golden_model_1.DPH [2]);
  nor (_08411_, _08410_, _08409_);
  and (_08412_, _08411_, _08408_);
  and (_08413_, _07958_, \oc8051_golden_model_1.TL1 [2]);
  not (_08414_, _08413_);
  and (_08415_, _07961_, \oc8051_golden_model_1.P1 [2]);
  and (_08416_, _07963_, \oc8051_golden_model_1.SCON [2]);
  nor (_08417_, _08416_, _08415_);
  and (_08418_, _08417_, _08414_);
  and (_08419_, _08418_, _08412_);
  and (_08420_, _08419_, _08406_);
  and (_08421_, _08420_, _08396_);
  or (_08422_, _07760_, _06181_);
  and (_08423_, _08422_, _08421_);
  not (_08424_, _08423_);
  and (_08425_, _08424_, _08375_);
  and (_08426_, _08425_, _08280_);
  and (_08427_, _07894_, \oc8051_golden_model_1.SBUF [4]);
  not (_08428_, _08427_);
  and (_08429_, _07876_, \oc8051_golden_model_1.P2 [4]);
  not (_08430_, _08429_);
  and (_08431_, _07885_, \oc8051_golden_model_1.P3 [4]);
  and (_08432_, _07881_, \oc8051_golden_model_1.IE [4]);
  nor (_08433_, _08432_, _08431_);
  and (_08434_, _08433_, _08430_);
  and (_08435_, _08434_, _08428_);
  and (_08436_, _07919_, \oc8051_golden_model_1.SP [4]);
  not (_08437_, _08436_);
  and (_08438_, _07950_, \oc8051_golden_model_1.DPL [4]);
  and (_08439_, _07953_, \oc8051_golden_model_1.DPH [4]);
  nor (_08440_, _08439_, _08438_);
  and (_08441_, _08440_, _08437_);
  and (_08442_, _07961_, \oc8051_golden_model_1.P1 [4]);
  and (_08443_, _07963_, \oc8051_golden_model_1.SCON [4]);
  nor (_08444_, _08443_, _08442_);
  and (_08445_, _07900_, \oc8051_golden_model_1.TH1 [4]);
  and (_08446_, _07958_, \oc8051_golden_model_1.TL1 [4]);
  nor (_08447_, _08446_, _08445_);
  and (_08448_, _08447_, _08444_);
  and (_08449_, _08448_, _08441_);
  and (_08450_, _08449_, _08435_);
  and (_08451_, _07937_, \oc8051_golden_model_1.IP [4]);
  not (_08452_, _08451_);
  and (_08453_, _07930_, \oc8051_golden_model_1.ACC [4]);
  and (_08454_, _07933_, \oc8051_golden_model_1.B [4]);
  nor (_08455_, _08454_, _08453_);
  and (_08456_, _08455_, _08452_);
  and (_08457_, _07926_, \oc8051_golden_model_1.PSW [4]);
  and (_08458_, _07942_, \oc8051_golden_model_1.PCON [4]);
  nor (_08459_, _08458_, _08457_);
  and (_08460_, _08459_, _08456_);
  and (_08461_, _07904_, \oc8051_golden_model_1.TMOD [4]);
  not (_08462_, _08461_);
  and (_08463_, _07912_, \oc8051_golden_model_1.TL0 [4]);
  and (_08464_, _07908_, \oc8051_golden_model_1.TH0 [4]);
  nor (_08465_, _08464_, _08463_);
  and (_08466_, _08465_, _08462_);
  and (_08467_, _07916_, \oc8051_golden_model_1.TCON [4]);
  and (_08468_, _07946_, \oc8051_golden_model_1.P0 [4]);
  nor (_08469_, _08468_, _08467_);
  and (_08470_, _08469_, _08466_);
  and (_08471_, _08470_, _08460_);
  and (_08472_, _08471_, _08450_);
  not (_08473_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_08474_, _06929_, _08473_);
  not (_08475_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_08476_, _07078_, _08475_);
  and (_08477_, _08476_, _07076_);
  nand (_08478_, _08477_, _08474_);
  not (_08479_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_08480_, _07078_, _08479_);
  not (_08481_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_08482_, _06929_, _08481_);
  and (_08483_, _08482_, _07084_);
  nand (_08484_, _08483_, _08480_);
  nand (_08485_, _08484_, _08478_);
  nand (_08486_, _08485_, _06738_);
  not (_08487_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_08488_, _07078_, _08487_);
  not (_08489_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_08490_, _06929_, _08489_);
  and (_08491_, _08490_, _07084_);
  nand (_08492_, _08491_, _08488_);
  not (_08493_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_08494_, _06929_, _08493_);
  not (_08495_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_08496_, _07078_, _08495_);
  and (_08497_, _08496_, _07076_);
  nand (_08498_, _08497_, _08494_);
  nand (_08499_, _08498_, _08492_);
  nand (_08500_, _08499_, _07091_);
  nand (_08501_, _08500_, _08486_);
  nand (_08502_, _08501_, _06573_);
  nand (_08503_, _06929_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_08504_, _07078_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_08505_, _08504_, _07084_);
  nand (_08506_, _08505_, _08503_);
  nand (_08507_, _07078_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_08508_, _06929_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_08509_, _08508_, _07076_);
  nand (_08510_, _08509_, _08507_);
  nand (_08511_, _08510_, _08506_);
  nand (_08512_, _08511_, _06738_);
  nand (_08513_, _06929_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_08514_, _07078_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_08515_, _08514_, _07084_);
  nand (_08516_, _08515_, _08513_);
  nand (_08517_, _07078_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_08518_, _06929_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_08519_, _08518_, _07076_);
  nand (_08520_, _08519_, _08517_);
  nand (_08521_, _08520_, _08516_);
  nand (_08522_, _08521_, _07091_);
  nand (_08523_, _08522_, _08512_);
  nand (_08524_, _08523_, _07108_);
  nand (_08525_, _08524_, _08502_);
  or (_08526_, _08525_, _06181_);
  and (_08527_, _08526_, _08472_);
  not (_08528_, _08527_);
  and (_08529_, _08528_, _08426_);
  and (_08530_, _08529_, _08231_);
  and (_08531_, _08530_, _08128_);
  nor (_08532_, _08531_, _08026_);
  and (_08533_, _08531_, _08026_);
  nor (_08534_, _08533_, _08532_);
  and (_08535_, _08534_, _07265_);
  and (_08536_, _08022_, _07999_);
  and (_08537_, _07334_, _07157_);
  and (_08538_, _08537_, _07760_);
  and (_08539_, _08538_, _07578_);
  and (_08540_, _08539_, _08525_);
  and (_08541_, _08540_, _08228_);
  and (_08542_, _08541_, _08125_);
  or (_08543_, _08542_, _08536_);
  nand (_08544_, _08542_, _08536_);
  and (_08545_, _08544_, _08543_);
  nor (_08546_, _07486_, _07465_);
  and (_08547_, _08546_, _07411_);
  or (_08548_, _08547_, _08545_);
  not (_08549_, _07218_);
  nor (_08550_, _07219_, _06181_);
  and (_08551_, _06462_, _04418_);
  not (_08552_, _08551_);
  and (_08553_, _06494_, _04400_);
  and (_08554_, _06496_, _04395_);
  nor (_08555_, _08554_, _08553_);
  and (_08556_, _06502_, _04413_);
  and (_08557_, _06500_, _04382_);
  nor (_08558_, _08557_, _08556_);
  and (_08559_, _08558_, _08555_);
  and (_08560_, _06506_, _04416_);
  and (_08561_, _06511_, _04388_);
  and (_08562_, _06509_, _04391_);
  or (_08563_, _08562_, _08561_);
  nor (_08564_, _08563_, _08560_);
  and (_08565_, _08564_, _08559_);
  and (_08566_, _06477_, _04432_);
  and (_08567_, _06474_, _04346_);
  nor (_08568_, _08567_, _08566_);
  and (_08569_, _06466_, _04404_);
  and (_08570_, _06469_, _04429_);
  nor (_08571_, _08570_, _08569_);
  and (_08572_, _08571_, _08568_);
  and (_08573_, _06481_, _04378_);
  and (_08574_, _06483_, _04373_);
  nor (_08575_, _08574_, _08573_);
  and (_08576_, _06487_, _04408_);
  and (_08577_, _06489_, _04423_);
  nor (_08578_, _08577_, _08576_);
  and (_08579_, _08578_, _08575_);
  and (_08580_, _08579_, _08572_);
  and (_08581_, _08580_, _08565_);
  and (_08582_, _08581_, _08552_);
  nor (_08583_, _08582_, _08025_);
  and (_08584_, _08583_, _08550_);
  not (_08585_, _07178_);
  nor (_08586_, _06962_, _06605_);
  and (_08587_, _08586_, _06213_);
  and (_08588_, _08587_, _06378_);
  and (_08589_, _08588_, _07884_);
  and (_08590_, _08589_, \oc8051_golden_model_1.IP [7]);
  and (_08591_, _08587_, _06328_);
  and (_08592_, _08591_, _07925_);
  and (_08593_, _08592_, \oc8051_golden_model_1.PSW [7]);
  and (_08594_, _08591_, _07932_);
  and (_08595_, _08594_, \oc8051_golden_model_1.B [7]);
  and (_08596_, _08591_, _07929_);
  and (_08597_, _08596_, \oc8051_golden_model_1.ACC [7]);
  or (_08598_, _08597_, _08595_);
  or (_08599_, _08598_, _08593_);
  and (_08600_, _08588_, _07897_);
  and (_08601_, _08600_, \oc8051_golden_model_1.TCON [7]);
  and (_08602_, _07939_, \oc8051_golden_model_1.P0 [7]);
  and (_08603_, _08591_, _07891_);
  and (_08604_, _08603_, \oc8051_golden_model_1.P1 [7]);
  or (_08605_, _08604_, _08602_);
  or (_08606_, _08605_, _08601_);
  and (_08607_, _08591_, _07884_);
  and (_08608_, _08607_, \oc8051_golden_model_1.P3 [7]);
  and (_08609_, _08588_, _07875_);
  and (_08610_, _08609_, \oc8051_golden_model_1.IE [7]);
  or (_08611_, _08610_, _08608_);
  and (_08612_, _08588_, _07891_);
  and (_08613_, _08612_, \oc8051_golden_model_1.SCON [7]);
  and (_08614_, _08591_, _07875_);
  and (_08615_, _08614_, \oc8051_golden_model_1.P2 [7]);
  or (_08616_, _08615_, _08613_);
  or (_08617_, _08616_, _08611_);
  or (_08618_, _08617_, _08606_);
  or (_08619_, _08618_, _08599_);
  nor (_08620_, _08619_, _08590_);
  and (_08621_, _08620_, _08024_);
  nor (_08622_, _08621_, _07941_);
  or (_08623_, _08622_, _08585_);
  not (_08624_, _06284_);
  not (_08625_, _07941_);
  nand (_08626_, _08621_, _08625_);
  or (_08627_, _08626_, _08624_);
  and (_08628_, _08527_, _08230_);
  not (_08629_, _08374_);
  and (_08630_, _08629_, _08324_);
  and (_08631_, _08423_, _08279_);
  and (_08632_, _08631_, _08630_);
  and (_08633_, _08632_, _08628_);
  and (_08634_, _08633_, _08127_);
  or (_08635_, _08634_, _08026_);
  nand (_08636_, _08634_, _08026_);
  and (_08637_, _08636_, _08635_);
  and (_08638_, _08637_, _06287_);
  not (_08639_, _07159_);
  not (_08640_, \oc8051_golden_model_1.SP [2]);
  nor (_08641_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_08642_, _08641_, _08640_);
  nor (_08643_, _08642_, _06353_);
  nor (_08644_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_08645_, _08644_, _06353_);
  and (_08646_, _08645_, _06766_);
  nor (_08647_, _08646_, _08643_);
  nor (_08648_, _06543_, _06290_);
  nor (_08649_, _08648_, _08647_);
  not (_08650_, _07197_);
  and (_08651_, _07578_, _08650_);
  and (_08652_, _07197_, _06212_);
  not (_08653_, _08652_);
  nand (_08654_, _08653_, _08648_);
  nor (_08655_, _08654_, _08651_);
  nor (_08656_, _08655_, _08649_);
  not (_08657_, _08656_);
  nor (_08658_, _08641_, _08640_);
  nor (_08659_, _08658_, _08642_);
  nor (_08660_, _08659_, _08648_);
  not (_08661_, _08660_);
  and (_08662_, _07759_, _07733_);
  or (_08663_, _08662_, _07197_);
  and (_08664_, _07197_, _06646_);
  not (_08665_, _08664_);
  and (_08666_, _08665_, _08648_);
  nand (_08667_, _08666_, _08663_);
  and (_08668_, _08667_, _08661_);
  or (_08669_, _07197_, _07135_);
  nor (_08670_, _08650_, _06248_);
  not (_08671_, _08670_);
  and (_08672_, _08671_, _08648_);
  nand (_08673_, _08672_, _08669_);
  nor (_08674_, _08648_, \oc8051_golden_model_1.SP [0]);
  not (_08675_, _08674_);
  and (_08676_, _08675_, _08673_);
  or (_08677_, _08676_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor (_08678_, _08648_, _07274_);
  not (_08679_, _08678_);
  or (_08680_, _07334_, _07197_);
  or (_08681_, _08650_, _06995_);
  and (_08682_, _08681_, _08648_);
  nand (_08683_, _08682_, _08680_);
  and (_08684_, _08683_, _08679_);
  not (_08685_, _08684_);
  not (_08686_, _08676_);
  or (_08687_, _08686_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_08688_, _08687_, _08685_);
  and (_08689_, _08688_, _08677_);
  nand (_08690_, _08676_, _08001_);
  or (_08691_, _08676_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_08692_, _08691_, _08684_);
  and (_08693_, _08692_, _08690_);
  nor (_08694_, _08693_, _08689_);
  nand (_08695_, _08694_, _08668_);
  not (_08696_, _08668_);
  or (_08697_, _08676_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_08698_, _08686_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_08699_, _08698_, _08685_);
  and (_08700_, _08699_, _08697_);
  or (_08701_, _08686_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_08702_, _08676_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_08703_, _08702_, _08684_);
  and (_08704_, _08703_, _08701_);
  nor (_08705_, _08704_, _08700_);
  nand (_08706_, _08705_, _08696_);
  nand (_08707_, _08706_, _08695_);
  nand (_08708_, _08707_, _08657_);
  or (_08709_, _08676_, _07972_);
  nand (_08710_, _08676_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_08711_, _08710_, _08685_);
  nand (_08712_, _08711_, _08709_);
  nand (_08713_, _08676_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_08714_, _08676_, _07976_);
  and (_08715_, _08714_, _08684_);
  nand (_08716_, _08715_, _08713_);
  nand (_08717_, _08716_, _08712_);
  nand (_08718_, _08717_, _08668_);
  nand (_08719_, _08676_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_08720_, _08676_, _07992_);
  and (_08721_, _08720_, _08685_);
  nand (_08722_, _08721_, _08719_);
  nand (_08723_, _08676_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_08724_, _08676_, _07984_);
  and (_08725_, _08724_, _08684_);
  nand (_08726_, _08725_, _08723_);
  nand (_08727_, _08726_, _08722_);
  nand (_08728_, _08727_, _08696_);
  nand (_08729_, _08728_, _08718_);
  nand (_08730_, _08729_, _08656_);
  and (_08731_, _08730_, _08708_);
  or (_08732_, _08731_, _08639_);
  not (_08733_, _06287_);
  nor (_08734_, _05948_, _05880_);
  and (_08735_, _08734_, _08545_);
  not (_08736_, _08734_);
  not (_08737_, \oc8051_golden_model_1.ACC [7]);
  nor (_08738_, _07152_, _08737_);
  and (_08739_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_08740_, _08739_, \oc8051_golden_model_1.PC [6]);
  and (_08741_, _08740_, _06093_);
  and (_08742_, _08741_, \oc8051_golden_model_1.PC [7]);
  nor (_08743_, _08741_, \oc8051_golden_model_1.PC [7]);
  nor (_08744_, _08743_, _08742_);
  and (_08745_, _08744_, _07152_);
  or (_08746_, _08745_, _08738_);
  and (_08747_, _08746_, _08736_);
  or (_08748_, _08747_, _07159_);
  or (_08749_, _08748_, _08735_);
  and (_08750_, _08749_, _08733_);
  and (_08751_, _08750_, _08732_);
  or (_08752_, _08751_, _08638_);
  or (_08753_, _08752_, _06284_);
  and (_08754_, _08753_, _08627_);
  or (_08755_, _08754_, _07460_);
  nor (_08756_, _08744_, _05949_);
  nor (_08757_, _08756_, _07170_);
  and (_08758_, _08757_, _08755_);
  and (_08759_, _08536_, _07170_);
  or (_08760_, _08759_, _07178_);
  or (_08761_, _08760_, _08758_);
  and (_08762_, _08761_, _08623_);
  or (_08763_, _08762_, _06276_);
  nand (_08764_, _08025_, _06276_);
  and (_08765_, _08764_, _06274_);
  and (_08766_, _08765_, _08763_);
  nor (_08767_, _08621_, _08625_);
  not (_08768_, _08767_);
  and (_08769_, _08768_, _08626_);
  and (_08770_, _08769_, _06273_);
  or (_08771_, _08770_, _08766_);
  and (_08772_, _08771_, _05946_);
  not (_08773_, _08744_);
  or (_08774_, _08773_, _05946_);
  nand (_08775_, _08774_, _06343_);
  or (_08776_, _08775_, _08772_);
  nand (_08777_, _08025_, _06344_);
  and (_08778_, _08777_, _08776_);
  or (_08779_, _08778_, _07197_);
  not (_08780_, _07196_);
  and (_08781_, _08731_, _06294_);
  nand (_08782_, _07969_, _07197_);
  or (_08783_, _08782_, _08781_);
  and (_08784_, _08783_, _08780_);
  and (_08785_, _08784_, _08779_);
  and (_08786_, _06248_, \oc8051_golden_model_1.PSW [7]);
  and (_08787_, _08786_, _06996_);
  and (_08788_, _08787_, _06647_);
  or (_08789_, _08788_, _08622_);
  and (_08790_, _08789_, _07196_);
  or (_08791_, _08790_, _05974_);
  or (_08792_, _08791_, _08785_);
  nor (_08793_, _06260_, _06181_);
  and (_08794_, _08773_, _05974_);
  nor (_08795_, _08794_, _08793_);
  and (_08796_, _08795_, _08792_);
  nor (_08797_, _06258_, _06181_);
  and (_08798_, _08536_, _08793_);
  or (_08799_, _08798_, _08797_);
  or (_08800_, _08799_, _08796_);
  not (_08801_, _07506_);
  not (_08802_, _08797_);
  or (_08803_, _08731_, _08802_);
  and (_08804_, _08803_, _08801_);
  and (_08805_, _08804_, _08800_);
  not (_08806_, _08582_);
  nor (_08807_, _08806_, _08023_);
  and (_08808_, _07031_, _06850_);
  not (_08809_, _06517_);
  and (_08810_, _06689_, _08809_);
  and (_08811_, _08810_, _08808_);
  and (_08812_, _06462_, _04833_);
  not (_08813_, _08812_);
  and (_08814_, _06469_, _04835_);
  and (_08815_, _06466_, _04820_);
  nor (_08816_, _08815_, _08814_);
  and (_08817_, _06474_, _04825_);
  and (_08818_, _06477_, _04842_);
  nor (_08819_, _08818_, _08817_);
  and (_08820_, _08819_, _08816_);
  and (_08821_, _06481_, _04809_);
  and (_08822_, _06483_, _04812_);
  nor (_08823_, _08822_, _08821_);
  and (_08824_, _06489_, _04814_);
  and (_08825_, _06487_, _04831_);
  nor (_08826_, _08825_, _08824_);
  and (_08827_, _08826_, _08823_);
  and (_08828_, _08827_, _08820_);
  and (_08829_, _06494_, _04840_);
  and (_08830_, _06496_, _04823_);
  nor (_08831_, _08830_, _08829_);
  and (_08832_, _06500_, _04829_);
  and (_08833_, _06502_, _04818_);
  nor (_08834_, _08833_, _08832_);
  and (_08835_, _08834_, _08831_);
  and (_08836_, _06506_, _04847_);
  not (_08837_, _08836_);
  and (_08838_, _06511_, _04849_);
  and (_08839_, _06509_, _04807_);
  nor (_08840_, _08839_, _08838_);
  and (_08841_, _08840_, _08837_);
  and (_08842_, _08841_, _08835_);
  and (_08843_, _08842_, _08828_);
  and (_08844_, _08843_, _08813_);
  not (_08845_, _08844_);
  nor (_08846_, _08845_, _08582_);
  and (_08847_, _06462_, _04715_);
  not (_08848_, _08847_);
  and (_08849_, _06494_, _04726_);
  and (_08850_, _06496_, _04724_);
  nor (_08851_, _08850_, _08849_);
  and (_08852_, _06500_, _04731_);
  and (_08853_, _06502_, _04729_);
  nor (_08854_, _08853_, _08852_);
  and (_08855_, _08854_, _08851_);
  and (_08856_, _06506_, _04719_);
  and (_08857_, _06511_, _04722_);
  and (_08858_, _06509_, _04717_);
  or (_08859_, _08858_, _08857_);
  nor (_08860_, _08859_, _08856_);
  and (_08861_, _08860_, _08855_);
  and (_08862_, _06466_, _04737_);
  and (_08863_, _06469_, _04739_);
  nor (_08864_, _08863_, _08862_);
  and (_08865_, _06474_, _04742_);
  and (_08866_, _06477_, _04744_);
  nor (_08867_, _08866_, _08865_);
  and (_08868_, _08867_, _08864_);
  and (_08869_, _06481_, _04748_);
  and (_08870_, _06483_, _04750_);
  nor (_08871_, _08870_, _08869_);
  and (_08873_, _06489_, _04753_);
  and (_08874_, _06487_, _04755_);
  nor (_08875_, _08874_, _08873_);
  and (_08876_, _08875_, _08871_);
  and (_08877_, _08876_, _08868_);
  and (_08878_, _08877_, _08861_);
  and (_08879_, _08878_, _08848_);
  and (_08880_, _06511_, _04803_);
  and (_08881_, _06487_, _04785_);
  or (_08882_, _08881_, _08880_);
  and (_08884_, _06509_, _04768_);
  and (_08885_, _06481_, _04763_);
  or (_08886_, _08885_, _08884_);
  or (_08887_, _08886_, _08882_);
  and (_08888_, _06506_, _04801_);
  and (_08889_, _06483_, _04761_);
  or (_08890_, _08889_, _08888_);
  and (_08891_, _06502_, _04796_);
  and (_08892_, _06489_, _04766_);
  or (_08893_, _08892_, _08891_);
  or (_08895_, _08893_, _08890_);
  or (_08896_, _08895_, _08887_);
  and (_08897_, _06477_, _04794_);
  and (_08898_, _06474_, _04777_);
  or (_08899_, _08898_, _08897_);
  and (_08900_, _06462_, _04787_);
  and (_08901_, _06466_, _04772_);
  or (_08902_, _08901_, _08900_);
  or (_08903_, _08902_, _08899_);
  and (_08904_, _06494_, _04774_);
  and (_08906_, _06500_, _04783_);
  or (_08907_, _08906_, _08904_);
  and (_08908_, _06496_, _04779_);
  and (_08909_, _06469_, _04789_);
  or (_08910_, _08909_, _08908_);
  or (_08911_, _08910_, _08907_);
  or (_08912_, _08911_, _08903_);
  or (_08913_, _08912_, _08896_);
  nor (_08914_, _08913_, _08879_);
  and (_08915_, _08914_, _08846_);
  and (_08917_, _08915_, _08811_);
  and (_08918_, _08917_, \oc8051_golden_model_1.SCON [7]);
  not (_08919_, _08879_);
  and (_08920_, _08913_, _08919_);
  and (_08921_, _06689_, _06517_);
  and (_08922_, _08921_, _08808_);
  nor (_08923_, _08844_, _08582_);
  and (_08924_, _08923_, _08922_);
  and (_08925_, _08924_, _08920_);
  and (_08926_, _08925_, \oc8051_golden_model_1.B [7]);
  or (_08928_, _08926_, _08918_);
  not (_08929_, _06850_);
  and (_08930_, _07031_, _08929_);
  and (_08931_, _08930_, _08810_);
  and (_08932_, _08931_, _08915_);
  and (_08933_, _08932_, \oc8051_golden_model_1.SBUF [7]);
  and (_08934_, _08913_, _08879_);
  and (_08935_, _08934_, _08924_);
  and (_08936_, _08935_, \oc8051_golden_model_1.ACC [7]);
  or (_08937_, _08936_, _08933_);
  or (_08939_, _08937_, _08928_);
  nor (_08940_, _08913_, _08919_);
  and (_08941_, _08940_, _08846_);
  and (_08942_, _08941_, _08811_);
  and (_08943_, _08942_, \oc8051_golden_model_1.TCON [7]);
  and (_08944_, _08922_, _08915_);
  and (_08945_, _08944_, \oc8051_golden_model_1.P1 [7]);
  or (_08946_, _08945_, _08943_);
  and (_08947_, _08941_, _08922_);
  and (_08948_, _08947_, \oc8051_golden_model_1.P0 [7]);
  nor (_08949_, _07031_, _08929_);
  and (_08950_, _08949_, _08810_);
  and (_08951_, _08950_, _08941_);
  and (_08952_, _08951_, \oc8051_golden_model_1.TL0 [7]);
  or (_08953_, _08952_, _08948_);
  or (_08954_, _08953_, _08946_);
  and (_08955_, _08934_, _08846_);
  and (_08956_, _08955_, _08922_);
  and (_08957_, _08956_, \oc8051_golden_model_1.P2 [7]);
  and (_08958_, _08920_, _08846_);
  and (_08959_, _08958_, _08922_);
  and (_08960_, _08959_, \oc8051_golden_model_1.P3 [7]);
  or (_08961_, _08960_, _08957_);
  and (_08962_, _08955_, _08811_);
  and (_08963_, _08962_, \oc8051_golden_model_1.IE [7]);
  and (_08964_, _08958_, _08811_);
  and (_08965_, _08964_, \oc8051_golden_model_1.IP [7]);
  or (_08966_, _08965_, _08963_);
  or (_08967_, _08966_, _08961_);
  and (_08968_, _08941_, _08931_);
  and (_08969_, _08968_, \oc8051_golden_model_1.TMOD [7]);
  and (_08970_, _08924_, _08914_);
  and (_08971_, _08970_, \oc8051_golden_model_1.PSW [7]);
  or (_08972_, _08971_, _08969_);
  or (_08973_, _08972_, _08967_);
  or (_08974_, _08973_, _08954_);
  or (_08975_, _08974_, _08939_);
  nor (_08976_, _07031_, _06850_);
  and (_08977_, _08976_, _08941_);
  and (_08978_, _08977_, _08921_);
  and (_08979_, _08978_, \oc8051_golden_model_1.DPH [7]);
  not (_08980_, _06689_);
  and (_08981_, _08980_, _06517_);
  and (_08982_, _08981_, _08977_);
  and (_08983_, _08982_, \oc8051_golden_model_1.PCON [7]);
  nor (_08984_, _06689_, _06517_);
  and (_08985_, _08984_, _08941_);
  and (_08986_, _08985_, _08808_);
  and (_08987_, _08986_, \oc8051_golden_model_1.TH0 [7]);
  or (_08988_, _08987_, _08983_);
  or (_08989_, _08988_, _08979_);
  and (_08990_, _08977_, _08810_);
  and (_08991_, _08990_, \oc8051_golden_model_1.TL1 [7]);
  and (_08992_, _08941_, _08921_);
  and (_08993_, _08992_, _08930_);
  and (_08994_, _08993_, \oc8051_golden_model_1.SP [7]);
  or (_08995_, _08994_, _08991_);
  and (_08996_, _08949_, _08992_);
  and (_08997_, _08996_, \oc8051_golden_model_1.DPL [7]);
  and (_08998_, _08985_, _08930_);
  and (_08999_, _08998_, \oc8051_golden_model_1.TH1 [7]);
  or (_09000_, _08999_, _08997_);
  or (_09001_, _09000_, _08995_);
  or (_09002_, _09001_, _08989_);
  or (_09003_, _09002_, _08975_);
  or (_09004_, _09003_, _08807_);
  and (_09005_, _09004_, _07506_);
  and (_09006_, _05882_, _05968_);
  not (_09007_, _09006_);
  nand (_09008_, _07446_, _09007_);
  and (_09009_, _09008_, _06003_);
  not (_09010_, _09009_);
  not (_09011_, _06256_);
  and (_09012_, _07138_, _09011_);
  nor (_09013_, _09012_, _07205_);
  nor (_09014_, _09013_, _07467_);
  and (_09015_, _09014_, _09010_);
  not (_09016_, _09015_);
  or (_09017_, _09016_, _09005_);
  or (_09018_, _09017_, _08805_);
  nor (_09019_, _09015_, _06181_);
  nor (_09020_, _09019_, _06217_);
  and (_09021_, _09020_, _09018_);
  and (_09022_, _08806_, _06217_);
  or (_09023_, _09022_, _06004_);
  or (_09024_, _09023_, _09021_);
  not (_09025_, _06398_);
  nor (_09026_, _09025_, _06181_);
  and (_09027_, _08773_, _06004_);
  nor (_09028_, _09027_, _09026_);
  and (_09029_, _09028_, _09024_);
  not (_09030_, _06524_);
  nor (_09031_, _09030_, _06181_);
  not (_09032_, _08583_);
  nand (_09033_, _08582_, _08025_);
  and (_09034_, _09033_, _09032_);
  and (_09035_, _09034_, _09026_);
  or (_09036_, _09035_, _09031_);
  or (_09037_, _09036_, _09029_);
  not (_09038_, _08550_);
  not (_09039_, _09031_);
  nor (_09040_, _08025_, _08737_);
  and (_09041_, _08025_, _08737_);
  nor (_09042_, _09041_, _09040_);
  or (_09043_, _09042_, _09039_);
  and (_09044_, _09043_, _09038_);
  and (_09045_, _09044_, _09037_);
  or (_09046_, _09045_, _08584_);
  and (_09047_, _09046_, _08549_);
  and (_09048_, _09040_, _07218_);
  or (_09049_, _09048_, _06013_);
  or (_09050_, _09049_, _09047_);
  and (_09051_, _08773_, _06013_);
  nor (_09052_, _09051_, _07230_);
  and (_09053_, _09052_, _09050_);
  and (_09054_, _09033_, _07230_);
  or (_09055_, _09054_, _07232_);
  or (_09056_, _09055_, _09053_);
  not (_09057_, _06011_);
  nand (_09058_, _09041_, _07232_);
  and (_09059_, _09058_, _09057_);
  and (_09060_, _09059_, _09056_);
  nand (_09061_, _08744_, _06011_);
  nand (_09062_, _09061_, _08547_);
  or (_09063_, _09062_, _09060_);
  and (_09064_, _09063_, _08548_);
  or (_09065_, _09064_, _07245_);
  not (_09066_, _07241_);
  nand (_09067_, _08730_, _08708_);
  or (_09068_, _08676_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_09069_, _08686_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_09070_, _09069_, _08685_);
  and (_09071_, _09070_, _09068_);
  or (_09072_, _08686_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_09073_, _08676_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_09074_, _09073_, _08684_);
  and (_09075_, _09074_, _09072_);
  nor (_09076_, _09075_, _09071_);
  nand (_09077_, _09076_, _08668_);
  or (_09078_, _08676_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_09079_, _08686_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_09080_, _09079_, _08685_);
  and (_09081_, _09080_, _09078_);
  or (_09082_, _08686_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_09083_, _08676_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_09084_, _09083_, _08684_);
  and (_09085_, _09084_, _09082_);
  nor (_09086_, _09085_, _09081_);
  nand (_09087_, _09086_, _08696_);
  nand (_09088_, _09087_, _09077_);
  nand (_09089_, _09088_, _08657_);
  or (_09090_, _08676_, _08075_);
  nand (_09091_, _08676_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_09092_, _09091_, _08685_);
  nand (_09093_, _09092_, _09090_);
  nand (_09094_, _08676_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_09095_, _08676_, _08079_);
  and (_09096_, _09095_, _08684_);
  nand (_09097_, _09096_, _09094_);
  nand (_09098_, _09097_, _09093_);
  nand (_09099_, _09098_, _08668_);
  nand (_09100_, _08676_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_09101_, _08676_, _08095_);
  and (_09102_, _09101_, _08685_);
  nand (_09103_, _09102_, _09100_);
  nand (_09104_, _08676_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_09105_, _08676_, _08087_);
  and (_09106_, _09105_, _08684_);
  nand (_09107_, _09106_, _09104_);
  nand (_09108_, _09107_, _09103_);
  nand (_09109_, _09108_, _08696_);
  nand (_09110_, _09109_, _09099_);
  nand (_09111_, _09110_, _08656_);
  nand (_09112_, _09111_, _09089_);
  or (_09113_, _08676_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_09114_, _08686_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_09115_, _09114_, _08685_);
  and (_09116_, _09115_, _09113_);
  or (_09117_, _08686_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_09118_, _08676_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_09119_, _09118_, _08684_);
  and (_09120_, _09119_, _09117_);
  nor (_09121_, _09120_, _09116_);
  nand (_09122_, _09121_, _08668_);
  or (_09123_, _08676_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_09124_, _08686_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_09125_, _09124_, _08685_);
  and (_09126_, _09125_, _09123_);
  or (_09127_, _08686_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_09128_, _08676_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_09129_, _09128_, _08684_);
  and (_09130_, _09129_, _09127_);
  nor (_09131_, _09130_, _09126_);
  nand (_09132_, _09131_, _08696_);
  nand (_09133_, _09132_, _09122_);
  nand (_09134_, _09133_, _08657_);
  or (_09135_, _08676_, _08177_);
  nand (_09136_, _08676_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_09137_, _09136_, _08685_);
  nand (_09138_, _09137_, _09135_);
  nand (_09139_, _08676_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_09140_, _08676_, _08181_);
  and (_09141_, _09140_, _08684_);
  nand (_09142_, _09141_, _09139_);
  nand (_09143_, _09142_, _09138_);
  nand (_09144_, _09143_, _08668_);
  nand (_09145_, _08676_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_09146_, _08676_, _08197_);
  and (_09147_, _09146_, _08685_);
  nand (_09148_, _09147_, _09145_);
  nand (_09149_, _08676_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_09150_, _08676_, _08189_);
  and (_09151_, _09150_, _08684_);
  nand (_09152_, _09151_, _09149_);
  nand (_09153_, _09152_, _09148_);
  nand (_09154_, _09153_, _08696_);
  nand (_09155_, _09154_, _09144_);
  nand (_09156_, _09155_, _08656_);
  nand (_09157_, _09156_, _09134_);
  or (_09158_, _08676_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_09159_, _08686_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_09160_, _09159_, _08685_);
  and (_09161_, _09160_, _09158_);
  or (_09162_, _08686_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_09163_, _08676_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_09164_, _09163_, _08684_);
  and (_09165_, _09164_, _09162_);
  nor (_09166_, _09165_, _09161_);
  nand (_09167_, _09166_, _08668_);
  or (_09168_, _08676_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_09169_, _08686_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_09170_, _09169_, _08685_);
  and (_09171_, _09170_, _09168_);
  or (_09172_, _08686_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_09173_, _08676_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_09174_, _09173_, _08684_);
  and (_09175_, _09174_, _09172_);
  nor (_09176_, _09175_, _09171_);
  nand (_09177_, _09176_, _08696_);
  nand (_09178_, _09177_, _09167_);
  nand (_09179_, _09178_, _08657_);
  or (_09180_, _08676_, _08475_);
  nand (_09181_, _08676_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_09182_, _09181_, _08685_);
  nand (_09183_, _09182_, _09180_);
  nand (_09184_, _08676_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_09185_, _08676_, _08479_);
  and (_09186_, _09185_, _08684_);
  nand (_09187_, _09186_, _09184_);
  nand (_09188_, _09187_, _09183_);
  nand (_09189_, _09188_, _08668_);
  nand (_09190_, _08676_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_09191_, _08676_, _08495_);
  and (_09192_, _09191_, _08685_);
  nand (_09193_, _09192_, _09190_);
  nand (_09194_, _08676_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_09195_, _08676_, _08487_);
  and (_09196_, _09195_, _08684_);
  nand (_09197_, _09196_, _09194_);
  nand (_09198_, _09197_, _09193_);
  nand (_09199_, _09198_, _08696_);
  nand (_09200_, _09199_, _09189_);
  nand (_09201_, _09200_, _08656_);
  nand (_09202_, _09201_, _09179_);
  or (_09203_, _08676_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_09204_, _08686_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_09205_, _09204_, _08685_);
  and (_09206_, _09205_, _09203_);
  or (_09207_, _08686_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_09208_, _08676_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_09209_, _09208_, _08684_);
  and (_09210_, _09209_, _09207_);
  nor (_09211_, _09210_, _09206_);
  nand (_09212_, _09211_, _08668_);
  or (_09213_, _08676_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_09214_, _08686_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_09215_, _09214_, _08685_);
  and (_09216_, _09215_, _09213_);
  or (_09217_, _08686_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_09218_, _08676_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_09219_, _09218_, _08684_);
  and (_09220_, _09219_, _09217_);
  nor (_09221_, _09220_, _09216_);
  nand (_09222_, _09221_, _08696_);
  nand (_09223_, _09222_, _09212_);
  nand (_09224_, _09223_, _08657_);
  or (_09225_, _08676_, _07528_);
  nand (_09226_, _08676_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_09227_, _09226_, _08685_);
  nand (_09228_, _09227_, _09225_);
  nand (_09229_, _08676_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_09230_, _08676_, _07532_);
  and (_09231_, _09230_, _08684_);
  nand (_09232_, _09231_, _09229_);
  nand (_09233_, _09232_, _09228_);
  nand (_09234_, _09233_, _08668_);
  nand (_09235_, _08676_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_09236_, _08676_, _07548_);
  and (_09237_, _09236_, _08685_);
  nand (_09238_, _09237_, _09235_);
  nand (_09239_, _08676_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_09240_, _08676_, _07540_);
  and (_09241_, _09240_, _08684_);
  nand (_09242_, _09241_, _09239_);
  nand (_09243_, _09242_, _09238_);
  nand (_09244_, _09243_, _08696_);
  nand (_09245_, _09244_, _09234_);
  nand (_09246_, _09245_, _08656_);
  and (_09247_, _09246_, _09224_);
  not (_09248_, _09247_);
  and (_09249_, _08684_, _07736_);
  nor (_09250_, _08684_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_09251_, _09250_, _09249_);
  and (_09252_, _09251_, _08676_);
  and (_09253_, _08684_, _07734_);
  nor (_09254_, _08684_, \oc8051_golden_model_1.IRAM[9] [2]);
  or (_09255_, _09254_, _09253_);
  and (_09256_, _09255_, _08686_);
  or (_09257_, _09256_, _09252_);
  nand (_09258_, _09257_, _08668_);
  and (_09259_, _08684_, _07748_);
  nor (_09260_, _08684_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_09261_, _09260_, _09259_);
  and (_09262_, _09261_, _08676_);
  and (_09263_, _08684_, _07746_);
  nor (_09264_, _08684_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_09265_, _09264_, _09263_);
  and (_09266_, _09265_, _08686_);
  or (_09267_, _09266_, _09262_);
  nand (_09268_, _09267_, _08696_);
  nand (_09269_, _09268_, _09258_);
  nand (_09270_, _09269_, _08657_);
  or (_09271_, _08676_, _07706_);
  nand (_09272_, _08676_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_09273_, _09272_, _08685_);
  nand (_09274_, _09273_, _09271_);
  nand (_09275_, _08676_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_09276_, _08676_, _07710_);
  and (_09277_, _09276_, _08684_);
  nand (_09278_, _09277_, _09275_);
  nand (_09279_, _09278_, _09274_);
  nand (_09280_, _09279_, _08668_);
  nand (_09281_, _08676_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_09282_, _08676_, _07726_);
  and (_09283_, _09282_, _08685_);
  nand (_09284_, _09283_, _09281_);
  nand (_09285_, _08676_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_09286_, _08676_, _07718_);
  and (_09287_, _09286_, _08684_);
  nand (_09288_, _09287_, _09285_);
  nand (_09289_, _09288_, _09284_);
  nand (_09290_, _09289_, _08696_);
  nand (_09291_, _09290_, _09280_);
  nand (_09292_, _09291_, _08656_);
  and (_09293_, _09292_, _09270_);
  not (_09294_, _09293_);
  or (_09295_, _08676_, \oc8051_golden_model_1.IRAM[9] [1]);
  or (_09296_, _08686_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_09297_, _09296_, _08685_);
  and (_09298_, _09297_, _09295_);
  or (_09299_, _08686_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_09300_, _08676_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_09301_, _09300_, _08684_);
  and (_09302_, _09301_, _09299_);
  nor (_09303_, _09302_, _09298_);
  nand (_09304_, _09303_, _08668_);
  or (_09305_, _08676_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_09306_, _08686_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_09307_, _09306_, _08685_);
  and (_09308_, _09307_, _09305_);
  or (_09309_, _08686_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_09310_, _08676_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_09311_, _09310_, _08684_);
  and (_09312_, _09311_, _09309_);
  nor (_09313_, _09312_, _09308_);
  nand (_09314_, _09313_, _08696_);
  nand (_09315_, _09314_, _09304_);
  nand (_09316_, _09315_, _08657_);
  or (_09317_, _08676_, _07284_);
  nand (_09318_, _08676_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_09319_, _09318_, _08685_);
  nand (_09320_, _09319_, _09317_);
  nand (_09321_, _08676_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_09322_, _08676_, _07288_);
  and (_09323_, _09322_, _08684_);
  nand (_09324_, _09323_, _09321_);
  nand (_09325_, _09324_, _09320_);
  nand (_09326_, _09325_, _08668_);
  nand (_09327_, _08676_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_09328_, _08676_, _07304_);
  and (_09329_, _09328_, _08685_);
  nand (_09330_, _09329_, _09327_);
  nand (_09331_, _08676_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_09332_, _08676_, _07296_);
  and (_09333_, _09332_, _08684_);
  nand (_09334_, _09333_, _09331_);
  nand (_09335_, _09334_, _09330_);
  nand (_09336_, _09335_, _08696_);
  nand (_09337_, _09336_, _09326_);
  nand (_09338_, _09337_, _08656_);
  and (_09339_, _09338_, _09316_);
  and (_09340_, _08684_, _07111_);
  nor (_09341_, _08684_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_09342_, _09341_, _09340_);
  and (_09343_, _09342_, _08676_);
  and (_09344_, _08684_, _07109_);
  nor (_09345_, _08684_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_09346_, _09345_, _09344_);
  and (_09347_, _09346_, _08686_);
  or (_09348_, _09347_, _09343_);
  nand (_09349_, _09348_, _08668_);
  and (_09350_, _08684_, _07123_);
  nor (_09351_, _08684_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_09352_, _09351_, _09350_);
  and (_09353_, _09352_, _08676_);
  and (_09354_, _08684_, _07121_);
  nor (_09355_, _08684_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_09356_, _09355_, _09354_);
  and (_09357_, _09356_, _08686_);
  or (_09358_, _09357_, _09353_);
  nand (_09359_, _09358_, _08696_);
  nand (_09360_, _09359_, _09349_);
  nand (_09361_, _09360_, _08657_);
  or (_09362_, _08676_, _07077_);
  nand (_09363_, _08676_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_09364_, _09363_, _08685_);
  nand (_09365_, _09364_, _09362_);
  nand (_09366_, _08676_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_09367_, _08676_, _07082_);
  and (_09368_, _09367_, _08684_);
  nand (_09369_, _09368_, _09366_);
  nand (_09370_, _09369_, _09365_);
  nand (_09371_, _09370_, _08668_);
  nand (_09372_, _08676_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_09373_, _08676_, _07100_);
  and (_09374_, _09373_, _08685_);
  nand (_09375_, _09374_, _09372_);
  nand (_09376_, _08676_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_09377_, _08676_, _07092_);
  and (_09378_, _09377_, _08684_);
  nand (_09379_, _09378_, _09376_);
  nand (_09380_, _09379_, _09375_);
  nand (_09381_, _09380_, _08696_);
  nand (_09382_, _09381_, _09371_);
  nand (_09383_, _09382_, _08656_);
  and (_09384_, _09383_, _09361_);
  nor (_09385_, _09384_, _09339_);
  and (_09386_, _09385_, _09294_);
  and (_09387_, _09386_, _09248_);
  and (_09388_, _09387_, _09202_);
  and (_09389_, _09388_, _09157_);
  and (_09390_, _09389_, _09112_);
  nor (_09391_, _09390_, _09067_);
  and (_09392_, _09390_, _09067_);
  or (_09393_, _09392_, _07244_);
  or (_09394_, _09393_, _09391_);
  and (_09395_, _09394_, _09066_);
  and (_09396_, _09395_, _09065_);
  and (_09397_, _08637_, _07241_);
  or (_09398_, _09397_, _06432_);
  or (_09399_, _09398_, _09396_);
  and (_09400_, _05625_, \oc8051_golden_model_1.PC [2]);
  and (_09401_, _09400_, \oc8051_golden_model_1.PC [3]);
  and (_09402_, _09401_, _08740_);
  and (_09403_, _09402_, \oc8051_golden_model_1.PC [7]);
  nor (_09404_, _09402_, \oc8051_golden_model_1.PC [7]);
  nor (_09405_, _09404_, _09403_);
  or (_09406_, _09405_, _06433_);
  and (_09407_, _09406_, _09399_);
  or (_09408_, _09407_, _05991_);
  and (_09409_, _08773_, _05991_);
  nor (_09410_, _09409_, _07251_);
  and (_09411_, _09410_, _09408_);
  and (_09412_, _08622_, _07251_);
  and (_09413_, _05766_, _05879_);
  nor (_09414_, _09413_, _09412_);
  not (_09415_, _09414_);
  nor (_09416_, _09415_, _09411_);
  not (_09417_, _09413_);
  and (_09418_, _08124_, _08102_);
  and (_09419_, _08227_, _08204_);
  and (_09420_, _08524_, _08502_);
  and (_09421_, _07577_, _07555_);
  and (_09422_, _07333_, _07311_);
  and (_09423_, _09422_, _07135_);
  and (_09424_, _09423_, _08662_);
  and (_09425_, _09424_, _09421_);
  and (_09426_, _09425_, _09420_);
  and (_09427_, _09426_, _09419_);
  and (_09428_, _09427_, _09418_);
  nor (_09429_, _09428_, _08023_);
  and (_09430_, _09428_, _08023_);
  or (_09431_, _09430_, _09429_);
  nor (_09432_, _09431_, _09417_);
  nor (_09433_, _09432_, _09416_);
  nor (_09434_, _09433_, _07261_);
  and (_09435_, _09111_, _09089_);
  and (_09436_, _09156_, _09134_);
  and (_09437_, _09201_, _09179_);
  and (_09438_, _09384_, _09339_);
  and (_09439_, _09438_, _09293_);
  and (_09440_, _09439_, _09247_);
  and (_09441_, _09440_, _09437_);
  and (_09442_, _09441_, _09436_);
  and (_09443_, _09442_, _09435_);
  nor (_09444_, _09443_, _09067_);
  and (_09445_, _09443_, _09067_);
  or (_09446_, _09445_, _09444_);
  nor (_09447_, _09446_, _07439_);
  nor (_09448_, _09447_, _07265_);
  not (_09449_, _09448_);
  nor (_09450_, _09449_, _09434_);
  nor (_09451_, _09450_, _08535_);
  nor (_09452_, _09451_, _07523_);
  or (_09453_, _09452_, _07868_);
  and (_09454_, _09453_, _07867_);
  not (_09455_, \oc8051_golden_model_1.PC [15]);
  and (_09456_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and (_09457_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_09458_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_09459_, _09458_, _09457_);
  and (_09460_, _09459_, _09403_);
  and (_09461_, _09460_, _09456_);
  and (_09462_, _09461_, \oc8051_golden_model_1.PC [14]);
  and (_09463_, _09462_, _09455_);
  nor (_09464_, _09462_, _09455_);
  or (_09465_, _09464_, _09463_);
  and (_09466_, _09465_, _06432_);
  and (_09467_, _09459_, _08742_);
  and (_09468_, _09467_, _09456_);
  and (_09469_, _09468_, \oc8051_golden_model_1.PC [14]);
  and (_09470_, _09469_, _09455_);
  nor (_09471_, _09469_, _09455_);
  or (_09472_, _09471_, _09470_);
  not (_09473_, _09472_);
  nor (_09474_, _09473_, _06432_);
  or (_09475_, _09474_, _09466_);
  and (_09476_, _09475_, _07862_);
  and (_09477_, _09476_, _07865_);
  or (_40310_, _09477_, _09454_);
  not (_09478_, \oc8051_golden_model_1.B [7]);
  nor (_09479_, _01320_, _09478_);
  and (_09480_, _06418_, _05971_);
  not (_09481_, _09480_);
  nor (_09482_, _07933_, _09478_);
  and (_09483_, _09004_, _07933_);
  or (_09484_, _09483_, _09482_);
  and (_09485_, _09484_, _05972_);
  not (_09486_, _06258_);
  and (_09487_, _08536_, _07933_);
  or (_09489_, _09487_, _09482_);
  or (_09490_, _09489_, _06260_);
  nor (_09491_, _08594_, _09478_);
  and (_09492_, _08622_, _08594_);
  or (_09493_, _09492_, _09491_);
  and (_09494_, _09493_, _06277_);
  and (_09495_, _08637_, _07933_);
  or (_09496_, _09495_, _09482_);
  or (_09497_, _09496_, _06286_);
  and (_09498_, _07933_, \oc8051_golden_model_1.ACC [7]);
  or (_09499_, _09498_, _09482_);
  and (_09500_, _09499_, _07143_);
  nor (_09501_, _07143_, _09478_);
  or (_09502_, _09501_, _06285_);
  or (_09503_, _09502_, _09500_);
  and (_09504_, _09503_, _06282_);
  and (_09505_, _09504_, _09497_);
  and (_09506_, _08626_, _08594_);
  or (_09507_, _09506_, _09491_);
  and (_09508_, _09507_, _06281_);
  or (_09510_, _09508_, _06354_);
  or (_09511_, _09510_, _09505_);
  or (_09512_, _09489_, _07169_);
  and (_09513_, _09512_, _09511_);
  or (_09514_, _09513_, _06345_);
  or (_09515_, _09499_, _06346_);
  and (_09516_, _09515_, _06278_);
  and (_09517_, _09516_, _09514_);
  or (_09518_, _09517_, _09494_);
  and (_09519_, _09518_, _06271_);
  and (_09520_, _06418_, _06336_);
  or (_09521_, _09491_, _08768_);
  and (_09522_, _09521_, _06270_);
  and (_09523_, _09522_, _09507_);
  or (_09524_, _09523_, _09520_);
  or (_09525_, _09524_, _09519_);
  and (_09526_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_09527_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_09528_, _09527_, _09526_);
  and (_09529_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and (_09530_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_09531_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_09532_, _09531_, _09530_);
  nor (_09533_, _09532_, _09528_);
  and (_09534_, _09533_, _09529_);
  nor (_09535_, _09534_, _09528_);
  and (_09536_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_09537_, _09536_, _09531_);
  and (_09538_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_09539_, _09538_, _09526_);
  nor (_09540_, _09539_, _09537_);
  not (_09541_, _09540_);
  nor (_09542_, _09541_, _09535_);
  and (_09543_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_09544_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and (_09545_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and (_09546_, _09545_, _09544_);
  nor (_09547_, _09545_, _09544_);
  nor (_09548_, _09547_, _09546_);
  and (_09549_, _09548_, _09543_);
  nor (_09550_, _09548_, _09543_);
  nor (_09551_, _09550_, _09549_);
  and (_09552_, _09541_, _09535_);
  nor (_09553_, _09552_, _09542_);
  and (_09554_, _09553_, _09551_);
  nor (_09555_, _09554_, _09542_);
  not (_09556_, _09531_);
  and (_09557_, _09536_, _09556_);
  and (_09558_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and (_09559_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_09560_, _09559_, _09544_);
  and (_09561_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  and (_09562_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_09563_, _09562_, _09561_);
  nor (_09564_, _09563_, _09560_);
  and (_09565_, _09564_, _09558_);
  nor (_09566_, _09564_, _09558_);
  nor (_09567_, _09566_, _09565_);
  and (_09568_, _09567_, _09557_);
  nor (_09569_, _09567_, _09557_);
  nor (_09570_, _09569_, _09568_);
  not (_09571_, _09570_);
  nor (_09572_, _09571_, _09555_);
  and (_09573_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_09574_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and (_09575_, _09574_, _09573_);
  nor (_09576_, _09549_, _09546_);
  and (_09577_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and (_09578_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_09579_, _09578_, _09577_);
  nor (_09580_, _09578_, _09577_);
  nor (_09581_, _09580_, _09579_);
  not (_09582_, _09581_);
  nor (_09583_, _09582_, _09576_);
  and (_09584_, _09582_, _09576_);
  nor (_09585_, _09584_, _09583_);
  and (_09586_, _09585_, _09575_);
  nor (_09587_, _09585_, _09575_);
  nor (_09588_, _09587_, _09586_);
  and (_09589_, _09571_, _09555_);
  nor (_09590_, _09589_, _09572_);
  and (_09591_, _09590_, _09588_);
  nor (_09592_, _09591_, _09572_);
  nor (_09593_, _09565_, _09560_);
  and (_09594_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and (_09595_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and (_09596_, _09595_, _09594_);
  nor (_09597_, _09595_, _09594_);
  nor (_09598_, _09597_, _09596_);
  not (_09599_, _09598_);
  nor (_09600_, _09599_, _09593_);
  and (_09601_, _09599_, _09593_);
  nor (_09602_, _09601_, _09600_);
  and (_09603_, _09602_, _09579_);
  nor (_09604_, _09602_, _09579_);
  nor (_09605_, _09604_, _09603_);
  nor (_09606_, _09568_, _09537_);
  and (_09607_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  and (_09608_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_09609_, _09608_, _09559_);
  nor (_09610_, _09608_, _09559_);
  nor (_09611_, _09610_, _09609_);
  and (_09612_, _09611_, _09607_);
  nor (_09613_, _09611_, _09607_);
  nor (_09614_, _09613_, _09612_);
  not (_09615_, _09614_);
  nor (_09616_, _09615_, _09606_);
  and (_09617_, _09615_, _09606_);
  nor (_09618_, _09617_, _09616_);
  and (_09619_, _09618_, _09605_);
  nor (_09620_, _09618_, _09605_);
  nor (_09621_, _09620_, _09619_);
  not (_09622_, _09621_);
  nor (_09623_, _09622_, _09592_);
  nor (_09624_, _09586_, _09583_);
  not (_09625_, _09624_);
  and (_09626_, _09622_, _09592_);
  nor (_09627_, _09626_, _09623_);
  and (_09628_, _09627_, _09625_);
  nor (_09629_, _09628_, _09623_);
  nor (_09630_, _09603_, _09600_);
  not (_09631_, _09630_);
  nor (_09632_, _09619_, _09616_);
  not (_09633_, _09632_);
  and (_09634_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_09635_, _09634_, _09559_);
  and (_09636_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_09637_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_09638_, _09637_, _09636_);
  nor (_09639_, _09638_, _09635_);
  nor (_09640_, _09612_, _09609_);
  and (_09641_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and (_09642_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and (_09643_, _09642_, _09641_);
  nor (_09644_, _09642_, _09641_);
  nor (_09645_, _09644_, _09643_);
  not (_09646_, _09645_);
  nor (_09647_, _09646_, _09640_);
  and (_09648_, _09646_, _09640_);
  nor (_09649_, _09648_, _09647_);
  and (_09650_, _09649_, _09596_);
  nor (_09651_, _09649_, _09596_);
  nor (_09652_, _09651_, _09650_);
  and (_09653_, _09652_, _09639_);
  nor (_09654_, _09652_, _09639_);
  nor (_09655_, _09654_, _09653_);
  and (_09656_, _09655_, _09633_);
  nor (_09657_, _09655_, _09633_);
  nor (_09658_, _09657_, _09656_);
  and (_09659_, _09658_, _09631_);
  nor (_09660_, _09658_, _09631_);
  nor (_09661_, _09660_, _09659_);
  not (_09662_, _09661_);
  nor (_09663_, _09662_, _09629_);
  nor (_09665_, _09659_, _09656_);
  nor (_09666_, _09650_, _09647_);
  not (_09668_, _09666_);
  and (_09669_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and (_09671_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_09672_, _09671_, _09669_);
  nor (_09674_, _09671_, _09669_);
  nor (_09675_, _09674_, _09672_);
  and (_09677_, _09675_, _09635_);
  nor (_09678_, _09675_, _09635_);
  nor (_09680_, _09678_, _09677_);
  and (_09681_, _09680_, _09643_);
  nor (_09683_, _09680_, _09643_);
  nor (_09684_, _09683_, _09681_);
  and (_09686_, _09684_, _09634_);
  nor (_09687_, _09684_, _09634_);
  nor (_09689_, _09687_, _09686_);
  and (_09690_, _09689_, _09653_);
  nor (_09692_, _09689_, _09653_);
  nor (_09693_, _09692_, _09690_);
  and (_09695_, _09693_, _09668_);
  nor (_09696_, _09693_, _09668_);
  nor (_09698_, _09696_, _09695_);
  not (_09699_, _09698_);
  nor (_09701_, _09699_, _09665_);
  and (_09702_, _09699_, _09665_);
  nor (_09703_, _09702_, _09701_);
  and (_09704_, _09703_, _09663_);
  nor (_09705_, _09695_, _09690_);
  nor (_09706_, _09681_, _09677_);
  not (_09707_, _09706_);
  and (_09708_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and (_09709_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_09710_, _09709_, _09708_);
  nor (_09711_, _09709_, _09708_);
  nor (_09712_, _09711_, _09710_);
  and (_09713_, _09712_, _09672_);
  nor (_09714_, _09712_, _09672_);
  nor (_09715_, _09714_, _09713_);
  and (_09716_, _09715_, _09686_);
  nor (_09717_, _09715_, _09686_);
  nor (_09718_, _09717_, _09716_);
  and (_09719_, _09718_, _09707_);
  nor (_09720_, _09718_, _09707_);
  nor (_09721_, _09720_, _09719_);
  not (_09722_, _09721_);
  nor (_09723_, _09722_, _09705_);
  and (_09724_, _09722_, _09705_);
  nor (_09725_, _09724_, _09723_);
  and (_09726_, _09725_, _09701_);
  nor (_09727_, _09725_, _09701_);
  nor (_09728_, _09727_, _09726_);
  and (_09729_, _09728_, _09704_);
  nor (_09730_, _09728_, _09704_);
  nor (_09731_, _09730_, _09729_);
  and (_09732_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and (_09733_, _09732_, _09531_);
  and (_09734_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and (_09735_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor (_09736_, _09735_, _09527_);
  nor (_09737_, _09736_, _09733_);
  and (_09738_, _09737_, _09734_);
  nor (_09739_, _09738_, _09733_);
  not (_09740_, _09739_);
  nor (_09741_, _09533_, _09529_);
  nor (_09742_, _09741_, _09534_);
  and (_09743_, _09742_, _09740_);
  and (_09744_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_09745_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and (_09746_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_09747_, _09746_, _09745_);
  nor (_09748_, _09746_, _09745_);
  nor (_09749_, _09748_, _09747_);
  and (_09750_, _09749_, _09744_);
  nor (_09751_, _09749_, _09744_);
  nor (_09752_, _09751_, _09750_);
  nor (_09753_, _09742_, _09740_);
  nor (_09754_, _09753_, _09743_);
  and (_09755_, _09754_, _09752_);
  nor (_09756_, _09755_, _09743_);
  nor (_09757_, _09553_, _09551_);
  nor (_09758_, _09757_, _09554_);
  not (_09760_, _09758_);
  nor (_09762_, _09760_, _09756_);
  and (_09763_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_09765_, _09763_, _09574_);
  nor (_09766_, _09750_, _09747_);
  nor (_09768_, _09574_, _09573_);
  nor (_09769_, _09768_, _09575_);
  not (_09771_, _09769_);
  nor (_09772_, _09771_, _09766_);
  and (_09774_, _09771_, _09766_);
  nor (_09775_, _09774_, _09772_);
  and (_09777_, _09775_, _09765_);
  nor (_09778_, _09775_, _09765_);
  nor (_09780_, _09778_, _09777_);
  and (_09781_, _09760_, _09756_);
  nor (_09783_, _09781_, _09762_);
  and (_09784_, _09783_, _09780_);
  nor (_09786_, _09784_, _09762_);
  nor (_09787_, _09590_, _09588_);
  nor (_09789_, _09787_, _09591_);
  not (_09790_, _09789_);
  nor (_09792_, _09790_, _09786_);
  nor (_09793_, _09777_, _09772_);
  not (_09795_, _09793_);
  and (_09796_, _09790_, _09786_);
  nor (_09797_, _09796_, _09792_);
  and (_09798_, _09797_, _09795_);
  nor (_09799_, _09798_, _09792_);
  nor (_09800_, _09627_, _09625_);
  nor (_09801_, _09800_, _09628_);
  not (_09802_, _09801_);
  nor (_09803_, _09802_, _09799_);
  and (_09804_, _09662_, _09629_);
  nor (_09805_, _09804_, _09663_);
  and (_09806_, _09805_, _09803_);
  nor (_09807_, _09703_, _09663_);
  nor (_09808_, _09807_, _09704_);
  nand (_09809_, _09808_, _09806_);
  and (_09810_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and (_09811_, _09810_, _09732_);
  and (_09812_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_09813_, _09810_, _09732_);
  nor (_09814_, _09813_, _09811_);
  and (_09815_, _09814_, _09812_);
  nor (_09816_, _09815_, _09811_);
  not (_09817_, _09816_);
  nor (_09818_, _09737_, _09734_);
  nor (_09819_, _09818_, _09738_);
  and (_09820_, _09819_, _09817_);
  and (_09821_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and (_09822_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_09823_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_09824_, _09823_, _09822_);
  nor (_09825_, _09823_, _09822_);
  nor (_09826_, _09825_, _09824_);
  and (_09827_, _09826_, _09821_);
  nor (_09828_, _09826_, _09821_);
  nor (_09829_, _09828_, _09827_);
  nor (_09830_, _09819_, _09817_);
  nor (_09831_, _09830_, _09820_);
  and (_09832_, _09831_, _09829_);
  nor (_09833_, _09832_, _09820_);
  not (_09834_, _09833_);
  nor (_09835_, _09754_, _09752_);
  nor (_09836_, _09835_, _09755_);
  and (_09837_, _09836_, _09834_);
  nor (_09838_, _09827_, _09824_);
  and (_09839_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and (_09840_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor (_09841_, _09840_, _09839_);
  nor (_09842_, _09841_, _09765_);
  not (_09843_, _09842_);
  nor (_09844_, _09843_, _09838_);
  and (_09845_, _09843_, _09838_);
  nor (_09846_, _09845_, _09844_);
  nor (_09847_, _09836_, _09834_);
  nor (_09848_, _09847_, _09837_);
  and (_09849_, _09848_, _09846_);
  nor (_09850_, _09849_, _09837_);
  nor (_09851_, _09783_, _09780_);
  nor (_09852_, _09851_, _09784_);
  not (_09853_, _09852_);
  nor (_09854_, _09853_, _09850_);
  and (_09855_, _09853_, _09850_);
  nor (_09856_, _09855_, _09854_);
  and (_09857_, _09856_, _09844_);
  nor (_09858_, _09857_, _09854_);
  nor (_09859_, _09797_, _09795_);
  nor (_09860_, _09859_, _09798_);
  not (_09861_, _09860_);
  nor (_09862_, _09861_, _09858_);
  and (_09863_, _09802_, _09799_);
  nor (_09864_, _09863_, _09803_);
  and (_09865_, _09864_, _09862_);
  nor (_09866_, _09805_, _09803_);
  nor (_09867_, _09866_, _09806_);
  and (_09868_, _09867_, _09865_);
  nor (_09869_, _09867_, _09865_);
  nor (_09870_, _09869_, _09868_);
  and (_09871_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and (_09872_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_09873_, _09872_, _09871_);
  and (_09874_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_09875_, _09872_, _09871_);
  nor (_09876_, _09875_, _09873_);
  and (_09877_, _09876_, _09874_);
  nor (_09878_, _09877_, _09873_);
  not (_09879_, _09878_);
  nor (_09880_, _09814_, _09812_);
  nor (_09881_, _09880_, _09815_);
  and (_09882_, _09881_, _09879_);
  and (_09883_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_09884_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_09885_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and (_09886_, _09885_, _09884_);
  nor (_09887_, _09885_, _09884_);
  nor (_09888_, _09887_, _09886_);
  and (_09889_, _09888_, _09883_);
  nor (_09890_, _09888_, _09883_);
  nor (_09891_, _09890_, _09889_);
  nor (_09892_, _09881_, _09879_);
  nor (_09893_, _09892_, _09882_);
  and (_09894_, _09893_, _09891_);
  nor (_09895_, _09894_, _09882_);
  not (_09896_, _09895_);
  nor (_09897_, _09831_, _09829_);
  nor (_09898_, _09897_, _09832_);
  and (_09899_, _09898_, _09896_);
  not (_09900_, _09763_);
  nor (_09901_, _09889_, _09886_);
  nor (_09902_, _09901_, _09900_);
  and (_09903_, _09901_, _09900_);
  nor (_09904_, _09903_, _09902_);
  nor (_09905_, _09898_, _09896_);
  nor (_09906_, _09905_, _09899_);
  and (_09907_, _09906_, _09904_);
  nor (_09908_, _09907_, _09899_);
  not (_09909_, _09908_);
  nor (_09910_, _09848_, _09846_);
  nor (_09911_, _09910_, _09849_);
  and (_09912_, _09911_, _09909_);
  nor (_09913_, _09911_, _09909_);
  nor (_09914_, _09913_, _09912_);
  and (_09915_, _09914_, _09902_);
  nor (_09916_, _09915_, _09912_);
  nor (_09917_, _09856_, _09844_);
  nor (_09918_, _09917_, _09857_);
  not (_09919_, _09918_);
  nor (_09920_, _09919_, _09916_);
  and (_09921_, _09861_, _09858_);
  nor (_09922_, _09921_, _09862_);
  and (_09923_, _09922_, _09920_);
  nor (_09924_, _09864_, _09862_);
  nor (_09925_, _09924_, _09865_);
  nand (_09926_, _09925_, _09923_);
  or (_09927_, _09925_, _09923_);
  and (_09928_, _09927_, _09926_);
  and (_09929_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_09930_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_09931_, _09930_, _09929_);
  and (_09932_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor (_09933_, _09930_, _09929_);
  nor (_09934_, _09933_, _09931_);
  and (_09935_, _09934_, _09932_);
  nor (_09936_, _09935_, _09931_);
  not (_09937_, _09936_);
  nor (_09938_, _09876_, _09874_);
  nor (_09939_, _09938_, _09877_);
  and (_09940_, _09939_, _09937_);
  and (_09941_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_09942_, _09941_, _09885_);
  and (_09943_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and (_09944_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_09945_, _09944_, _09943_);
  nor (_09946_, _09945_, _09942_);
  nor (_09947_, _09939_, _09937_);
  nor (_09948_, _09947_, _09940_);
  and (_09949_, _09948_, _09946_);
  nor (_09950_, _09949_, _09940_);
  not (_09951_, _09950_);
  nor (_09952_, _09893_, _09891_);
  nor (_09953_, _09952_, _09894_);
  and (_09954_, _09953_, _09951_);
  nor (_09955_, _09953_, _09951_);
  nor (_09956_, _09955_, _09954_);
  and (_09957_, _09956_, _09942_);
  nor (_09958_, _09957_, _09954_);
  not (_09959_, _09958_);
  nor (_09960_, _09906_, _09904_);
  nor (_09961_, _09960_, _09907_);
  and (_09962_, _09961_, _09959_);
  nor (_09963_, _09914_, _09902_);
  nor (_09964_, _09963_, _09915_);
  and (_09965_, _09964_, _09962_);
  and (_09966_, _09919_, _09916_);
  nor (_09967_, _09966_, _09920_);
  and (_09968_, _09967_, _09965_);
  nor (_09969_, _09922_, _09920_);
  nor (_09970_, _09969_, _09923_);
  nor (_09971_, _09970_, _09968_);
  and (_09972_, _09970_, _09968_);
  not (_09973_, _09972_);
  and (_09974_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_09975_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and (_09976_, _09975_, _09974_);
  and (_09977_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_09978_, _09975_, _09974_);
  nor (_09979_, _09978_, _09976_);
  and (_09980_, _09979_, _09977_);
  nor (_09981_, _09980_, _09976_);
  not (_09982_, _09981_);
  nor (_09983_, _09934_, _09932_);
  nor (_09984_, _09983_, _09935_);
  and (_09985_, _09984_, _09982_);
  nor (_09986_, _09984_, _09982_);
  nor (_09987_, _09986_, _09985_);
  and (_09988_, _09987_, _09941_);
  nor (_09989_, _09988_, _09985_);
  not (_09990_, _09989_);
  nor (_09991_, _09948_, _09946_);
  nor (_09992_, _09991_, _09949_);
  and (_09993_, _09992_, _09990_);
  nor (_09994_, _09956_, _09942_);
  nor (_09995_, _09994_, _09957_);
  and (_09996_, _09995_, _09993_);
  nor (_09997_, _09961_, _09959_);
  nor (_09998_, _09997_, _09962_);
  and (_09999_, _09998_, _09996_);
  nor (_10000_, _09964_, _09962_);
  nor (_10001_, _10000_, _09965_);
  and (_10002_, _10001_, _09999_);
  nor (_10003_, _09967_, _09965_);
  nor (_10004_, _10003_, _09968_);
  and (_10005_, _10004_, _10002_);
  and (_10006_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and (_10007_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and (_10008_, _10007_, _10006_);
  nor (_10009_, _09979_, _09977_);
  nor (_10010_, _10009_, _09980_);
  and (_10011_, _10010_, _10008_);
  nor (_10012_, _09987_, _09941_);
  nor (_10013_, _10012_, _09988_);
  and (_10014_, _10013_, _10011_);
  nor (_10015_, _09992_, _09990_);
  nor (_10016_, _10015_, _09993_);
  and (_10017_, _10016_, _10014_);
  nor (_10018_, _09995_, _09993_);
  nor (_10019_, _10018_, _09996_);
  and (_10020_, _10019_, _10017_);
  nor (_10021_, _09998_, _09996_);
  nor (_10022_, _10021_, _09999_);
  and (_10023_, _10022_, _10020_);
  nor (_10024_, _10001_, _09999_);
  nor (_10025_, _10024_, _10002_);
  and (_10026_, _10025_, _10023_);
  nor (_10027_, _10004_, _10002_);
  nor (_10028_, _10027_, _10005_);
  and (_10029_, _10028_, _10026_);
  nor (_10030_, _10029_, _10005_);
  and (_10031_, _10030_, _09973_);
  nor (_10032_, _10031_, _09971_);
  nand (_10033_, _10032_, _09928_);
  and (_10034_, _10033_, _09926_);
  not (_10035_, _10034_);
  and (_10036_, _10035_, _09870_);
  or (_10037_, _10036_, _09868_);
  or (_10038_, _09808_, _09806_);
  and (_10039_, _10038_, _09809_);
  nand (_10040_, _10039_, _10037_);
  and (_10041_, _10040_, _09809_);
  not (_10042_, _10041_);
  and (_10043_, _10042_, _09731_);
  or (_10044_, _10043_, _09729_);
  and (_10045_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not (_10046_, _10045_);
  nor (_10047_, _10046_, _09671_);
  nor (_10048_, _10047_, _09713_);
  nor (_10049_, _09719_, _09716_);
  nor (_10050_, _10049_, _10048_);
  and (_10051_, _10049_, _10048_);
  nor (_10052_, _10051_, _10050_);
  not (_10053_, _10052_);
  nor (_10054_, _09726_, _09723_);
  and (_10055_, _10054_, _10053_);
  nor (_10056_, _10054_, _10053_);
  nor (_10057_, _10056_, _10055_);
  and (_10058_, _10057_, _10044_);
  not (_10059_, _09520_);
  or (_10060_, _10050_, _09710_);
  or (_10061_, _10060_, _10056_);
  or (_10062_, _10061_, _10059_);
  or (_10063_, _10062_, _10058_);
  and (_10064_, _10063_, _06267_);
  and (_10065_, _10064_, _09525_);
  and (_10066_, _08789_, _08594_);
  or (_10067_, _10066_, _09491_);
  and (_10068_, _10067_, _06266_);
  or (_10069_, _10068_, _06259_);
  or (_10070_, _10069_, _10065_);
  and (_10071_, _10070_, _09490_);
  or (_10072_, _10071_, _09486_);
  and (_10073_, _08731_, _07933_);
  or (_10074_, _09482_, _06258_);
  or (_10075_, _10074_, _10073_);
  and (_10076_, _10075_, _06251_);
  and (_10077_, _10076_, _10072_);
  or (_10078_, _10077_, _09485_);
  and (_10079_, _10078_, _09481_);
  not (_10080_, _06399_);
  not (_10081_, \oc8051_golden_model_1.B [1]);
  nor (_10082_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_10083_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_10084_, _10083_, _10082_);
  and (_10085_, _10084_, _10081_);
  not (_10086_, \oc8051_golden_model_1.B [0]);
  and (_10087_, _10086_, \oc8051_golden_model_1.ACC [7]);
  nor (_10088_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_10089_, _10088_, _10087_);
  and (_10090_, _10089_, _10085_);
  not (_10091_, _10088_);
  and (_10092_, \oc8051_golden_model_1.B [0], _08737_);
  nor (_10093_, _10092_, _10091_);
  and (_10094_, _10093_, _10085_);
  or (_10095_, _10094_, _08737_);
  not (_10096_, \oc8051_golden_model_1.B [2]);
  not (_10097_, \oc8051_golden_model_1.B [3]);
  not (_10098_, \oc8051_golden_model_1.B [4]);
  not (_10099_, \oc8051_golden_model_1.B [5]);
  nor (_10100_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_10101_, _10100_, _10099_);
  and (_10102_, _10101_, _10098_);
  and (_10103_, _10102_, _10097_);
  and (_10104_, _10103_, _10096_);
  not (_10105_, \oc8051_golden_model_1.ACC [6]);
  and (_10106_, \oc8051_golden_model_1.B [0], _10105_);
  nor (_10107_, _10106_, _08737_);
  nor (_10108_, _10107_, _10081_);
  not (_10109_, _10108_);
  and (_10110_, _10109_, _10104_);
  nor (_10111_, _10110_, _10095_);
  nor (_10112_, _10111_, _10090_);
  and (_10113_, _10110_, \oc8051_golden_model_1.B [0]);
  nor (_10114_, _10113_, _10105_);
  and (_10115_, _10114_, _10081_);
  nor (_10116_, _10114_, _10081_);
  nor (_10117_, _10116_, _10115_);
  nor (_10118_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor (_10119_, _10118_, _09732_);
  nor (_10120_, _10119_, \oc8051_golden_model_1.ACC [4]);
  and (_10121_, \oc8051_golden_model_1.ACC [4], _10086_);
  nor (_10122_, _10121_, \oc8051_golden_model_1.ACC [5]);
  not (_10123_, \oc8051_golden_model_1.ACC [4]);
  and (_10124_, _10123_, \oc8051_golden_model_1.B [0]);
  nor (_10125_, _10124_, _10122_);
  nor (_10126_, _10125_, _10120_);
  not (_10127_, _10126_);
  and (_10128_, _10127_, _10117_);
  nor (_10129_, _10112_, \oc8051_golden_model_1.B [2]);
  nor (_10130_, _10129_, _10115_);
  not (_10131_, _10130_);
  nor (_10132_, _10131_, _10128_);
  and (_10133_, \oc8051_golden_model_1.B [2], _08737_);
  nor (_10134_, _10133_, \oc8051_golden_model_1.B [7]);
  and (_10135_, _10134_, _10084_);
  not (_10136_, _10135_);
  nor (_10137_, _10136_, _10132_);
  nor (_10138_, _10137_, _10112_);
  nor (_10139_, _10138_, _10090_);
  and (_10140_, _10102_, \oc8051_golden_model_1.ACC [7]);
  nor (_10141_, _10140_, _10103_);
  nor (_10142_, _10127_, _10117_);
  nor (_10143_, _10142_, _10128_);
  not (_10144_, _10143_);
  and (_10145_, _10144_, _10137_);
  nor (_10146_, _10137_, _10114_);
  nor (_10147_, _10146_, _10145_);
  and (_10148_, _10147_, _10096_);
  nor (_10149_, _10147_, _10096_);
  nor (_10150_, _10149_, _10148_);
  not (_10151_, _10150_);
  not (_10152_, \oc8051_golden_model_1.ACC [5]);
  nor (_10153_, _10137_, _10152_);
  and (_10154_, _10137_, _10119_);
  or (_10155_, _10154_, _10153_);
  and (_10156_, _10155_, _10081_);
  nor (_10157_, _10155_, _10081_);
  nor (_10158_, _10157_, _10124_);
  nor (_10159_, _10158_, _10156_);
  nor (_10160_, _10159_, _10151_);
  nor (_10161_, _10139_, \oc8051_golden_model_1.B [3]);
  nor (_10162_, _10161_, _10148_);
  not (_10163_, _10162_);
  nor (_10164_, _10163_, _10160_);
  nor (_10165_, _10164_, _10141_);
  nor (_10166_, _10165_, _10139_);
  nor (_10167_, _10166_, _10090_);
  nor (_10168_, _10167_, \oc8051_golden_model_1.B [4]);
  not (_10169_, _10165_);
  and (_10170_, _10159_, _10151_);
  nor (_10171_, _10170_, _10160_);
  nor (_10172_, _10171_, _10169_);
  nor (_10173_, _10165_, _10147_);
  nor (_10174_, _10173_, _10172_);
  and (_10175_, _10174_, _10097_);
  nor (_10176_, _10174_, _10097_);
  nor (_10177_, _10176_, _10175_);
  not (_10178_, _10177_);
  nor (_10179_, _10165_, _10155_);
  nor (_10180_, _10157_, _10156_);
  and (_10181_, _10180_, _10124_);
  nor (_10182_, _10180_, _10124_);
  nor (_10183_, _10182_, _10181_);
  and (_10184_, _10183_, _10165_);
  or (_10185_, _10184_, _10179_);
  nor (_10186_, _10185_, \oc8051_golden_model_1.B [2]);
  and (_10187_, _10185_, \oc8051_golden_model_1.B [2]);
  nor (_10188_, _10124_, _10121_);
  and (_10189_, _10165_, _10188_);
  nor (_10190_, _10165_, \oc8051_golden_model_1.ACC [4]);
  nor (_10191_, _10190_, _10189_);
  and (_10192_, _10191_, _10081_);
  nor (_10193_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_10194_, _10193_, _09929_);
  nor (_10195_, _10194_, \oc8051_golden_model_1.ACC [2]);
  and (_10196_, _10086_, \oc8051_golden_model_1.ACC [2]);
  nor (_10197_, _10196_, \oc8051_golden_model_1.ACC [3]);
  not (_10198_, \oc8051_golden_model_1.ACC [2]);
  and (_10199_, \oc8051_golden_model_1.B [0], _10198_);
  nor (_10200_, _10199_, _10197_);
  nor (_10201_, _10200_, _10195_);
  not (_10202_, _10201_);
  nor (_10203_, _10191_, _10081_);
  nor (_10204_, _10203_, _10192_);
  and (_10205_, _10204_, _10202_);
  nor (_10206_, _10205_, _10192_);
  nor (_10207_, _10206_, _10187_);
  nor (_10208_, _10207_, _10186_);
  nor (_10209_, _10208_, _10178_);
  or (_10210_, _10209_, _10175_);
  nor (_10211_, _10210_, _10168_);
  and (_10212_, _10101_, \oc8051_golden_model_1.ACC [7]);
  or (_10213_, _10212_, _10102_);
  not (_10214_, _10213_);
  nor (_10215_, _10214_, _10211_);
  nor (_10216_, _10215_, _10167_);
  nor (_10217_, _10216_, _10090_);
  and (_10218_, _10100_, \oc8051_golden_model_1.ACC [7]);
  nor (_10219_, _10218_, _10101_);
  nor (_10220_, _10217_, \oc8051_golden_model_1.B [5]);
  and (_10221_, _10208_, _10178_);
  nor (_10222_, _10221_, _10209_);
  not (_10223_, _10222_);
  and (_10224_, _10223_, _10215_);
  nor (_10225_, _10215_, _10174_);
  nor (_10226_, _10225_, _10224_);
  and (_10227_, _10226_, _10098_);
  nor (_10228_, _10226_, _10098_);
  nor (_10229_, _10228_, _10227_);
  not (_10230_, _10229_);
  nor (_10231_, _10215_, _10185_);
  nor (_10232_, _10187_, _10186_);
  and (_10233_, _10232_, _10206_);
  nor (_10234_, _10232_, _10206_);
  nor (_10235_, _10234_, _10233_);
  not (_10236_, _10235_);
  and (_10237_, _10236_, _10215_);
  nor (_10238_, _10237_, _10231_);
  nor (_10239_, _10238_, \oc8051_golden_model_1.B [3]);
  and (_10240_, _10238_, \oc8051_golden_model_1.B [3]);
  nor (_10241_, _10204_, _10202_);
  nor (_10242_, _10241_, _10205_);
  not (_10243_, _10242_);
  and (_10244_, _10243_, _10215_);
  nor (_10245_, _10215_, _10191_);
  nor (_10246_, _10245_, _10244_);
  and (_10247_, _10246_, _10096_);
  not (_10248_, \oc8051_golden_model_1.ACC [3]);
  nor (_10249_, _10215_, _10248_);
  and (_10250_, _10215_, _10194_);
  or (_10251_, _10250_, _10249_);
  and (_10252_, _10251_, _10081_);
  nor (_10253_, _10251_, _10081_);
  nor (_10254_, _10253_, _10199_);
  nor (_10255_, _10254_, _10252_);
  nor (_10256_, _10246_, _10096_);
  nor (_10257_, _10256_, _10247_);
  not (_10258_, _10257_);
  nor (_10259_, _10258_, _10255_);
  nor (_10260_, _10259_, _10247_);
  nor (_10261_, _10260_, _10240_);
  nor (_10262_, _10261_, _10239_);
  nor (_10263_, _10262_, _10230_);
  or (_10264_, _10263_, _10227_);
  nor (_10265_, _10264_, _10220_);
  nor (_10266_, _10265_, _10219_);
  nor (_10267_, _10266_, _10217_);
  not (_10268_, _10266_);
  and (_10269_, _10262_, _10230_);
  nor (_10270_, _10269_, _10263_);
  nor (_10271_, _10270_, _10268_);
  nor (_10272_, _10266_, _10226_);
  nor (_10273_, _10272_, _10271_);
  and (_10274_, _10273_, _10099_);
  nor (_10275_, _10273_, _10099_);
  nor (_10276_, _10275_, _10274_);
  not (_10277_, _10276_);
  nor (_10278_, _10266_, _10238_);
  nor (_10279_, _10240_, _10239_);
  nor (_10280_, _10279_, _10260_);
  and (_10281_, _10279_, _10260_);
  or (_10282_, _10281_, _10280_);
  and (_10283_, _10282_, _10266_);
  or (_10284_, _10283_, _10278_);
  and (_10285_, _10284_, _10098_);
  nor (_10286_, _10284_, _10098_);
  and (_10287_, _10258_, _10255_);
  nor (_10288_, _10287_, _10259_);
  nor (_10289_, _10288_, _10268_);
  nor (_10290_, _10266_, _10246_);
  nor (_10291_, _10290_, _10289_);
  and (_10292_, _10291_, _10097_);
  nor (_10293_, _10253_, _10252_);
  nor (_10294_, _10293_, _10199_);
  and (_10295_, _10293_, _10199_);
  or (_10296_, _10295_, _10294_);
  nor (_10297_, _10296_, _10268_);
  nor (_10298_, _10266_, _10251_);
  nor (_10299_, _10298_, _10297_);
  and (_10300_, _10299_, _10096_);
  nor (_10301_, _10299_, _10096_);
  nor (_10302_, _10266_, \oc8051_golden_model_1.ACC [2]);
  nor (_10303_, _10199_, _10196_);
  and (_10304_, _10266_, _10303_);
  nor (_10305_, _10304_, _10302_);
  and (_10306_, _10305_, _10081_);
  and (_10307_, _06044_, \oc8051_golden_model_1.B [0]);
  not (_10308_, _10307_);
  nor (_10309_, _10305_, _10081_);
  nor (_10310_, _10309_, _10306_);
  and (_10311_, _10310_, _10308_);
  nor (_10312_, _10311_, _10306_);
  nor (_10313_, _10312_, _10301_);
  nor (_10314_, _10313_, _10300_);
  nor (_10315_, _10291_, _10097_);
  nor (_10316_, _10315_, _10292_);
  not (_10317_, _10316_);
  nor (_10318_, _10317_, _10314_);
  nor (_10319_, _10318_, _10292_);
  nor (_10320_, _10319_, _10286_);
  nor (_10321_, _10320_, _10285_);
  nor (_10322_, _10321_, _10277_);
  nor (_10323_, _10322_, _10274_);
  and (_10324_, \oc8051_golden_model_1.ACC [7], _09478_);
  nor (_10325_, _10324_, _10100_);
  nor (_10326_, _10325_, _10323_);
  not (_10327_, _10100_);
  nor (_10328_, _10267_, _10090_);
  nor (_10329_, _10328_, _10327_);
  nor (_10330_, _10329_, _10326_);
  and (_10331_, _10330_, _10267_);
  or (_10332_, _10331_, _10090_);
  nor (_10333_, _10332_, _09478_);
  nor (_10334_, _10332_, \oc8051_golden_model_1.B [7]);
  nor (_10335_, _10334_, _10045_);
  not (_10336_, _10335_);
  not (_10337_, \oc8051_golden_model_1.B [6]);
  and (_10338_, _10321_, _10277_);
  nor (_10339_, _10338_, _10322_);
  nor (_10340_, _10339_, _10330_);
  not (_10341_, _10330_);
  nor (_10342_, _10341_, _10273_);
  nor (_10343_, _10342_, _10340_);
  nor (_10344_, _10343_, _10337_);
  and (_10345_, _10343_, _10337_);
  nor (_10346_, _10286_, _10285_);
  nor (_10347_, _10346_, _10319_);
  and (_10348_, _10346_, _10319_);
  or (_10349_, _10348_, _10347_);
  nor (_10350_, _10349_, _10330_);
  nor (_10351_, _10341_, _10284_);
  nor (_10352_, _10351_, _10350_);
  nor (_10353_, _10352_, _10099_);
  and (_10354_, _10352_, _10099_);
  not (_10355_, _10354_);
  and (_10356_, _10317_, _10314_);
  nor (_10357_, _10356_, _10318_);
  nor (_10358_, _10357_, _10330_);
  nor (_10359_, _10341_, _10291_);
  nor (_10360_, _10359_, _10358_);
  nor (_10361_, _10360_, _10098_);
  and (_10362_, _10330_, _10299_);
  nor (_10363_, _10301_, _10300_);
  and (_10364_, _10363_, _10312_);
  nor (_10365_, _10363_, _10312_);
  nor (_10366_, _10365_, _10364_);
  nor (_10367_, _10366_, _10330_);
  or (_10368_, _10367_, _10362_);
  nor (_10369_, _10368_, _10097_);
  and (_10370_, _10368_, _10097_);
  nor (_10371_, _10370_, _10369_);
  nor (_10372_, _10310_, _10308_);
  or (_10373_, _10372_, _10311_);
  nor (_10374_, _10373_, _10330_);
  and (_10375_, _10330_, _10305_);
  nor (_10376_, _10375_, _10374_);
  and (_10377_, _10376_, \oc8051_golden_model_1.B [2]);
  nor (_10378_, _10376_, \oc8051_golden_model_1.B [2]);
  nor (_10379_, _10378_, _10377_);
  and (_10380_, _10379_, _10371_);
  and (_10381_, _10330_, _06044_);
  nor (_10382_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  nor (_10383_, _10382_, _10006_);
  nor (_10384_, _10330_, _10383_);
  nor (_10385_, _10384_, _10381_);
  and (_10386_, _10385_, _10081_);
  nor (_10387_, _10385_, _10081_);
  and (_10388_, _10086_, \oc8051_golden_model_1.ACC [0]);
  not (_10389_, _10388_);
  nor (_10390_, _10389_, _10387_);
  nor (_10391_, _10390_, _10386_);
  and (_10392_, _10391_, _10380_);
  not (_10393_, _10392_);
  and (_10394_, _10377_, _10371_);
  nor (_10395_, _10394_, _10369_);
  and (_10396_, _10395_, _10393_);
  and (_10397_, _10360_, _10098_);
  nor (_10398_, _10397_, _10396_);
  or (_10399_, _10398_, _10361_);
  and (_10400_, _10399_, _10355_);
  nor (_10401_, _10400_, _10353_);
  nor (_10402_, _10401_, _10345_);
  or (_10403_, _10402_, _10344_);
  and (_10404_, _10403_, _10336_);
  nor (_10405_, _10404_, _10333_);
  nor (_10406_, _10345_, _10344_);
  and (_10407_, _10406_, _10336_);
  nor (_10408_, _10397_, _10361_);
  nor (_10409_, _10354_, _10353_);
  and (_10410_, _10409_, _10408_);
  and (_10411_, _10410_, _10407_);
  and (_10412_, \oc8051_golden_model_1.B [0], _06018_);
  not (_10413_, _10412_);
  nor (_10414_, _10387_, _10386_);
  and (_10415_, _10414_, _10413_);
  and (_10416_, _10415_, _10389_);
  and (_10417_, _10416_, _10380_);
  and (_10418_, _10417_, _10411_);
  nor (_10419_, _10418_, _10405_);
  or (_10420_, _10419_, _10090_);
  and (_10421_, _10332_, _09480_);
  and (_10422_, _10421_, _10420_);
  or (_10423_, _10422_, _10080_);
  or (_10424_, _10423_, _10079_);
  and (_10425_, _09034_, _07933_);
  or (_10426_, _09482_, _09025_);
  or (_10427_, _10426_, _10425_);
  and (_10428_, _08806_, _07933_);
  or (_10429_, _10428_, _09482_);
  or (_10430_, _10429_, _06216_);
  and (_10431_, _10430_, _09030_);
  and (_10432_, _10431_, _10427_);
  and (_10433_, _10432_, _10424_);
  and (_10434_, _09042_, _07933_);
  or (_10435_, _10434_, _09482_);
  and (_10436_, _10435_, _06524_);
  or (_10437_, _10436_, _10433_);
  and (_10438_, _10437_, _07219_);
  or (_10439_, _09482_, _08026_);
  and (_10440_, _10429_, _06426_);
  and (_10441_, _10440_, _10439_);
  or (_10442_, _10441_, _10438_);
  and (_10443_, _10442_, _07217_);
  and (_10444_, _09499_, _06532_);
  and (_10445_, _10444_, _10439_);
  or (_10446_, _10445_, _06437_);
  or (_10447_, _10446_, _10443_);
  and (_10448_, _09033_, _07933_);
  or (_10449_, _09482_, _07229_);
  or (_10450_, _10449_, _10448_);
  and (_10451_, _10450_, _07231_);
  and (_10452_, _10451_, _10447_);
  not (_10453_, _07933_);
  nor (_10454_, _09041_, _10453_);
  or (_10455_, _10454_, _09482_);
  and (_10456_, _10455_, _06535_);
  or (_10457_, _10456_, _06559_);
  or (_10458_, _10457_, _10452_);
  or (_10459_, _09496_, _07240_);
  and (_10460_, _10459_, _05933_);
  and (_10461_, _10460_, _10458_);
  and (_10462_, _09493_, _05932_);
  or (_10463_, _10462_, _06566_);
  or (_10464_, _10463_, _10461_);
  and (_10465_, _08534_, _07933_);
  or (_10466_, _09482_, _06570_);
  or (_10467_, _10466_, _10465_);
  and (_10468_, _10467_, _01320_);
  and (_10469_, _10468_, _10464_);
  or (_10470_, _10469_, _09479_);
  and (_40311_, _10470_, _42355_);
  nor (_10471_, _01320_, _08737_);
  and (_10472_, _05993_, _06397_);
  nand (_10473_, _10472_, _10105_);
  and (_10474_, _06418_, _05993_);
  not (_10475_, _10474_);
  nor (_10476_, _07446_, _06904_);
  nor (_10477_, _07930_, _08737_);
  and (_10478_, _09033_, _07930_);
  or (_10479_, _10478_, _10477_);
  and (_10480_, _10479_, _06437_);
  and (_10481_, _06418_, _06000_);
  or (_10482_, _06181_, _05985_);
  and (_10483_, _08536_, _07930_);
  or (_10484_, _10483_, _10477_);
  or (_10485_, _10484_, _06260_);
  and (_10486_, _06418_, _05938_);
  not (_10487_, _10486_);
  and (_10488_, _08374_, \oc8051_golden_model_1.PSW [7]);
  and (_10489_, _10488_, _08325_);
  and (_10490_, _10489_, _08424_);
  and (_10491_, _10490_, _08280_);
  and (_10492_, _10491_, _08528_);
  and (_10493_, _10492_, _08231_);
  and (_10494_, _10493_, _08128_);
  nor (_10495_, _10494_, _08025_);
  and (_10496_, _10494_, _08025_);
  nor (_10497_, _10496_, _10495_);
  and (_10498_, _10497_, \oc8051_golden_model_1.ACC [7]);
  nor (_10499_, _10497_, \oc8051_golden_model_1.ACC [7]);
  nor (_10500_, _10499_, _10498_);
  not (_10501_, _10500_);
  nor (_10502_, _10493_, _08128_);
  nor (_10503_, _10502_, _10494_);
  nor (_10504_, _10503_, _10105_);
  nor (_10505_, _10492_, _08231_);
  nor (_10506_, _10505_, _10493_);
  and (_10507_, _10506_, _10152_);
  nor (_10508_, _10506_, _10152_);
  nor (_10509_, _10491_, _08528_);
  nor (_10510_, _10509_, _10492_);
  nor (_10511_, _10510_, _10123_);
  nor (_10512_, _10511_, _10508_);
  nor (_10513_, _10512_, _10507_);
  nor (_10514_, _10508_, _10507_);
  not (_10515_, _10514_);
  and (_10516_, _10510_, _10123_);
  or (_10517_, _10516_, _10511_);
  or (_10518_, _10517_, _10515_);
  nor (_10519_, _10490_, _08280_);
  nor (_10520_, _10519_, _10491_);
  nor (_10521_, _10520_, _10248_);
  and (_10522_, _10520_, _10248_);
  nor (_10523_, _10522_, _10521_);
  nor (_10524_, _10489_, _08424_);
  nor (_10525_, _10524_, _10490_);
  nor (_10526_, _10525_, _10198_);
  and (_10527_, _10525_, _10198_);
  nor (_10528_, _10527_, _10526_);
  and (_10529_, _10528_, _10523_);
  nor (_10530_, _10488_, _08325_);
  nor (_10531_, _10530_, _10489_);
  nor (_10532_, _10531_, _06044_);
  and (_10533_, _10531_, _06044_);
  nor (_10534_, _08374_, \oc8051_golden_model_1.PSW [7]);
  nor (_10535_, _10534_, _10488_);
  and (_10536_, _10535_, _06018_);
  nor (_10537_, _10536_, _10533_);
  or (_10538_, _10537_, _10532_);
  and (_10539_, _10538_, _10529_);
  and (_10540_, _10526_, _10523_);
  or (_10541_, _10540_, _10521_);
  nor (_10542_, _10541_, _10539_);
  nor (_10543_, _10542_, _10518_);
  nor (_10544_, _10543_, _10513_);
  and (_10545_, _10503_, _10105_);
  nor (_10546_, _10504_, _10545_);
  not (_10547_, _10546_);
  nor (_10548_, _10547_, _10544_);
  or (_10549_, _10548_, _10504_);
  and (_10550_, _10549_, _10501_);
  nor (_10551_, _10549_, _10501_);
  or (_10552_, _10551_, _10550_);
  and (_10553_, _10552_, _06380_);
  and (_10554_, _06256_, _05938_);
  nor (_10555_, _10554_, _06805_);
  and (_10556_, _09384_, \oc8051_golden_model_1.PSW [7]);
  and (_10557_, _10556_, _09339_);
  and (_10558_, _10557_, _09293_);
  and (_10559_, _10558_, _09247_);
  and (_10560_, _10559_, _09437_);
  and (_10561_, _10560_, _09436_);
  and (_10562_, _10561_, _09435_);
  nor (_10563_, _10562_, _09067_);
  and (_10564_, _10562_, _09067_);
  nor (_10565_, _10564_, _10563_);
  and (_10566_, _10565_, \oc8051_golden_model_1.ACC [7]);
  nor (_10567_, _10565_, \oc8051_golden_model_1.ACC [7]);
  nor (_10568_, _10567_, _10566_);
  not (_10569_, _10568_);
  nor (_10570_, _10561_, _09435_);
  nor (_10571_, _10570_, _10562_);
  nor (_10572_, _10571_, _10105_);
  nor (_10573_, _10560_, _09436_);
  nor (_10574_, _10573_, _10561_);
  and (_10575_, _10574_, _10152_);
  nor (_10576_, _10574_, _10152_);
  nor (_10577_, _10559_, _09437_);
  nor (_10578_, _10577_, _10560_);
  nor (_10579_, _10578_, _10123_);
  nor (_10580_, _10579_, _10576_);
  nor (_10581_, _10580_, _10575_);
  nor (_10582_, _10576_, _10575_);
  not (_10583_, _10582_);
  and (_10584_, _10578_, _10123_);
  or (_10585_, _10584_, _10579_);
  or (_10586_, _10585_, _10583_);
  nor (_10587_, _10558_, _09247_);
  nor (_10588_, _10587_, _10559_);
  nor (_10589_, _10588_, _10248_);
  and (_10590_, _10588_, _10248_);
  nor (_10591_, _10590_, _10589_);
  nor (_10592_, _10557_, _09293_);
  nor (_10593_, _10592_, _10558_);
  nor (_10594_, _10593_, _10198_);
  and (_10595_, _10593_, _10198_);
  nor (_10596_, _10595_, _10594_);
  and (_10597_, _10596_, _10591_);
  nor (_10598_, _10556_, _09339_);
  nor (_10599_, _10598_, _10557_);
  nor (_10600_, _10599_, _06044_);
  and (_10601_, _10599_, _06044_);
  nor (_10602_, _09384_, \oc8051_golden_model_1.PSW [7]);
  nor (_10603_, _10602_, _10556_);
  and (_10604_, _10603_, _06018_);
  nor (_10605_, _10604_, _10601_);
  or (_10606_, _10605_, _10600_);
  and (_10607_, _10606_, _10597_);
  and (_10608_, _10594_, _10591_);
  or (_10609_, _10608_, _10589_);
  nor (_10610_, _10609_, _10607_);
  nor (_10611_, _10610_, _10586_);
  nor (_10612_, _10611_, _10581_);
  and (_10613_, _10571_, _10105_);
  nor (_10614_, _10572_, _10613_);
  not (_10615_, _10614_);
  nor (_10616_, _10615_, _10612_);
  or (_10617_, _10616_, _10572_);
  and (_10618_, _10617_, _10569_);
  nor (_10619_, _10617_, _10569_);
  or (_10620_, _10619_, _10618_);
  or (_10621_, _10620_, _10555_);
  nor (_10622_, _05954_, _05880_);
  not (_10623_, _10622_);
  or (_10624_, _10623_, _08536_);
  nor (_10625_, _08596_, _08737_);
  and (_10626_, _08626_, _08596_);
  or (_10627_, _10626_, _10625_);
  or (_10628_, _10627_, _06282_);
  and (_10629_, _10628_, _07169_);
  and (_10630_, _08637_, _07930_);
  or (_10631_, _10630_, _10477_);
  and (_10632_, _10631_, _06285_);
  and (_10633_, _06418_, _06357_);
  not (_10634_, _10633_);
  or (_10635_, _10634_, _08731_);
  and (_10636_, _06286_, _05960_);
  and (_10637_, _06256_, _06357_);
  not (_10638_, _10637_);
  and (_10639_, _06253_, _06357_);
  nor (_10640_, _10639_, _06358_);
  and (_10641_, _10640_, _10638_);
  nor (_10642_, _07446_, _05959_);
  and (_10643_, _06414_, _06357_);
  nor (_10644_, _10643_, _10642_);
  nand (_10645_, _10644_, _10641_);
  and (_10646_, _10645_, _08536_);
  nor (_10647_, _06755_, _08737_);
  and (_10648_, _06755_, _08737_);
  nor (_10649_, _10648_, _10647_);
  nor (_10650_, _10649_, _10645_);
  or (_10651_, _10650_, _10633_);
  or (_10652_, _10651_, _10646_);
  and (_10653_, _10652_, _10636_);
  and (_10654_, _10653_, _10635_);
  or (_10655_, _10654_, _10632_);
  and (_10656_, _06418_, _06280_);
  not (_10657_, _10656_);
  and (_10658_, _10657_, _10655_);
  nor (_10659_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor (_10660_, _10659_, _10248_);
  and (_10661_, _10660_, \oc8051_golden_model_1.ACC [4]);
  and (_10662_, _10661_, \oc8051_golden_model_1.ACC [5]);
  and (_10663_, _10662_, \oc8051_golden_model_1.ACC [6]);
  and (_10664_, _10663_, \oc8051_golden_model_1.ACC [7]);
  nor (_10666_, _10663_, \oc8051_golden_model_1.ACC [7]);
  nor (_10667_, _10666_, _10664_);
  nor (_10668_, _10661_, \oc8051_golden_model_1.ACC [5]);
  nor (_10669_, _10668_, _10662_);
  nor (_10670_, _10662_, \oc8051_golden_model_1.ACC [6]);
  nor (_10671_, _10670_, _10663_);
  nor (_10672_, _10671_, _10669_);
  not (_10673_, _10672_);
  and (_10674_, _10673_, _10667_);
  not (_10675_, _10674_);
  nor (_10677_, _10664_, \oc8051_golden_model_1.PSW [7]);
  and (_10678_, _10677_, _10675_);
  nor (_10679_, _10678_, _10672_);
  or (_10680_, _10679_, _10667_);
  and (_10681_, _10675_, _10656_);
  and (_10682_, _10681_, _10680_);
  or (_10683_, _10682_, _06281_);
  or (_10684_, _10683_, _10658_);
  and (_10685_, _10684_, _10629_);
  and (_10686_, _10484_, _06354_);
  or (_10688_, _10686_, _10622_);
  or (_10689_, _10688_, _10685_);
  and (_10690_, _10689_, _10624_);
  or (_10691_, _10690_, _07174_);
  not (_10692_, _07174_);
  or (_10693_, _08731_, _10692_);
  and (_10694_, _10693_, _06346_);
  and (_10695_, _10694_, _10691_);
  and (_10696_, _06418_, _06275_);
  nor (_10697_, _08025_, _06346_);
  or (_10699_, _10697_, _10696_);
  or (_10700_, _10699_, _10695_);
  nand (_10701_, _10696_, _10248_);
  and (_10702_, _10701_, _10700_);
  or (_10703_, _10702_, _06277_);
  and (_10704_, _08622_, _08596_);
  or (_10705_, _10704_, _10625_);
  or (_10706_, _10705_, _06278_);
  and (_10707_, _10706_, _06271_);
  and (_10708_, _10707_, _10703_);
  or (_10710_, _10625_, _08768_);
  and (_10711_, _10710_, _06270_);
  and (_10712_, _10711_, _10627_);
  or (_10713_, _10712_, _09520_);
  or (_10714_, _10713_, _10708_);
  nor (_10715_, _10025_, _10023_);
  nor (_10716_, _10715_, _10026_);
  or (_10717_, _10716_, _10059_);
  and (_10718_, _07466_, _05938_);
  not (_10719_, _10718_);
  nand (_10721_, _06414_, _05938_);
  or (_10722_, _07446_, _05939_);
  and (_10723_, _10722_, _10721_);
  and (_10724_, _10723_, _10719_);
  and (_10725_, _10724_, _10717_);
  and (_10726_, _10725_, _10714_);
  not (_10727_, _10555_);
  and (_10728_, _09428_, \oc8051_golden_model_1.PSW [7]);
  and (_10729_, _10728_, _08536_);
  nor (_10730_, _10728_, _08536_);
  or (_10732_, _10730_, _10729_);
  and (_10733_, _10732_, \oc8051_golden_model_1.ACC [7]);
  nor (_10734_, _10732_, \oc8051_golden_model_1.ACC [7]);
  nor (_10735_, _10734_, _10733_);
  and (_10736_, _09427_, \oc8051_golden_model_1.PSW [7]);
  nor (_10737_, _10736_, _09418_);
  nor (_10738_, _10737_, _10728_);
  nor (_10739_, _10738_, _10105_);
  and (_10740_, _09426_, \oc8051_golden_model_1.PSW [7]);
  nor (_10741_, _10740_, _09419_);
  nor (_10742_, _10741_, _10736_);
  and (_10743_, _10742_, _10152_);
  nor (_10744_, _10742_, _10152_);
  and (_10745_, _09425_, \oc8051_golden_model_1.PSW [7]);
  nor (_10746_, _10745_, _09420_);
  nor (_10747_, _10746_, _10740_);
  nor (_10748_, _10747_, _10123_);
  nor (_10749_, _10748_, _10744_);
  nor (_10750_, _10749_, _10743_);
  nor (_10751_, _10744_, _10743_);
  not (_10752_, _10751_);
  and (_10753_, _10747_, _10123_);
  or (_10754_, _10753_, _10748_);
  or (_10755_, _10754_, _10752_);
  and (_10756_, _09424_, \oc8051_golden_model_1.PSW [7]);
  nor (_10757_, _10756_, _09421_);
  nor (_10758_, _10757_, _10745_);
  nor (_10759_, _10758_, _10248_);
  and (_10760_, _10758_, _10248_);
  nor (_10761_, _10760_, _10759_);
  and (_10762_, _09423_, \oc8051_golden_model_1.PSW [7]);
  nor (_10763_, _10762_, _08662_);
  nor (_10764_, _10763_, _10756_);
  nor (_10765_, _10764_, _10198_);
  and (_10766_, _10764_, _10198_);
  nor (_10767_, _10766_, _10765_);
  and (_10768_, _10767_, _10761_);
  and (_10769_, _07135_, \oc8051_golden_model_1.PSW [7]);
  nor (_10770_, _10769_, _09422_);
  nor (_10771_, _10770_, _10762_);
  nor (_10772_, _10771_, _06044_);
  and (_10773_, _10771_, _06044_);
  not (_10774_, \oc8051_golden_model_1.PSW [7]);
  and (_10775_, _07157_, _10774_);
  nor (_10776_, _10775_, _10769_);
  and (_10777_, _10776_, _06018_);
  nor (_10778_, _10777_, _10773_);
  or (_10779_, _10778_, _10772_);
  nand (_10780_, _10779_, _10768_);
  and (_10781_, _10765_, _10761_);
  nor (_10782_, _10781_, _10759_);
  and (_10783_, _10782_, _10780_);
  nor (_10784_, _10783_, _10755_);
  nor (_10785_, _10784_, _10750_);
  and (_10786_, _10738_, _10105_);
  nor (_10787_, _10739_, _10786_);
  not (_10788_, _10787_);
  nor (_10789_, _10788_, _10785_);
  or (_10790_, _10789_, _10739_);
  nor (_10791_, _10790_, _10735_);
  and (_10792_, _10790_, _10735_);
  or (_10793_, _10792_, _10791_);
  nor (_10794_, _10793_, _10724_);
  or (_10795_, _10794_, _10727_);
  or (_10796_, _10795_, _10726_);
  and (_10797_, _10796_, _06386_);
  and (_10798_, _10797_, _10621_);
  or (_10799_, _10798_, _10553_);
  and (_10800_, _10799_, _10487_);
  and (_10801_, _08787_, _07898_);
  and (_10802_, _10801_, _07932_);
  and (_10803_, _10801_, _07883_);
  and (_10804_, _10803_, _07589_);
  nor (_10805_, _10804_, _06181_);
  nor (_10806_, _10805_, _10802_);
  nor (_10807_, _10806_, _08737_);
  and (_10808_, _10806_, _08737_);
  nor (_10809_, _10808_, _10807_);
  nor (_10810_, _10803_, _07589_);
  nor (_10811_, _10810_, _10804_);
  nor (_10812_, _10811_, _10105_);
  and (_10813_, _10801_, _07889_);
  nor (_10814_, _10813_, _07873_);
  nor (_10815_, _10814_, _10803_);
  and (_10816_, _10815_, _10152_);
  nor (_10817_, _10815_, _10152_);
  nor (_10818_, _10817_, _10816_);
  not (_10819_, _10818_);
  nor (_10820_, _10801_, _07889_);
  nor (_10821_, _10820_, _10813_);
  nor (_10822_, _10821_, _10123_);
  and (_10823_, _10821_, _10123_);
  or (_10824_, _10823_, _10822_);
  or (_10825_, _10824_, _10819_);
  nor (_10826_, _08788_, _06356_);
  nor (_10827_, _10826_, _10801_);
  nor (_10828_, _10827_, _10248_);
  and (_10829_, _10827_, _10248_);
  nor (_10830_, _10829_, _10828_);
  nor (_10831_, _08787_, _06647_);
  or (_10832_, _10831_, _08788_);
  and (_10833_, _10832_, \oc8051_golden_model_1.ACC [2]);
  nor (_10834_, _10832_, \oc8051_golden_model_1.ACC [2]);
  nor (_10835_, _10834_, _10833_);
  and (_10836_, _10835_, _10830_);
  nor (_10837_, _08786_, _06996_);
  nor (_10838_, _10837_, _08787_);
  nor (_10839_, _10838_, _06044_);
  and (_10840_, _10838_, _06044_);
  nor (_10841_, _06248_, \oc8051_golden_model_1.PSW [7]);
  nor (_10842_, _10841_, _08786_);
  and (_10843_, _10842_, _06018_);
  nor (_10844_, _10843_, _10840_);
  or (_10845_, _10844_, _10839_);
  nand (_10846_, _10845_, _10836_);
  and (_10847_, _10833_, _10830_);
  nor (_10848_, _10847_, _10828_);
  and (_10849_, _10848_, _10846_);
  nor (_10850_, _10849_, _10825_);
  and (_10851_, _10822_, _10818_);
  nor (_10852_, _10851_, _10817_);
  not (_10853_, _10852_);
  nor (_10854_, _10853_, _10850_);
  and (_10855_, _10811_, _10105_);
  nor (_10856_, _10812_, _10855_);
  not (_10857_, _10856_);
  nor (_10858_, _10857_, _10854_);
  or (_10859_, _10858_, _10812_);
  nor (_10860_, _10859_, _10809_);
  and (_10861_, _10859_, _10809_);
  or (_10862_, _10861_, _10860_);
  nor (_10863_, _10862_, _10487_);
  or (_10864_, _10863_, _10800_);
  and (_10865_, _10864_, _05940_);
  and (_10866_, _06181_, _05976_);
  or (_10867_, _10866_, _10865_);
  and (_10868_, _10867_, _06267_);
  and (_10869_, _08789_, _08596_);
  or (_10870_, _10869_, _10625_);
  and (_10871_, _10870_, _06266_);
  or (_10872_, _10871_, _06259_);
  or (_10873_, _10872_, _10868_);
  and (_10874_, _10873_, _10485_);
  or (_10875_, _10874_, _09486_);
  and (_10876_, _08731_, _07930_);
  or (_10877_, _10477_, _06258_);
  or (_10878_, _10877_, _10876_);
  and (_10879_, _10878_, _06251_);
  and (_10880_, _10879_, _10875_);
  and (_10881_, _09004_, _07930_);
  or (_10882_, _10881_, _10477_);
  and (_10883_, _10882_, _05972_);
  or (_10884_, _10883_, _09480_);
  or (_10885_, _10884_, _10880_);
  or (_10886_, _10094_, _09481_);
  and (_10887_, _10886_, _10885_);
  or (_10888_, _10887_, _05984_);
  and (_10889_, _10888_, _10482_);
  or (_10890_, _10889_, _06215_);
  and (_10891_, _06418_, _06003_);
  not (_10892_, _10891_);
  and (_10893_, _08806_, _07930_);
  or (_10894_, _10893_, _10477_);
  or (_10895_, _10894_, _06216_);
  and (_10896_, _10895_, _10892_);
  and (_10897_, _10896_, _10890_);
  and (_10898_, _10891_, _06181_);
  and (_10899_, _07466_, _06000_);
  or (_10900_, _10899_, _10898_);
  or (_10901_, _10900_, _10897_);
  and (_10902_, _08023_, _08737_);
  and (_10903_, _08536_, \oc8051_golden_model_1.ACC [7]);
  nor (_10904_, _10903_, _10902_);
  not (_10905_, _10899_);
  or (_10906_, _10905_, _10904_);
  not (_10907_, _06000_);
  nor (_10908_, _07446_, _10907_);
  not (_10909_, _10908_);
  and (_10910_, _10909_, _10906_);
  and (_10911_, _10910_, _10901_);
  and (_10912_, _10908_, _10904_);
  and (_10913_, _06414_, _06000_);
  or (_10914_, _10913_, _10912_);
  or (_10915_, _10914_, _10911_);
  and (_10916_, _06256_, _06000_);
  or (_10917_, _10916_, _06868_);
  not (_10918_, _10917_);
  not (_10919_, _10913_);
  or (_10920_, _10919_, _10904_);
  and (_10921_, _10920_, _10918_);
  and (_10922_, _10921_, _10915_);
  and (_10923_, _09067_, _08737_);
  and (_10924_, _08731_, \oc8051_golden_model_1.ACC [7]);
  nor (_10925_, _10924_, _10923_);
  and (_10926_, _10917_, _10925_);
  or (_10927_, _10926_, _06526_);
  or (_10928_, _10927_, _10922_);
  or (_10929_, _09042_, _06527_);
  and (_10930_, _10929_, _10928_);
  or (_10931_, _10930_, _10481_);
  nor (_10932_, _06181_, \oc8051_golden_model_1.ACC [7]);
  and (_10933_, _06181_, \oc8051_golden_model_1.ACC [7]);
  nor (_10934_, _10933_, _10932_);
  not (_10935_, _10481_);
  or (_10936_, _10935_, _10934_);
  and (_10937_, _10936_, _10931_);
  or (_10938_, _10937_, _06398_);
  and (_10939_, _09034_, _07930_);
  or (_10940_, _10939_, _10477_);
  or (_10941_, _10940_, _09025_);
  and (_10942_, _10941_, _09030_);
  and (_10943_, _10942_, _10938_);
  and (_10944_, _06702_, _06012_);
  and (_10945_, _10477_, _06524_);
  or (_10946_, _10945_, _10944_);
  or (_10947_, _10946_, _10943_);
  not (_10948_, _10944_);
  or (_10949_, _10903_, _10948_);
  and (_10950_, _06801_, _06012_);
  not (_10951_, _10950_);
  not (_10952_, _05928_);
  and (_10953_, _05882_, _10952_);
  nor (_10954_, _10953_, _06714_);
  or (_10955_, _10954_, _06875_);
  and (_10956_, _10955_, _10951_);
  and (_10957_, _10956_, _10949_);
  and (_10958_, _10957_, _10947_);
  nor (_10959_, _07158_, _06875_);
  not (_10960_, _10956_);
  and (_10961_, _10960_, _10903_);
  or (_10962_, _10961_, _10959_);
  or (_10963_, _10962_, _10958_);
  not (_10964_, _10959_);
  or (_10965_, _10964_, _10924_);
  and (_10966_, _10965_, _06531_);
  and (_10967_, _10966_, _10963_);
  and (_10968_, _06418_, _06012_);
  nor (_10969_, _10968_, _06530_);
  not (_10970_, _10969_);
  or (_10971_, _10968_, _09040_);
  and (_10972_, _10971_, _10970_);
  or (_10973_, _10972_, _10967_);
  not (_10974_, _10968_);
  or (_10975_, _10974_, _10933_);
  and (_10976_, _10975_, _07219_);
  and (_10977_, _10976_, _10973_);
  nand (_10978_, _10894_, _06426_);
  nor (_10979_, _10978_, _09041_);
  or (_10980_, _10979_, _10977_);
  and (_10981_, _06702_, _06007_);
  not (_10982_, _10981_);
  and (_10983_, _06339_, _06007_);
  nor (_10984_, _07472_, _07059_);
  nor (_10985_, _10984_, _10983_);
  nand (_10986_, _10985_, _10982_);
  not (_10987_, _10986_);
  and (_10988_, _10987_, _10980_);
  and (_10989_, _09006_, _06007_);
  nor (_10990_, _10989_, _06882_);
  not (_10991_, _10990_);
  nor (_10992_, _10987_, _10902_);
  or (_10993_, _10992_, _10991_);
  or (_10994_, _10993_, _10988_);
  not (_10995_, _06881_);
  nand (_10996_, _10991_, _10902_);
  and (_10997_, _10996_, _10995_);
  and (_10998_, _10997_, _10994_);
  nor (_10999_, _10902_, _10995_);
  nor (_11000_, _07158_, _07059_);
  or (_11001_, _11000_, _10999_);
  or (_11002_, _11001_, _10998_);
  nand (_11003_, _11000_, _10923_);
  and (_11004_, _11003_, _06538_);
  and (_11005_, _11004_, _11002_);
  and (_11006_, _06418_, _06007_);
  nor (_11007_, _11006_, _06537_);
  not (_11008_, _11007_);
  not (_11009_, _11006_);
  nand (_11010_, _11009_, _09041_);
  and (_11011_, _11010_, _11008_);
  or (_11012_, _11011_, _11005_);
  nand (_11013_, _11006_, _10932_);
  and (_11014_, _11013_, _07229_);
  and (_11015_, _11014_, _11012_);
  nor (_11016_, _11015_, _10480_);
  and (_11017_, _07466_, _06010_);
  not (_11018_, _11017_);
  and (_11019_, _06414_, _06010_);
  not (_11020_, _11019_);
  or (_11021_, _07446_, _06889_);
  and (_11022_, _11021_, _11020_);
  and (_11023_, _11022_, _11018_);
  not (_11024_, _11023_);
  or (_11025_, _11024_, _11016_);
  and (_11026_, _06256_, _06010_);
  nor (_11027_, _11026_, _06892_);
  and (_11028_, _10738_, \oc8051_golden_model_1.ACC [6]);
  and (_11029_, _10742_, \oc8051_golden_model_1.ACC [5]);
  nand (_11030_, _10747_, \oc8051_golden_model_1.ACC [4]);
  and (_11031_, _10758_, \oc8051_golden_model_1.ACC [3]);
  and (_11032_, _10764_, \oc8051_golden_model_1.ACC [2]);
  and (_11033_, _10771_, \oc8051_golden_model_1.ACC [1]);
  nor (_11034_, _10773_, _10772_);
  not (_11035_, _11034_);
  and (_11036_, _10776_, \oc8051_golden_model_1.ACC [0]);
  and (_11037_, _11036_, _11035_);
  nor (_11038_, _11037_, _11033_);
  nor (_11039_, _11038_, _10767_);
  nor (_11040_, _11039_, _11032_);
  nor (_11041_, _11040_, _10761_);
  or (_11042_, _11041_, _11031_);
  nand (_11043_, _11042_, _10754_);
  and (_11044_, _11043_, _11030_);
  nor (_11045_, _11044_, _10751_);
  or (_11046_, _11045_, _11029_);
  and (_11047_, _11046_, _10788_);
  nor (_11048_, _11047_, _11028_);
  nor (_11049_, _11048_, _10735_);
  and (_11050_, _11048_, _10735_);
  nor (_11051_, _11050_, _11049_);
  nand (_11052_, _11051_, _11024_);
  and (_11053_, _11052_, _11027_);
  and (_11054_, _11053_, _11025_);
  nand (_11055_, _10571_, \oc8051_golden_model_1.ACC [6]);
  and (_11056_, _10574_, \oc8051_golden_model_1.ACC [5]);
  nand (_11057_, _10578_, \oc8051_golden_model_1.ACC [4]);
  and (_11058_, _10588_, \oc8051_golden_model_1.ACC [3]);
  and (_11059_, _10593_, \oc8051_golden_model_1.ACC [2]);
  and (_11060_, _10599_, \oc8051_golden_model_1.ACC [1]);
  nor (_11061_, _10601_, _10600_);
  not (_11062_, _11061_);
  and (_11063_, _10603_, \oc8051_golden_model_1.ACC [0]);
  and (_11064_, _11063_, _11062_);
  nor (_11065_, _11064_, _11060_);
  nor (_11066_, _11065_, _10596_);
  nor (_11067_, _11066_, _11059_);
  nor (_11068_, _11067_, _10591_);
  or (_11069_, _11068_, _11058_);
  nand (_11070_, _11069_, _10585_);
  and (_11071_, _11070_, _11057_);
  nor (_11072_, _11071_, _10582_);
  or (_11073_, _11072_, _11056_);
  nand (_11074_, _11073_, _10615_);
  and (_11075_, _11074_, _11055_);
  nor (_11076_, _11075_, _10568_);
  and (_11077_, _11075_, _10568_);
  nor (_11078_, _11077_, _11076_);
  nor (_11079_, _11078_, _11027_);
  or (_11080_, _11079_, _06522_);
  or (_11081_, _11080_, _11054_);
  and (_11082_, _06418_, _06010_);
  not (_11083_, _11082_);
  nand (_11084_, _10503_, \oc8051_golden_model_1.ACC [6]);
  and (_11085_, _10506_, \oc8051_golden_model_1.ACC [5]);
  nand (_11086_, _10510_, \oc8051_golden_model_1.ACC [4]);
  and (_11087_, _10520_, \oc8051_golden_model_1.ACC [3]);
  and (_11088_, _10525_, \oc8051_golden_model_1.ACC [2]);
  and (_11089_, _10531_, \oc8051_golden_model_1.ACC [1]);
  nor (_11090_, _10533_, _10532_);
  not (_11091_, _11090_);
  and (_11092_, _10535_, \oc8051_golden_model_1.ACC [0]);
  and (_11093_, _11092_, _11091_);
  nor (_11094_, _11093_, _11089_);
  nor (_11095_, _11094_, _10528_);
  nor (_11096_, _11095_, _11088_);
  nor (_11097_, _11096_, _10523_);
  or (_11098_, _11097_, _11087_);
  nand (_11099_, _11098_, _10517_);
  and (_11100_, _11099_, _11086_);
  nor (_11101_, _11100_, _10514_);
  or (_11102_, _11101_, _11085_);
  nand (_11103_, _11102_, _10547_);
  and (_11104_, _11103_, _11084_);
  nor (_11105_, _11104_, _10500_);
  and (_11106_, _11104_, _10500_);
  nor (_11107_, _11106_, _11105_);
  nand (_11108_, _11107_, _06522_);
  and (_11109_, _11108_, _11083_);
  and (_11110_, _11109_, _11081_);
  and (_11111_, _06010_, _06397_);
  nand (_11112_, _10811_, \oc8051_golden_model_1.ACC [6]);
  and (_11113_, _10815_, \oc8051_golden_model_1.ACC [5]);
  nand (_11114_, _10821_, \oc8051_golden_model_1.ACC [4]);
  and (_11115_, _10827_, \oc8051_golden_model_1.ACC [3]);
  nor (_11116_, _10832_, _10198_);
  and (_11117_, _10838_, \oc8051_golden_model_1.ACC [1]);
  nor (_11118_, _10840_, _10839_);
  not (_11119_, _11118_);
  and (_11120_, _10842_, \oc8051_golden_model_1.ACC [0]);
  and (_11121_, _11120_, _11119_);
  nor (_11122_, _11121_, _11117_);
  nor (_11123_, _11122_, _10835_);
  nor (_11124_, _11123_, _11116_);
  nor (_11125_, _11124_, _10830_);
  or (_11126_, _11125_, _11115_);
  nand (_11127_, _11126_, _10824_);
  and (_11128_, _11127_, _11114_);
  nor (_11129_, _11128_, _10818_);
  or (_11130_, _11129_, _11113_);
  nand (_11131_, _11130_, _10857_);
  and (_11132_, _11131_, _11112_);
  nor (_11133_, _11132_, _10809_);
  and (_11134_, _11132_, _10809_);
  nor (_11135_, _11134_, _11133_);
  nor (_11136_, _11135_, _11083_);
  or (_11137_, _11136_, _11111_);
  or (_11138_, _11137_, _11110_);
  and (_11139_, _11111_, \oc8051_golden_model_1.ACC [6]);
  and (_11140_, _07466_, _05993_);
  nor (_11141_, _11140_, _11139_);
  nand (_11142_, _11141_, _11138_);
  or (_11143_, _11142_, _10476_);
  and (_11144_, _06414_, _05993_);
  and (_11145_, _09418_, \oc8051_golden_model_1.ACC [6]);
  not (_11146_, _11145_);
  or (_11147_, _09418_, \oc8051_golden_model_1.ACC [6]);
  and (_11148_, _11147_, _11146_);
  and (_11149_, _09419_, \oc8051_golden_model_1.ACC [5]);
  and (_11150_, _08228_, _10152_);
  nor (_11151_, _11150_, _11149_);
  and (_11152_, _09420_, \oc8051_golden_model_1.ACC [4]);
  not (_11153_, _11152_);
  or (_11154_, _09420_, \oc8051_golden_model_1.ACC [4]);
  and (_11155_, _11154_, _11153_);
  and (_11156_, _09421_, \oc8051_golden_model_1.ACC [3]);
  and (_11157_, _07578_, _10248_);
  and (_11158_, _08662_, \oc8051_golden_model_1.ACC [2]);
  and (_11159_, _07760_, _10198_);
  nor (_11160_, _11159_, _11158_);
  and (_11161_, _09422_, \oc8051_golden_model_1.ACC [1]);
  and (_11162_, _07334_, _06044_);
  nor (_11163_, _11162_, _11161_);
  and (_11164_, _07135_, \oc8051_golden_model_1.ACC [0]);
  and (_11165_, _11164_, _11163_);
  nor (_11166_, _11165_, _11161_);
  not (_11167_, _11166_);
  and (_11168_, _11167_, _11160_);
  nor (_11169_, _11168_, _11158_);
  nor (_11170_, _11169_, _11157_);
  or (_11171_, _11170_, _11156_);
  and (_11172_, _11171_, _11155_);
  nor (_11173_, _11172_, _11152_);
  not (_11174_, _11173_);
  and (_11175_, _11174_, _11151_);
  or (_11176_, _11175_, _11149_);
  and (_11177_, _11176_, _11148_);
  nor (_11178_, _11177_, _11145_);
  nor (_11179_, _11178_, _10904_);
  and (_11180_, _11178_, _10904_);
  or (_11181_, _11180_, _11179_);
  not (_11182_, _11181_);
  nor (_11183_, _11182_, _11144_);
  and (_11184_, _05993_, _05879_);
  not (_11185_, _11184_);
  or (_11186_, _11185_, _11183_);
  and (_11187_, _11186_, _11143_);
  and (_11188_, _06253_, _05993_);
  and (_11189_, _06256_, _05993_);
  nor (_11190_, _11189_, _11188_);
  not (_11191_, _11190_);
  and (_11192_, _11181_, _11144_);
  or (_11193_, _11192_, _11191_);
  or (_11194_, _11193_, _11187_);
  and (_11195_, _09435_, \oc8051_golden_model_1.ACC [6]);
  not (_11196_, _11195_);
  or (_11197_, _09435_, \oc8051_golden_model_1.ACC [6]);
  and (_11198_, _11197_, _11196_);
  and (_11199_, _09436_, \oc8051_golden_model_1.ACC [5]);
  and (_11200_, _09157_, _10152_);
  or (_11201_, _11200_, _11199_);
  and (_11202_, _09437_, \oc8051_golden_model_1.ACC [4]);
  not (_11203_, _11202_);
  or (_11204_, _09437_, \oc8051_golden_model_1.ACC [4]);
  and (_11205_, _11204_, _11203_);
  and (_11206_, _09247_, \oc8051_golden_model_1.ACC [3]);
  nor (_11207_, _09247_, \oc8051_golden_model_1.ACC [3]);
  and (_11208_, _09293_, \oc8051_golden_model_1.ACC [2]);
  not (_11209_, _11208_);
  or (_11210_, _09293_, \oc8051_golden_model_1.ACC [2]);
  and (_11211_, _11210_, _11209_);
  not (_11212_, _11211_);
  and (_11213_, _09339_, \oc8051_golden_model_1.ACC [1]);
  not (_11214_, _11213_);
  or (_11215_, _09339_, \oc8051_golden_model_1.ACC [1]);
  and (_11216_, _11215_, _11214_);
  and (_11217_, _09384_, \oc8051_golden_model_1.ACC [0]);
  and (_11218_, _11217_, _11216_);
  nor (_11219_, _11218_, _11213_);
  nor (_11220_, _11219_, _11212_);
  nor (_11221_, _11220_, _11208_);
  nor (_11222_, _11221_, _11207_);
  or (_11223_, _11222_, _11206_);
  nand (_11224_, _11223_, _11205_);
  and (_11225_, _11224_, _11203_);
  nor (_11226_, _11225_, _11201_);
  or (_11227_, _11226_, _11199_);
  and (_11228_, _11227_, _11198_);
  nor (_11229_, _11228_, _11195_);
  and (_11230_, _11229_, _10925_);
  nor (_11231_, _11229_, _10925_);
  or (_11232_, _11231_, _11230_);
  or (_11233_, _11232_, _11190_);
  and (_11234_, _11233_, _06293_);
  and (_11235_, _11234_, _11194_);
  nor (_11236_, _08127_, _10105_);
  not (_11237_, _11236_);
  and (_11238_, _08127_, _10105_);
  nor (_11239_, _11238_, _11236_);
  nor (_11240_, _08230_, _10152_);
  and (_11241_, _08230_, _10152_);
  nor (_11242_, _08527_, _10123_);
  not (_11243_, _11242_);
  and (_11244_, _08527_, _10123_);
  nor (_11245_, _11244_, _11242_);
  nor (_11246_, _08279_, _10248_);
  and (_11247_, _08279_, _10248_);
  nor (_11248_, _08423_, _10198_);
  and (_11249_, _08423_, _10198_);
  nor (_11250_, _11249_, _11248_);
  nor (_11251_, _08324_, _06044_);
  and (_11252_, _08324_, _06044_);
  nor (_11253_, _11252_, _11251_);
  and (_11254_, _08374_, \oc8051_golden_model_1.ACC [0]);
  and (_11255_, _11254_, _11253_);
  nor (_11256_, _11255_, _11251_);
  not (_11257_, _11256_);
  and (_11258_, _11257_, _11250_);
  nor (_11259_, _11258_, _11248_);
  nor (_11260_, _11259_, _11247_);
  or (_11261_, _11260_, _11246_);
  nand (_11262_, _11261_, _11245_);
  and (_11263_, _11262_, _11243_);
  nor (_11264_, _11263_, _11241_);
  or (_11265_, _11264_, _11240_);
  nand (_11266_, _11265_, _11239_);
  and (_11267_, _11266_, _11237_);
  nor (_11268_, _11267_, _09042_);
  and (_11269_, _11267_, _09042_);
  or (_11270_, _11269_, _11268_);
  and (_11271_, _11270_, _06292_);
  or (_11272_, _11271_, _11235_);
  and (_11273_, _11272_, _10475_);
  nor (_11274_, _06325_, _10105_);
  and (_11275_, _06325_, _10105_);
  nor (_11276_, _11274_, _11275_);
  nor (_11277_, _06604_, _10152_);
  and (_11278_, _06604_, _10152_);
  nor (_11279_, _06961_, _10123_);
  not (_11280_, _11279_);
  and (_11281_, _06961_, _10123_);
  or (_11282_, _11281_, _11279_);
  not (_11283_, _11282_);
  nor (_11284_, _06212_, _10248_);
  nand (_11285_, _06212_, _10248_);
  nor (_11286_, _06646_, _10198_);
  and (_11287_, _06646_, \oc8051_golden_model_1.ACC [2]);
  nor (_11288_, _06646_, \oc8051_golden_model_1.ACC [2]);
  nor (_11289_, _11288_, _11287_);
  nor (_11290_, _06995_, _06044_);
  and (_11291_, _06995_, _06044_);
  nor (_11292_, _11290_, _11291_);
  and (_11293_, _06248_, \oc8051_golden_model_1.ACC [0]);
  and (_11294_, _11293_, _11292_);
  nor (_11295_, _11294_, _11290_);
  nor (_11296_, _11295_, _11289_);
  nor (_11297_, _11296_, _11286_);
  not (_11298_, _11297_);
  and (_11299_, _11298_, _11285_);
  or (_11300_, _11299_, _11284_);
  nand (_11301_, _11300_, _11283_);
  and (_11302_, _11301_, _11280_);
  nor (_11303_, _11302_, _11278_);
  or (_11304_, _11303_, _11277_);
  and (_11305_, _11304_, _11276_);
  nor (_11306_, _11305_, _11274_);
  nor (_11307_, _11306_, _10934_);
  and (_11308_, _11306_, _10934_);
  or (_11309_, _11308_, _11307_);
  and (_11310_, _11309_, _10474_);
  or (_11311_, _11310_, _10472_);
  or (_11312_, _11311_, _11273_);
  and (_11313_, _11312_, _10473_);
  or (_11314_, _11313_, _06559_);
  and (_11315_, _06418_, _05895_);
  not (_11316_, _11315_);
  or (_11317_, _10631_, _07240_);
  and (_11318_, _11317_, _11316_);
  and (_11319_, _11318_, _11314_);
  and (_11320_, _06397_, _05895_);
  and (_11321_, _10659_, _06018_);
  and (_11322_, _11321_, _10248_);
  and (_11323_, _11322_, _10123_);
  and (_11324_, _11323_, _10152_);
  and (_11325_, _11324_, _10105_);
  nor (_11326_, _11325_, _08737_);
  and (_11327_, _11325_, _08737_);
  or (_11328_, _11327_, _11326_);
  and (_11329_, _11328_, _11315_);
  or (_11330_, _11329_, _11320_);
  or (_11331_, _11330_, _11319_);
  nand (_11332_, _11320_, _10774_);
  and (_11333_, _11332_, _05933_);
  and (_11334_, _11333_, _11331_);
  and (_11335_, _10705_, _05932_);
  or (_11336_, _11335_, _06566_);
  or (_11337_, _11336_, _11334_);
  and (_11338_, _06418_, _05766_);
  not (_11339_, _11338_);
  and (_11340_, _08534_, _07930_);
  or (_11341_, _11340_, _10477_);
  or (_11342_, _11341_, _06570_);
  and (_11343_, _11342_, _11339_);
  and (_11344_, _11343_, _11337_);
  and (_11345_, _05766_, _06397_);
  and (_11346_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and (_11347_, _11346_, \oc8051_golden_model_1.ACC [2]);
  and (_11348_, _11347_, \oc8051_golden_model_1.ACC [3]);
  and (_11349_, _11348_, \oc8051_golden_model_1.ACC [4]);
  and (_11350_, _11349_, \oc8051_golden_model_1.ACC [5]);
  and (_11351_, _11350_, \oc8051_golden_model_1.ACC [6]);
  or (_11352_, _11351_, \oc8051_golden_model_1.ACC [7]);
  nand (_11353_, _11351_, \oc8051_golden_model_1.ACC [7]);
  and (_11354_, _11353_, _11352_);
  and (_11355_, _11354_, _11338_);
  or (_11356_, _11355_, _11345_);
  or (_11357_, _11356_, _11344_);
  nand (_11358_, _11345_, _06018_);
  and (_11359_, _11358_, _01320_);
  and (_11360_, _11359_, _11357_);
  or (_11361_, _11360_, _10471_);
  and (_40312_, _11361_, _42355_);
  not (_11362_, _07942_);
  and (_11363_, _11362_, \oc8051_golden_model_1.PCON [7]);
  and (_11364_, _08536_, _07942_);
  or (_11365_, _11364_, _11363_);
  or (_11366_, _11365_, _06260_);
  and (_11367_, _08637_, _07942_);
  or (_11368_, _11367_, _11363_);
  or (_11369_, _11368_, _06286_);
  and (_11370_, _07942_, \oc8051_golden_model_1.ACC [7]);
  or (_11371_, _11370_, _11363_);
  and (_11372_, _11371_, _07143_);
  and (_11373_, _07144_, \oc8051_golden_model_1.PCON [7]);
  or (_11374_, _11373_, _06285_);
  or (_11375_, _11374_, _11372_);
  and (_11376_, _11375_, _07169_);
  and (_11377_, _11376_, _11369_);
  and (_11378_, _11365_, _06354_);
  or (_11379_, _11378_, _11377_);
  and (_11380_, _11379_, _06346_);
  and (_11381_, _11371_, _06345_);
  or (_11382_, _11381_, _06259_);
  or (_11383_, _11382_, _11380_);
  and (_11384_, _11383_, _11366_);
  or (_11385_, _11384_, _09486_);
  and (_11386_, _08731_, _07942_);
  or (_11387_, _11363_, _06258_);
  or (_11388_, _11387_, _11386_);
  and (_11389_, _11388_, _06251_);
  and (_11390_, _11389_, _11385_);
  and (_11391_, _09004_, _07942_);
  or (_11392_, _11391_, _11363_);
  and (_11393_, _11392_, _05972_);
  or (_11394_, _11393_, _11390_);
  or (_11395_, _11394_, _10080_);
  and (_11396_, _09034_, _07942_);
  or (_11397_, _11363_, _09025_);
  or (_11398_, _11397_, _11396_);
  and (_11399_, _08806_, _07942_);
  or (_11400_, _11399_, _11363_);
  or (_11401_, _11400_, _06216_);
  and (_11402_, _11401_, _09030_);
  and (_11403_, _11402_, _11398_);
  and (_11404_, _11403_, _11395_);
  and (_11405_, _09042_, _07942_);
  or (_11406_, _11405_, _11363_);
  and (_11407_, _11406_, _06524_);
  or (_11408_, _11407_, _11404_);
  and (_11409_, _11408_, _07219_);
  or (_11410_, _11363_, _08026_);
  and (_11411_, _11400_, _06426_);
  and (_11412_, _11411_, _11410_);
  or (_11413_, _11412_, _11409_);
  and (_11414_, _11413_, _07217_);
  and (_11415_, _11371_, _06532_);
  and (_11416_, _11415_, _11410_);
  or (_11417_, _11416_, _06437_);
  or (_11418_, _11417_, _11414_);
  and (_11419_, _09033_, _07942_);
  or (_11420_, _11363_, _07229_);
  or (_11421_, _11420_, _11419_);
  and (_11422_, _11421_, _07231_);
  and (_11423_, _11422_, _11418_);
  nor (_11424_, _09041_, _11362_);
  or (_11425_, _11424_, _11363_);
  and (_11426_, _11425_, _06535_);
  or (_11427_, _11426_, _06559_);
  or (_11428_, _11427_, _11423_);
  or (_11429_, _11368_, _07240_);
  and (_11430_, _11429_, _06570_);
  and (_11431_, _11430_, _11428_);
  and (_11432_, _08534_, _07942_);
  or (_11433_, _11432_, _11363_);
  and (_11434_, _11433_, _06566_);
  or (_11435_, _11434_, _01324_);
  or (_11436_, _11435_, _11431_);
  or (_11437_, _01320_, \oc8051_golden_model_1.PCON [7]);
  and (_11438_, _11437_, _42355_);
  and (_40313_, _11438_, _11436_);
  not (_11439_, _07904_);
  and (_11440_, _11439_, \oc8051_golden_model_1.TMOD [7]);
  and (_11441_, _08536_, _07904_);
  or (_11442_, _11441_, _11440_);
  or (_11443_, _11442_, _06260_);
  and (_11444_, _08637_, _07904_);
  or (_11445_, _11444_, _11440_);
  or (_11446_, _11445_, _06286_);
  and (_11447_, _07904_, \oc8051_golden_model_1.ACC [7]);
  or (_11448_, _11447_, _11440_);
  and (_11449_, _11448_, _07143_);
  and (_11450_, _07144_, \oc8051_golden_model_1.TMOD [7]);
  or (_11451_, _11450_, _06285_);
  or (_11452_, _11451_, _11449_);
  and (_11453_, _11452_, _07169_);
  and (_11454_, _11453_, _11446_);
  and (_11455_, _11442_, _06354_);
  or (_11456_, _11455_, _11454_);
  and (_11457_, _11456_, _06346_);
  and (_11458_, _11448_, _06345_);
  or (_11459_, _11458_, _06259_);
  or (_11460_, _11459_, _11457_);
  and (_11461_, _11460_, _11443_);
  or (_11462_, _11461_, _09486_);
  and (_11463_, _08731_, _07904_);
  or (_11464_, _11440_, _06258_);
  or (_11465_, _11464_, _11463_);
  and (_11466_, _11465_, _06251_);
  and (_11467_, _11466_, _11462_);
  and (_11468_, _09004_, _07904_);
  or (_11469_, _11468_, _11440_);
  and (_11470_, _11469_, _05972_);
  or (_11471_, _11470_, _11467_);
  or (_11472_, _11471_, _10080_);
  and (_11473_, _09034_, _07904_);
  or (_11474_, _11440_, _09025_);
  or (_11475_, _11474_, _11473_);
  and (_11476_, _08806_, _07904_);
  or (_11477_, _11476_, _11440_);
  or (_11478_, _11477_, _06216_);
  and (_11479_, _11478_, _09030_);
  and (_11480_, _11479_, _11475_);
  and (_11481_, _11480_, _11472_);
  and (_11482_, _09042_, _07904_);
  or (_11483_, _11482_, _11440_);
  and (_11484_, _11483_, _06524_);
  or (_11485_, _11484_, _11481_);
  and (_11486_, _11485_, _07219_);
  or (_11487_, _11440_, _08026_);
  and (_11488_, _11477_, _06426_);
  and (_11489_, _11488_, _11487_);
  or (_11490_, _11489_, _11486_);
  and (_11491_, _11490_, _07217_);
  and (_11492_, _11448_, _06532_);
  and (_11493_, _11492_, _11487_);
  or (_11494_, _11493_, _06437_);
  or (_11495_, _11494_, _11491_);
  and (_11496_, _09033_, _07904_);
  or (_11497_, _11440_, _07229_);
  or (_11498_, _11497_, _11496_);
  and (_11499_, _11498_, _07231_);
  and (_11500_, _11499_, _11495_);
  nor (_11501_, _09041_, _11439_);
  or (_11502_, _11501_, _11440_);
  and (_11503_, _11502_, _06535_);
  or (_11504_, _11503_, _06559_);
  or (_11505_, _11504_, _11500_);
  or (_11506_, _11445_, _07240_);
  and (_11507_, _11506_, _06570_);
  and (_11508_, _11507_, _11505_);
  and (_11509_, _08534_, _07904_);
  or (_11510_, _11509_, _11440_);
  and (_11511_, _11510_, _06566_);
  or (_11512_, _11511_, _01324_);
  or (_11513_, _11512_, _11508_);
  or (_11514_, _01320_, \oc8051_golden_model_1.TMOD [7]);
  and (_11515_, _11514_, _42355_);
  and (_40314_, _11515_, _11513_);
  not (_11516_, \oc8051_golden_model_1.DPL [7]);
  nor (_11517_, _07950_, _11516_);
  and (_11518_, _08536_, _07950_);
  or (_11519_, _11518_, _11517_);
  or (_11520_, _11519_, _06260_);
  and (_11521_, _08637_, _07950_);
  or (_11522_, _11521_, _11517_);
  or (_11523_, _11522_, _06286_);
  and (_11524_, _07950_, \oc8051_golden_model_1.ACC [7]);
  or (_11525_, _11524_, _11517_);
  and (_11526_, _11525_, _07143_);
  nor (_11527_, _07143_, _11516_);
  or (_11528_, _11527_, _06285_);
  or (_11529_, _11528_, _11526_);
  and (_11530_, _11529_, _07169_);
  and (_11531_, _11530_, _11523_);
  and (_11532_, _11519_, _06354_);
  or (_11533_, _11532_, _06345_);
  or (_11534_, _11533_, _11531_);
  nor (_11535_, _05952_, _05935_);
  not (_11536_, _11535_);
  or (_11537_, _11525_, _06346_);
  and (_11538_, _11537_, _11536_);
  and (_11539_, _11538_, _11534_);
  and (_11540_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_11541_, _11540_, \oc8051_golden_model_1.DPL [2]);
  and (_11542_, _11541_, \oc8051_golden_model_1.DPL [3]);
  and (_11543_, _11542_, \oc8051_golden_model_1.DPL [4]);
  and (_11544_, _11543_, \oc8051_golden_model_1.DPL [5]);
  and (_11545_, _11544_, \oc8051_golden_model_1.DPL [6]);
  nor (_11546_, _11545_, \oc8051_golden_model_1.DPL [7]);
  and (_11547_, _11545_, \oc8051_golden_model_1.DPL [7]);
  nor (_11548_, _11547_, _11546_);
  and (_11549_, _11548_, _11535_);
  or (_11550_, _11549_, _11539_);
  and (_11551_, _11550_, _06396_);
  nor (_11552_, _08582_, _06396_);
  or (_11553_, _11552_, _06259_);
  or (_11554_, _11553_, _11551_);
  and (_11555_, _11554_, _11520_);
  or (_11556_, _11555_, _09486_);
  and (_11557_, _08731_, _07950_);
  or (_11558_, _11517_, _06258_);
  or (_11559_, _11558_, _11557_);
  and (_11560_, _11559_, _06251_);
  and (_11561_, _11560_, _11556_);
  and (_11562_, _09004_, _07950_);
  or (_11563_, _11562_, _11517_);
  and (_11564_, _11563_, _05972_);
  or (_11565_, _11564_, _11561_);
  or (_11566_, _11565_, _10080_);
  and (_11567_, _09034_, _07950_);
  or (_11568_, _11517_, _09025_);
  or (_11569_, _11568_, _11567_);
  and (_11570_, _08806_, _07950_);
  or (_11571_, _11570_, _11517_);
  or (_11572_, _11571_, _06216_);
  and (_11573_, _11572_, _09030_);
  and (_11574_, _11573_, _11569_);
  and (_11575_, _11574_, _11566_);
  and (_11576_, _09042_, _07950_);
  or (_11577_, _11576_, _11517_);
  and (_11578_, _11577_, _06524_);
  or (_11579_, _11578_, _11575_);
  and (_11580_, _11579_, _07219_);
  or (_11581_, _11517_, _08026_);
  and (_11582_, _11571_, _06426_);
  and (_11583_, _11582_, _11581_);
  or (_11584_, _11583_, _11580_);
  and (_11585_, _11584_, _07217_);
  and (_11586_, _11525_, _06532_);
  and (_11587_, _11586_, _11581_);
  or (_11588_, _11587_, _06437_);
  or (_11589_, _11588_, _11585_);
  and (_11590_, _09033_, _07950_);
  or (_11591_, _11517_, _07229_);
  or (_11592_, _11591_, _11590_);
  and (_11593_, _11592_, _07231_);
  and (_11594_, _11593_, _11589_);
  not (_11595_, _07950_);
  nor (_11596_, _09041_, _11595_);
  or (_11597_, _11596_, _11517_);
  and (_11598_, _11597_, _06535_);
  or (_11599_, _11598_, _06559_);
  or (_11600_, _11599_, _11594_);
  or (_11601_, _11522_, _07240_);
  and (_11602_, _11601_, _06570_);
  and (_11603_, _11602_, _11600_);
  and (_11604_, _08534_, _07950_);
  or (_11605_, _11604_, _11517_);
  and (_11606_, _11605_, _06566_);
  or (_11607_, _11606_, _01324_);
  or (_11608_, _11607_, _11603_);
  or (_11609_, _01320_, \oc8051_golden_model_1.DPL [7]);
  and (_11610_, _11609_, _42355_);
  and (_40315_, _11610_, _11608_);
  not (_11611_, \oc8051_golden_model_1.DPH [7]);
  nor (_11612_, _07953_, _11611_);
  and (_11613_, _08536_, _08261_);
  or (_11614_, _11613_, _11612_);
  or (_11615_, _11614_, _06260_);
  and (_11616_, _08637_, _08261_);
  or (_11617_, _11616_, _11612_);
  or (_11618_, _11617_, _06286_);
  and (_11619_, _07953_, \oc8051_golden_model_1.ACC [7]);
  or (_11620_, _11619_, _11612_);
  and (_11621_, _11620_, _07143_);
  nor (_11622_, _07143_, _11611_);
  or (_11623_, _11622_, _06285_);
  or (_11624_, _11623_, _11621_);
  and (_11625_, _11624_, _07169_);
  and (_11626_, _11625_, _11618_);
  and (_11627_, _11614_, _06354_);
  or (_11628_, _11627_, _06345_);
  or (_11629_, _11628_, _11626_);
  or (_11630_, _11620_, _06346_);
  and (_11631_, _11630_, _11536_);
  and (_11632_, _11631_, _11629_);
  and (_11633_, _11547_, \oc8051_golden_model_1.DPH [0]);
  and (_11634_, _11633_, \oc8051_golden_model_1.DPH [1]);
  and (_11635_, _11634_, \oc8051_golden_model_1.DPH [2]);
  and (_11636_, _11635_, \oc8051_golden_model_1.DPH [3]);
  and (_11637_, _11636_, \oc8051_golden_model_1.DPH [4]);
  and (_11638_, _11637_, \oc8051_golden_model_1.DPH [5]);
  and (_11639_, _11638_, \oc8051_golden_model_1.DPH [6]);
  nand (_11640_, _11639_, \oc8051_golden_model_1.DPH [7]);
  or (_11641_, _11639_, \oc8051_golden_model_1.DPH [7]);
  and (_11642_, _11641_, _11640_);
  and (_11643_, _11642_, _11535_);
  or (_11644_, _11643_, _11632_);
  and (_11645_, _11644_, _06396_);
  and (_11646_, _06395_, _06181_);
  or (_11647_, _11646_, _06259_);
  or (_11648_, _11647_, _11645_);
  and (_11649_, _11648_, _11615_);
  or (_11650_, _11649_, _09486_);
  or (_11651_, _11612_, _06258_);
  and (_11652_, _08731_, _07953_);
  or (_11653_, _11652_, _11651_);
  and (_11654_, _11653_, _06251_);
  and (_11655_, _11654_, _11650_);
  and (_11656_, _09004_, _07953_);
  or (_11657_, _11656_, _11612_);
  and (_11658_, _11657_, _05972_);
  or (_11659_, _11658_, _11655_);
  or (_11660_, _11659_, _10080_);
  and (_11661_, _09034_, _08261_);
  or (_11662_, _11612_, _09025_);
  or (_11663_, _11662_, _11661_);
  and (_11664_, _08806_, _07953_);
  or (_11665_, _11664_, _11612_);
  or (_11666_, _11665_, _06216_);
  and (_11667_, _11666_, _09030_);
  and (_11668_, _11667_, _11663_);
  and (_11669_, _11668_, _11660_);
  and (_11670_, _09042_, _08261_);
  or (_11671_, _11670_, _11612_);
  and (_11672_, _11671_, _06524_);
  or (_11673_, _11672_, _11669_);
  and (_11674_, _11673_, _07219_);
  or (_11675_, _11612_, _08026_);
  and (_11676_, _11665_, _06426_);
  and (_11677_, _11676_, _11675_);
  or (_11678_, _11677_, _11674_);
  and (_11679_, _11678_, _07217_);
  and (_11680_, _11620_, _06532_);
  and (_11681_, _11680_, _11675_);
  or (_11682_, _11681_, _06437_);
  or (_11683_, _11682_, _11679_);
  and (_11684_, _09033_, _08261_);
  or (_11685_, _11612_, _07229_);
  or (_11686_, _11685_, _11684_);
  and (_11687_, _11686_, _07231_);
  and (_11688_, _11687_, _11683_);
  not (_11689_, _08261_);
  nor (_11690_, _09041_, _11689_);
  or (_11691_, _11690_, _11612_);
  and (_11692_, _11691_, _06535_);
  or (_11693_, _11692_, _06559_);
  or (_11694_, _11693_, _11688_);
  or (_11695_, _11617_, _07240_);
  and (_11696_, _11695_, _06570_);
  and (_11697_, _11696_, _11694_);
  and (_11698_, _08534_, _08261_);
  or (_11699_, _11698_, _11612_);
  and (_11700_, _11699_, _06566_);
  or (_11701_, _11700_, _01324_);
  or (_11702_, _11701_, _11697_);
  or (_11703_, _01320_, \oc8051_golden_model_1.DPH [7]);
  and (_11704_, _11703_, _42355_);
  and (_40318_, _11704_, _11702_);
  not (_11705_, _07958_);
  and (_11706_, _11705_, \oc8051_golden_model_1.TL1 [7]);
  and (_11707_, _08637_, _07958_);
  or (_11708_, _11707_, _11706_);
  or (_11709_, _11708_, _06286_);
  and (_11710_, _07958_, \oc8051_golden_model_1.ACC [7]);
  or (_11711_, _11710_, _11706_);
  and (_11712_, _11711_, _07143_);
  and (_11713_, _07144_, \oc8051_golden_model_1.TL1 [7]);
  or (_11714_, _11713_, _06285_);
  or (_11715_, _11714_, _11712_);
  and (_11716_, _11715_, _07169_);
  and (_11717_, _11716_, _11709_);
  and (_11718_, _08536_, _07958_);
  or (_11719_, _11718_, _11706_);
  and (_11720_, _11719_, _06354_);
  or (_11721_, _11720_, _11717_);
  and (_11722_, _11721_, _06346_);
  and (_11723_, _11711_, _06345_);
  or (_11724_, _11723_, _06259_);
  or (_11725_, _11724_, _11722_);
  or (_11726_, _11719_, _06260_);
  and (_11727_, _11726_, _11725_);
  or (_11728_, _11727_, _09486_);
  and (_11729_, _08731_, _07958_);
  or (_11730_, _11706_, _06258_);
  or (_11731_, _11730_, _11729_);
  and (_11732_, _11731_, _06251_);
  and (_11733_, _11732_, _11728_);
  and (_11734_, _09004_, _07958_);
  or (_11735_, _11734_, _11706_);
  and (_11736_, _11735_, _05972_);
  or (_11737_, _11736_, _11733_);
  or (_11738_, _11737_, _10080_);
  and (_11739_, _09034_, _07958_);
  or (_11740_, _11706_, _09025_);
  or (_11741_, _11740_, _11739_);
  and (_11742_, _08806_, _07958_);
  or (_11743_, _11742_, _11706_);
  or (_11744_, _11743_, _06216_);
  and (_11745_, _11744_, _09030_);
  and (_11746_, _11745_, _11741_);
  and (_11747_, _11746_, _11738_);
  and (_11748_, _09042_, _07958_);
  or (_11749_, _11748_, _11706_);
  and (_11750_, _11749_, _06524_);
  or (_11751_, _11750_, _11747_);
  and (_11752_, _11751_, _07219_);
  or (_11753_, _11706_, _08026_);
  and (_11754_, _11743_, _06426_);
  and (_11755_, _11754_, _11753_);
  or (_11756_, _11755_, _11752_);
  and (_11757_, _11756_, _07217_);
  and (_11758_, _11711_, _06532_);
  and (_11759_, _11758_, _11753_);
  or (_11760_, _11759_, _06437_);
  or (_11761_, _11760_, _11757_);
  and (_11762_, _09033_, _07958_);
  or (_11763_, _11706_, _07229_);
  or (_11764_, _11763_, _11762_);
  and (_11765_, _11764_, _07231_);
  and (_11766_, _11765_, _11761_);
  nor (_11767_, _09041_, _11705_);
  or (_11768_, _11767_, _11706_);
  and (_11769_, _11768_, _06535_);
  or (_11770_, _11769_, _06559_);
  or (_11771_, _11770_, _11766_);
  or (_11772_, _11708_, _07240_);
  and (_11773_, _11772_, _06570_);
  and (_11774_, _11773_, _11771_);
  and (_11775_, _08534_, _07958_);
  or (_11776_, _11775_, _11706_);
  and (_11777_, _11776_, _06566_);
  or (_11778_, _11777_, _01324_);
  or (_11779_, _11778_, _11774_);
  or (_11780_, _01320_, \oc8051_golden_model_1.TL1 [7]);
  and (_11781_, _11780_, _42355_);
  and (_40319_, _11781_, _11779_);
  not (_11782_, _07912_);
  and (_11783_, _11782_, \oc8051_golden_model_1.TL0 [7]);
  and (_11784_, _08536_, _07912_);
  or (_11785_, _11784_, _11783_);
  or (_11786_, _11785_, _06260_);
  and (_11787_, _08637_, _07912_);
  or (_11788_, _11787_, _11783_);
  or (_11789_, _11788_, _06286_);
  and (_11790_, _07912_, \oc8051_golden_model_1.ACC [7]);
  or (_11791_, _11790_, _11783_);
  and (_11792_, _11791_, _07143_);
  and (_11793_, _07144_, \oc8051_golden_model_1.TL0 [7]);
  or (_11794_, _11793_, _06285_);
  or (_11795_, _11794_, _11792_);
  and (_11796_, _11795_, _07169_);
  and (_11797_, _11796_, _11789_);
  and (_11798_, _11785_, _06354_);
  or (_11799_, _11798_, _11797_);
  and (_11800_, _11799_, _06346_);
  and (_11801_, _11791_, _06345_);
  or (_11802_, _11801_, _06259_);
  or (_11803_, _11802_, _11800_);
  and (_11804_, _11803_, _11786_);
  or (_11805_, _11804_, _09486_);
  and (_11806_, _08731_, _07912_);
  or (_11807_, _11783_, _06258_);
  or (_11808_, _11807_, _11806_);
  and (_11809_, _11808_, _06251_);
  and (_11810_, _11809_, _11805_);
  and (_11811_, _09004_, _07912_);
  or (_11812_, _11811_, _11783_);
  and (_11813_, _11812_, _05972_);
  or (_11814_, _11813_, _11810_);
  or (_11815_, _11814_, _10080_);
  and (_11816_, _09034_, _07912_);
  or (_11817_, _11783_, _09025_);
  or (_11818_, _11817_, _11816_);
  and (_11819_, _08806_, _07912_);
  or (_11820_, _11819_, _11783_);
  or (_11821_, _11820_, _06216_);
  and (_11822_, _11821_, _09030_);
  and (_11823_, _11822_, _11818_);
  and (_11824_, _11823_, _11815_);
  and (_11825_, _09042_, _07912_);
  or (_11826_, _11825_, _11783_);
  and (_11827_, _11826_, _06524_);
  or (_11828_, _11827_, _11824_);
  and (_11829_, _11828_, _07219_);
  or (_11830_, _11783_, _08026_);
  and (_11831_, _11820_, _06426_);
  and (_11832_, _11831_, _11830_);
  or (_11833_, _11832_, _11829_);
  and (_11834_, _11833_, _07217_);
  and (_11835_, _11791_, _06532_);
  and (_11836_, _11835_, _11830_);
  or (_11837_, _11836_, _06437_);
  or (_11838_, _11837_, _11834_);
  and (_11839_, _09033_, _07912_);
  or (_11840_, _11783_, _07229_);
  or (_11841_, _11840_, _11839_);
  and (_11842_, _11841_, _07231_);
  and (_11843_, _11842_, _11838_);
  nor (_11844_, _09041_, _11782_);
  or (_11845_, _11844_, _11783_);
  and (_11846_, _11845_, _06535_);
  or (_11847_, _11846_, _06559_);
  or (_11848_, _11847_, _11843_);
  or (_11849_, _11788_, _07240_);
  and (_11850_, _11849_, _06570_);
  and (_11851_, _11850_, _11848_);
  and (_11852_, _08534_, _07912_);
  or (_11853_, _11852_, _11783_);
  and (_11854_, _11853_, _06566_);
  or (_11855_, _11854_, _01324_);
  or (_11856_, _11855_, _11851_);
  or (_11857_, _01320_, \oc8051_golden_model_1.TL0 [7]);
  and (_11858_, _11857_, _42355_);
  and (_40320_, _11858_, _11856_);
  and (_11859_, _01324_, \oc8051_golden_model_1.TCON [7]);
  not (_11860_, _07916_);
  and (_11861_, _11860_, \oc8051_golden_model_1.TCON [7]);
  and (_11862_, _08536_, _07916_);
  or (_11863_, _11862_, _11861_);
  or (_11864_, _11863_, _06260_);
  not (_11865_, _08600_);
  and (_11866_, _11865_, \oc8051_golden_model_1.TCON [7]);
  and (_11867_, _08622_, _08600_);
  or (_11868_, _11867_, _11866_);
  and (_11869_, _11868_, _06277_);
  and (_11870_, _08637_, _07916_);
  or (_11871_, _11870_, _11861_);
  or (_11872_, _11871_, _06286_);
  and (_11873_, _07916_, \oc8051_golden_model_1.ACC [7]);
  or (_11874_, _11873_, _11861_);
  and (_11875_, _11874_, _07143_);
  and (_11876_, _07144_, \oc8051_golden_model_1.TCON [7]);
  or (_11877_, _11876_, _06285_);
  or (_11878_, _11877_, _11875_);
  and (_11879_, _11878_, _06282_);
  and (_11880_, _11879_, _11872_);
  and (_11881_, _08626_, _08600_);
  or (_11882_, _11881_, _11866_);
  and (_11883_, _11882_, _06281_);
  or (_11884_, _11883_, _06354_);
  or (_11885_, _11884_, _11880_);
  or (_11886_, _11863_, _07169_);
  and (_11887_, _11886_, _11885_);
  or (_11888_, _11887_, _06345_);
  or (_11889_, _11874_, _06346_);
  and (_11890_, _11889_, _06278_);
  and (_11891_, _11890_, _11888_);
  or (_11892_, _11891_, _11869_);
  and (_11893_, _11892_, _06271_);
  and (_11894_, _08769_, _08600_);
  or (_11895_, _11894_, _11866_);
  and (_11896_, _11895_, _06270_);
  or (_11897_, _11896_, _11893_);
  and (_11898_, _11897_, _06267_);
  and (_11899_, _08789_, _08600_);
  or (_11900_, _11899_, _11866_);
  and (_11901_, _11900_, _06266_);
  or (_11902_, _11901_, _06259_);
  or (_11903_, _11902_, _11898_);
  and (_11904_, _11903_, _11864_);
  or (_11905_, _11904_, _09486_);
  and (_11906_, _08731_, _07916_);
  or (_11907_, _11861_, _06258_);
  or (_11908_, _11907_, _11906_);
  and (_11909_, _11908_, _06251_);
  and (_11910_, _11909_, _11905_);
  and (_11911_, _09004_, _07916_);
  or (_11912_, _11911_, _11861_);
  and (_11913_, _11912_, _05972_);
  or (_11914_, _11913_, _10080_);
  or (_11915_, _11914_, _11910_);
  and (_11916_, _09034_, _07916_);
  or (_11917_, _11861_, _09025_);
  or (_11918_, _11917_, _11916_);
  and (_11919_, _08806_, _07916_);
  or (_11920_, _11919_, _11861_);
  or (_11921_, _11920_, _06216_);
  and (_11922_, _11921_, _09030_);
  and (_11923_, _11922_, _11918_);
  and (_11924_, _11923_, _11915_);
  and (_11925_, _09042_, _07916_);
  or (_11926_, _11925_, _11861_);
  and (_11927_, _11926_, _06524_);
  or (_11928_, _11927_, _11924_);
  and (_11929_, _11928_, _07219_);
  or (_11930_, _11861_, _08026_);
  and (_11931_, _11920_, _06426_);
  and (_11932_, _11931_, _11930_);
  or (_11933_, _11932_, _11929_);
  and (_11934_, _11933_, _07217_);
  and (_11935_, _11874_, _06532_);
  and (_11936_, _11935_, _11930_);
  or (_11937_, _11936_, _06437_);
  or (_11938_, _11937_, _11934_);
  and (_11939_, _09033_, _07916_);
  or (_11940_, _11861_, _07229_);
  or (_11941_, _11940_, _11939_);
  and (_11942_, _11941_, _07231_);
  and (_11943_, _11942_, _11938_);
  nor (_11944_, _09041_, _11860_);
  or (_11945_, _11944_, _11861_);
  and (_11946_, _11945_, _06535_);
  or (_11947_, _11946_, _06559_);
  or (_11948_, _11947_, _11943_);
  or (_11949_, _11871_, _07240_);
  and (_11950_, _11949_, _05933_);
  and (_11951_, _11950_, _11948_);
  and (_11952_, _11868_, _05932_);
  or (_11953_, _11952_, _06566_);
  or (_11954_, _11953_, _11951_);
  and (_11955_, _08534_, _07916_);
  or (_11956_, _11861_, _06570_);
  or (_11957_, _11956_, _11955_);
  and (_11958_, _11957_, _01320_);
  and (_11959_, _11958_, _11954_);
  or (_11960_, _11959_, _11859_);
  and (_40321_, _11960_, _42355_);
  not (_11961_, _07900_);
  and (_11962_, _11961_, \oc8051_golden_model_1.TH1 [7]);
  and (_11963_, _08536_, _07900_);
  or (_11964_, _11963_, _11962_);
  or (_11965_, _11964_, _06260_);
  and (_11966_, _08637_, _07900_);
  or (_11967_, _11966_, _11962_);
  or (_11968_, _11967_, _06286_);
  and (_11969_, _07900_, \oc8051_golden_model_1.ACC [7]);
  or (_11970_, _11969_, _11962_);
  and (_11971_, _11970_, _07143_);
  and (_11972_, _07144_, \oc8051_golden_model_1.TH1 [7]);
  or (_11973_, _11972_, _06285_);
  or (_11974_, _11973_, _11971_);
  and (_11975_, _11974_, _07169_);
  and (_11976_, _11975_, _11968_);
  and (_11977_, _11964_, _06354_);
  or (_11978_, _11977_, _11976_);
  and (_11979_, _11978_, _06346_);
  and (_11980_, _11970_, _06345_);
  or (_11981_, _11980_, _06259_);
  or (_11982_, _11981_, _11979_);
  and (_11983_, _11982_, _11965_);
  or (_11984_, _11983_, _09486_);
  and (_11985_, _08731_, _07900_);
  or (_11986_, _11962_, _06258_);
  or (_11987_, _11986_, _11985_);
  and (_11988_, _11987_, _06251_);
  and (_11989_, _11988_, _11984_);
  and (_11990_, _09004_, _07900_);
  or (_11991_, _11990_, _11962_);
  and (_11992_, _11991_, _05972_);
  or (_11993_, _11992_, _11989_);
  or (_11994_, _11993_, _10080_);
  and (_11995_, _09034_, _07900_);
  or (_11996_, _11962_, _09025_);
  or (_11997_, _11996_, _11995_);
  nor (_11998_, _08582_, _11961_);
  or (_11999_, _11998_, _11962_);
  or (_12000_, _11999_, _06216_);
  and (_12001_, _12000_, _09030_);
  and (_12002_, _12001_, _11997_);
  and (_12003_, _12002_, _11994_);
  and (_12004_, _09042_, _07900_);
  or (_12005_, _12004_, _11962_);
  and (_12006_, _12005_, _06524_);
  or (_12007_, _12006_, _12003_);
  and (_12008_, _12007_, _07219_);
  or (_12009_, _11962_, _08026_);
  and (_12010_, _11999_, _06426_);
  and (_12011_, _12010_, _12009_);
  or (_12012_, _12011_, _12008_);
  and (_12013_, _12012_, _07217_);
  and (_12014_, _11970_, _06532_);
  and (_12015_, _12014_, _12009_);
  or (_12016_, _12015_, _06437_);
  or (_12017_, _12016_, _12013_);
  and (_12018_, _09033_, _07900_);
  or (_12019_, _11962_, _07229_);
  or (_12020_, _12019_, _12018_);
  and (_12021_, _12020_, _07231_);
  and (_12022_, _12021_, _12017_);
  nor (_12023_, _09041_, _11961_);
  or (_12024_, _12023_, _11962_);
  and (_12025_, _12024_, _06535_);
  or (_12026_, _12025_, _06559_);
  or (_12027_, _12026_, _12022_);
  or (_12028_, _11967_, _07240_);
  and (_12029_, _12028_, _06570_);
  and (_12030_, _12029_, _12027_);
  and (_12031_, _08534_, _07900_);
  or (_12032_, _12031_, _11962_);
  and (_12033_, _12032_, _06566_);
  or (_12034_, _12033_, _01324_);
  or (_12035_, _12034_, _12030_);
  or (_12036_, _01320_, \oc8051_golden_model_1.TH1 [7]);
  and (_12037_, _12036_, _42355_);
  and (_40322_, _12037_, _12035_);
  not (_12038_, _07908_);
  and (_12039_, _12038_, \oc8051_golden_model_1.TH0 [7]);
  and (_12040_, _08536_, _07908_);
  or (_12041_, _12040_, _12039_);
  or (_12042_, _12041_, _06260_);
  and (_12043_, _08637_, _07908_);
  or (_12044_, _12043_, _12039_);
  or (_12045_, _12044_, _06286_);
  and (_12046_, _07908_, \oc8051_golden_model_1.ACC [7]);
  or (_12047_, _12046_, _12039_);
  and (_12048_, _12047_, _07143_);
  and (_12049_, _07144_, \oc8051_golden_model_1.TH0 [7]);
  or (_12050_, _12049_, _06285_);
  or (_12051_, _12050_, _12048_);
  and (_12052_, _12051_, _07169_);
  and (_12053_, _12052_, _12045_);
  and (_12054_, _12041_, _06354_);
  or (_12055_, _12054_, _12053_);
  and (_12056_, _12055_, _06346_);
  and (_12057_, _12047_, _06345_);
  or (_12058_, _12057_, _06259_);
  or (_12059_, _12058_, _12056_);
  and (_12060_, _12059_, _12042_);
  or (_12061_, _12060_, _09486_);
  and (_12062_, _08731_, _07908_);
  or (_12063_, _12039_, _06258_);
  or (_12064_, _12063_, _12062_);
  and (_12065_, _12064_, _06251_);
  and (_12066_, _12065_, _12061_);
  and (_12067_, _09004_, _07908_);
  or (_12068_, _12067_, _12039_);
  and (_12069_, _12068_, _05972_);
  or (_12070_, _12069_, _12066_);
  or (_12071_, _12070_, _10080_);
  and (_12072_, _09034_, _07908_);
  or (_12073_, _12039_, _09025_);
  or (_12074_, _12073_, _12072_);
  and (_12075_, _08806_, _07908_);
  or (_12076_, _12075_, _12039_);
  or (_12077_, _12076_, _06216_);
  and (_12078_, _12077_, _09030_);
  and (_12079_, _12078_, _12074_);
  and (_12080_, _12079_, _12071_);
  and (_12081_, _09042_, _07908_);
  or (_12082_, _12081_, _12039_);
  and (_12083_, _12082_, _06524_);
  or (_12084_, _12083_, _12080_);
  and (_12085_, _12084_, _07219_);
  or (_12086_, _12039_, _08026_);
  and (_12087_, _12076_, _06426_);
  and (_12088_, _12087_, _12086_);
  or (_12089_, _12088_, _12085_);
  and (_12090_, _12089_, _07217_);
  and (_12091_, _12047_, _06532_);
  and (_12092_, _12091_, _12086_);
  or (_12093_, _12092_, _06437_);
  or (_12094_, _12093_, _12090_);
  and (_12095_, _09033_, _07908_);
  or (_12096_, _12039_, _07229_);
  or (_12097_, _12096_, _12095_);
  and (_12098_, _12097_, _07231_);
  and (_12099_, _12098_, _12094_);
  nor (_12100_, _09041_, _12038_);
  or (_12101_, _12100_, _12039_);
  and (_12102_, _12101_, _06535_);
  or (_12103_, _12102_, _06559_);
  or (_12104_, _12103_, _12099_);
  or (_12105_, _12044_, _07240_);
  and (_12106_, _12105_, _06570_);
  and (_12107_, _12106_, _12104_);
  and (_12108_, _08534_, _07908_);
  or (_12109_, _12108_, _12039_);
  and (_12110_, _12109_, _06566_);
  or (_12111_, _12110_, _01324_);
  or (_12112_, _12111_, _12107_);
  or (_12113_, _01320_, \oc8051_golden_model_1.TH0 [7]);
  and (_12114_, _12113_, _42355_);
  and (_40324_, _12114_, _12112_);
  nor (_12115_, _01320_, _09455_);
  not (_12116_, _05602_);
  and (_12117_, _08740_, _12116_);
  and (_12118_, _12117_, \oc8051_golden_model_1.PC [7]);
  and (_12119_, _12118_, \oc8051_golden_model_1.PC [8]);
  and (_12120_, _12119_, \oc8051_golden_model_1.PC [9]);
  and (_12121_, _12120_, \oc8051_golden_model_1.PC [10]);
  and (_12122_, _12121_, \oc8051_golden_model_1.PC [11]);
  and (_12123_, _12122_, \oc8051_golden_model_1.PC [12]);
  and (_12124_, _12123_, \oc8051_golden_model_1.PC [13]);
  nand (_12125_, _12124_, \oc8051_golden_model_1.PC [14]);
  nand (_12126_, _12125_, _09455_);
  or (_12127_, _12125_, _09455_);
  and (_12128_, _12127_, _12126_);
  and (_12129_, _11190_, _11185_);
  or (_12130_, _12129_, _12128_);
  and (_12131_, _08742_, \oc8051_golden_model_1.PC [8]);
  and (_12132_, _12131_, \oc8051_golden_model_1.PC [9]);
  and (_12133_, _12132_, \oc8051_golden_model_1.PC [10]);
  and (_12134_, _12133_, \oc8051_golden_model_1.PC [11]);
  and (_12135_, _12134_, \oc8051_golden_model_1.PC [12]);
  and (_12136_, _12135_, \oc8051_golden_model_1.PC [13]);
  and (_12137_, _12136_, \oc8051_golden_model_1.PC [14]);
  nor (_12138_, _12136_, \oc8051_golden_model_1.PC [14]);
  nor (_12139_, _12138_, _12137_);
  nand (_12140_, _12139_, _06181_);
  or (_12141_, _12139_, _06181_);
  and (_12142_, _12141_, _12140_);
  nor (_12143_, _12135_, \oc8051_golden_model_1.PC [13]);
  nor (_12144_, _12143_, _12136_);
  and (_12145_, _12144_, _06181_);
  nor (_12146_, _12144_, _06181_);
  nor (_12147_, _12134_, \oc8051_golden_model_1.PC [12]);
  nor (_12148_, _12147_, _12135_);
  nand (_12149_, _12148_, _06181_);
  nor (_12150_, _12133_, \oc8051_golden_model_1.PC [11]);
  nor (_12151_, _12150_, _12134_);
  and (_12152_, _12151_, _06181_);
  nor (_12153_, _12151_, _06181_);
  nor (_12154_, _12153_, _12152_);
  nor (_12155_, _12132_, \oc8051_golden_model_1.PC [10]);
  nor (_12156_, _12155_, _12133_);
  and (_12157_, _12156_, _06181_);
  nor (_12158_, _12156_, _06181_);
  nor (_12159_, _12158_, _12157_);
  and (_12160_, _12159_, _12154_);
  nor (_12161_, _12131_, \oc8051_golden_model_1.PC [9]);
  nor (_12162_, _12161_, _12132_);
  and (_12163_, _12162_, _06181_);
  nor (_12164_, _12162_, _06181_);
  nor (_12165_, _12164_, _12163_);
  not (_12166_, _12165_);
  and (_12167_, _08744_, _06181_);
  nor (_12168_, _08744_, _06181_);
  and (_12169_, _08739_, _06093_);
  nor (_12170_, _12169_, \oc8051_golden_model_1.PC [6]);
  nor (_12171_, _12170_, _08741_);
  not (_12172_, _12171_);
  or (_12173_, _12172_, _06325_);
  nand (_12174_, _12172_, _06325_);
  and (_12175_, _12174_, _12173_);
  and (_12176_, _06093_, \oc8051_golden_model_1.PC [4]);
  nor (_12177_, _12176_, \oc8051_golden_model_1.PC [5]);
  nor (_12178_, _12177_, _12169_);
  not (_12179_, _12178_);
  nor (_12180_, _12179_, _06604_);
  and (_12181_, _12179_, _06604_);
  nor (_12182_, _06093_, \oc8051_golden_model_1.PC [4]);
  nor (_12183_, _12182_, _12176_);
  nand (_12184_, _12183_, _07889_);
  nor (_12185_, _06212_, _06456_);
  and (_12186_, _06212_, _06456_);
  nor (_12187_, _06646_, _06451_);
  nor (_12188_, _06995_, \oc8051_golden_model_1.PC [1]);
  and (_12189_, _06248_, \oc8051_golden_model_1.PC [0]);
  and (_12190_, _06995_, \oc8051_golden_model_1.PC [1]);
  nor (_12191_, _12190_, _12188_);
  and (_12192_, _12191_, _12189_);
  nor (_12193_, _12192_, _12188_);
  not (_12194_, _12193_);
  and (_12195_, _06646_, _06451_);
  nor (_12196_, _12195_, _12187_);
  and (_12197_, _12196_, _12194_);
  nor (_12198_, _12197_, _12187_);
  nor (_12199_, _12198_, _12186_);
  or (_12200_, _12199_, _12185_);
  or (_12201_, _12183_, _07889_);
  and (_12202_, _12201_, _12184_);
  nand (_12203_, _12202_, _12200_);
  and (_12204_, _12203_, _12184_);
  nor (_12205_, _12204_, _12181_);
  or (_12206_, _12205_, _12180_);
  nand (_12207_, _12206_, _12175_);
  and (_12208_, _12207_, _12173_);
  nor (_12209_, _12208_, _12168_);
  or (_12210_, _12209_, _12167_);
  nor (_12211_, _08742_, \oc8051_golden_model_1.PC [8]);
  nor (_12212_, _12211_, _12131_);
  and (_12213_, _12212_, _06181_);
  nor (_12214_, _12212_, _06181_);
  nor (_12215_, _12214_, _12213_);
  nand (_12216_, _12215_, _12210_);
  nor (_12217_, _12216_, _12166_);
  and (_12218_, _12217_, _12160_);
  or (_12219_, _12213_, _12163_);
  and (_12220_, _12219_, _12160_);
  or (_12221_, _12157_, _12152_);
  or (_12222_, _12221_, _12220_);
  or (_12223_, _12222_, _12218_);
  or (_12224_, _12148_, _06181_);
  and (_12225_, _12224_, _12149_);
  nand (_12226_, _12225_, _12223_);
  and (_12227_, _12226_, _12149_);
  nor (_12228_, _12227_, _12146_);
  or (_12229_, _12228_, _12145_);
  nand (_12230_, _12229_, _12142_);
  and (_12231_, _12230_, _12140_);
  nor (_12232_, _09472_, _06181_);
  and (_12233_, _09472_, _06181_);
  nor (_12234_, _12233_, _12232_);
  and (_12235_, _12234_, _12231_);
  nor (_12236_, _12234_, _12231_);
  or (_12237_, _12236_, _12235_);
  or (_12238_, _12237_, _10774_);
  and (_12239_, _06007_, _05931_);
  or (_12240_, _09472_, \oc8051_golden_model_1.PSW [7]);
  and (_12241_, _12240_, _12239_);
  and (_12242_, _12241_, _12238_);
  nand (_12243_, _06012_, _05879_);
  and (_12244_, _12243_, _10964_);
  or (_12245_, _12244_, _12128_);
  or (_12246_, _12237_, _11327_);
  and (_12247_, _06003_, _05931_);
  not (_12248_, _11327_);
  or (_12249_, _12248_, _09472_);
  and (_12250_, _12249_, _12247_);
  and (_12251_, _12250_, _12246_);
  nor (_12252_, _09480_, _05984_);
  and (_12253_, _09465_, _05972_);
  nor (_12254_, _05945_, _05935_);
  not (_12255_, _12254_);
  and (_12256_, _09403_, \oc8051_golden_model_1.PC [8]);
  and (_12257_, _12256_, \oc8051_golden_model_1.PC [9]);
  and (_12258_, _12257_, \oc8051_golden_model_1.PC [10]);
  and (_12259_, _12258_, \oc8051_golden_model_1.PC [11]);
  and (_12260_, _12259_, \oc8051_golden_model_1.PC [12]);
  and (_12261_, _12260_, \oc8051_golden_model_1.PC [13]);
  nand (_12262_, _12261_, \oc8051_golden_model_1.PC [14]);
  or (_12263_, _12261_, \oc8051_golden_model_1.PC [14]);
  and (_12264_, _12263_, _12262_);
  nand (_12265_, _12264_, _08806_);
  or (_12266_, _12264_, _08806_);
  and (_12267_, _12266_, _12265_);
  nor (_12268_, _12260_, \oc8051_golden_model_1.PC [13]);
  nor (_12269_, _12268_, _12261_);
  and (_12270_, _12269_, _08806_);
  nor (_12271_, _12269_, _08806_);
  nor (_12272_, _12259_, \oc8051_golden_model_1.PC [12]);
  nor (_12273_, _12272_, _12260_);
  nand (_12274_, _12273_, _08806_);
  nor (_12275_, _12258_, \oc8051_golden_model_1.PC [11]);
  nor (_12276_, _12275_, _12259_);
  and (_12277_, _12276_, _08806_);
  nor (_12278_, _12276_, _08806_);
  nor (_12279_, _12278_, _12277_);
  nor (_12280_, _12257_, \oc8051_golden_model_1.PC [10]);
  nor (_12281_, _12280_, _12258_);
  and (_12282_, _12281_, _08806_);
  nor (_12283_, _12281_, _08806_);
  nor (_12284_, _12283_, _12282_);
  and (_12285_, _12284_, _12279_);
  nor (_12286_, _12256_, \oc8051_golden_model_1.PC [9]);
  nor (_12287_, _12286_, _12257_);
  and (_12288_, _12287_, _08806_);
  nor (_12289_, _12287_, _08806_);
  nor (_12290_, _12289_, _12288_);
  not (_12291_, _12290_);
  and (_12292_, _09405_, _08806_);
  nor (_12293_, _09405_, _08806_);
  and (_12294_, _09401_, _08739_);
  nor (_12295_, _12294_, \oc8051_golden_model_1.PC [6]);
  nor (_12296_, _12295_, _09402_);
  not (_12297_, _12296_);
  or (_12298_, _12297_, _08844_);
  nand (_12299_, _12297_, _08844_);
  and (_12300_, _12299_, _12298_);
  and (_12301_, _09401_, \oc8051_golden_model_1.PC [4]);
  nor (_12302_, _12301_, \oc8051_golden_model_1.PC [5]);
  nor (_12303_, _12302_, _12294_);
  and (_12304_, _12303_, _08913_);
  nor (_12305_, _12303_, _08913_);
  nor (_12306_, _09401_, \oc8051_golden_model_1.PC [4]);
  nor (_12307_, _12306_, _12301_);
  nand (_12308_, _12307_, _08919_);
  nor (_12309_, _09400_, \oc8051_golden_model_1.PC [3]);
  nor (_12310_, _12309_, _09401_);
  and (_12311_, _12310_, _08809_);
  nor (_12312_, _12310_, _08809_);
  nor (_12313_, _05625_, \oc8051_golden_model_1.PC [2]);
  nor (_12314_, _12313_, _09400_);
  and (_12315_, _12314_, _08980_);
  not (_12316_, _12315_);
  nor (_12317_, _07031_, _06035_);
  not (_12318_, _12317_);
  nor (_12319_, _06850_, \oc8051_golden_model_1.PC [0]);
  and (_12320_, _07031_, _06035_);
  nor (_12321_, _12320_, _12317_);
  nand (_12322_, _12321_, _12319_);
  and (_12323_, _12322_, _12318_);
  not (_12324_, _12323_);
  nor (_12325_, _12314_, _08980_);
  nor (_12326_, _12325_, _12315_);
  nand (_12327_, _12326_, _12324_);
  and (_12328_, _12327_, _12316_);
  nor (_12329_, _12328_, _12312_);
  or (_12330_, _12329_, _12311_);
  or (_12331_, _12307_, _08919_);
  and (_12332_, _12331_, _12308_);
  nand (_12333_, _12332_, _12330_);
  and (_12334_, _12333_, _12308_);
  nor (_12335_, _12334_, _12305_);
  or (_12336_, _12335_, _12304_);
  nand (_12337_, _12336_, _12300_);
  and (_12338_, _12337_, _12298_);
  nor (_12339_, _12338_, _12293_);
  or (_12340_, _12339_, _12292_);
  nor (_12341_, _09403_, \oc8051_golden_model_1.PC [8]);
  nor (_12342_, _12341_, _12256_);
  and (_12343_, _12342_, _08806_);
  nor (_12344_, _12342_, _08806_);
  nor (_12345_, _12344_, _12343_);
  nand (_12346_, _12345_, _12340_);
  nor (_12347_, _12346_, _12291_);
  and (_12348_, _12347_, _12285_);
  or (_12349_, _12343_, _12288_);
  and (_12350_, _12349_, _12285_);
  or (_12351_, _12282_, _12277_);
  or (_12352_, _12351_, _12350_);
  or (_12353_, _12352_, _12348_);
  or (_12354_, _12273_, _08806_);
  and (_12355_, _12354_, _12274_);
  nand (_12356_, _12355_, _12353_);
  and (_12357_, _12356_, _12274_);
  nor (_12358_, _12357_, _12271_);
  or (_12359_, _12358_, _12270_);
  nand (_12360_, _12359_, _12267_);
  and (_12361_, _12360_, _12265_);
  not (_12362_, _09465_);
  and (_12363_, _12362_, _08582_);
  nor (_12364_, _12362_, _08582_);
  nor (_12365_, _12364_, _12363_);
  and (_12366_, _12365_, _12361_);
  nor (_12367_, _12365_, _12361_);
  nor (_12368_, _12367_, _12366_);
  or (_12369_, _09247_, _06212_);
  nand (_12370_, _09247_, _06212_);
  and (_12371_, _12370_, _12369_);
  and (_12372_, _09293_, _06646_);
  nor (_12373_, _09293_, _06646_);
  nor (_12374_, _12373_, _12372_);
  and (_12375_, _12374_, _12371_);
  nand (_12376_, _09384_, _06250_);
  nor (_12377_, _09339_, _06995_);
  and (_12378_, _09339_, _06995_);
  nor (_12379_, _12378_, _12377_);
  and (_12380_, _12379_, _12376_);
  and (_12381_, _12380_, _12375_);
  or (_12382_, _09384_, _06250_);
  and (_12383_, _09067_, _06181_);
  nor (_12384_, _12383_, _08781_);
  or (_12385_, _09435_, _06325_);
  or (_12386_, _09112_, _07589_);
  and (_12387_, _12386_, _12385_);
  and (_12388_, _12387_, _12384_);
  or (_12389_, _09157_, _07873_);
  or (_12390_, _09436_, _06604_);
  and (_12391_, _12390_, _12389_);
  or (_12392_, _09202_, _07889_);
  or (_12393_, _09437_, _06961_);
  and (_12394_, _12393_, _12392_);
  and (_12395_, _12394_, _12391_);
  and (_12396_, _12395_, _12388_);
  and (_12397_, _12396_, _12382_);
  nand (_12398_, _12397_, _12381_);
  and (_12399_, _12398_, _12368_);
  and (_12400_, _12397_, _12381_);
  and (_12401_, _12400_, _12362_);
  or (_12402_, _12401_, _06424_);
  nor (_12403_, _12402_, _12399_);
  nor (_12404_, _10622_, _07174_);
  or (_12405_, _12404_, _12128_);
  and (_12406_, _06361_, _05949_);
  not (_12407_, _12406_);
  nor (_12408_, _05948_, _05935_);
  nor (_12409_, _12408_, _10656_);
  not (_12410_, _12409_);
  nor (_12411_, _12410_, _07159_);
  or (_12412_, _12411_, _12128_);
  not (_12413_, _12368_);
  and (_12414_, _08374_, _08324_);
  and (_12415_, _08631_, _12414_);
  and (_12416_, _08127_, _08025_);
  and (_12417_, _12416_, _08628_);
  and (_12418_, _12417_, _12415_);
  or (_12419_, _12418_, _12413_);
  nand (_12420_, _12417_, _12415_);
  or (_12421_, _12420_, _09465_);
  and (_12422_, _12421_, _12419_);
  or (_12423_, _12422_, _06286_);
  or (_12424_, _09420_, _09419_);
  or (_12425_, _09418_, _08536_);
  nor (_12426_, _12425_, _12424_);
  or (_12427_, _08662_, _09421_);
  or (_12428_, _09422_, _07157_);
  nor (_12429_, _12428_, _12427_);
  and (_12430_, _12429_, _12426_);
  and (_12431_, _12430_, _09472_);
  nand (_12432_, _12429_, _12426_);
  and (_12433_, _12432_, _12237_);
  or (_12434_, _12433_, _12431_);
  and (_12435_, _12434_, _08734_);
  and (_12436_, _12128_, _06755_);
  and (_12437_, _12128_, _07455_);
  nor (_12438_, _06755_, _09455_);
  and (_12439_, _12438_, _07454_);
  or (_12440_, _12439_, _12437_);
  and (_12441_, _12440_, _07144_);
  or (_12442_, _12441_, _12436_);
  and (_12443_, _12442_, _07858_);
  nor (_12444_, _07137_, _05959_);
  nor (_12445_, _12444_, _10643_);
  and (_12446_, _12445_, _10641_);
  not (_12447_, _12446_);
  or (_12448_, _12447_, _10642_);
  or (_12449_, _07143_, _07152_);
  and (_12450_, _12449_, _09472_);
  or (_12451_, _12450_, _12448_);
  or (_12452_, _12451_, _12443_);
  not (_12453_, _12448_);
  or (_12454_, _12453_, _12128_);
  and (_12455_, _12454_, _08736_);
  nand (_12456_, _12455_, _12452_);
  nor (_12457_, _07159_, _06285_);
  nand (_12458_, _12457_, _12456_);
  or (_12459_, _12458_, _12435_);
  and (_12460_, _12459_, _12423_);
  nand (_12461_, _12409_, _12404_);
  or (_12462_, _12461_, _12460_);
  and (_12463_, _12462_, _12412_);
  or (_12464_, _12463_, _12407_);
  and (_12465_, _12464_, _12405_);
  or (_12466_, _12465_, _06345_);
  nor (_12467_, _05954_, _05935_);
  nor (_12468_, _12467_, _10696_);
  and (_12469_, _12406_, _06346_);
  or (_12470_, _12469_, _09472_);
  and (_12471_, _12470_, _12468_);
  and (_12472_, _12471_, _12466_);
  not (_12473_, _12468_);
  and (_12474_, _12473_, _12128_);
  not (_12475_, _05955_);
  nor (_12476_, _06276_, _12475_);
  and (_12477_, _12476_, _06278_);
  not (_12478_, _12477_);
  or (_12479_, _12478_, _12474_);
  or (_12480_, _12479_, _12472_);
  or (_12481_, _12477_, _09472_);
  and (_12482_, _12481_, _12480_);
  nor (_12483_, _07509_, _05945_);
  nor (_12484_, _12483_, _06415_);
  not (_12485_, _12484_);
  or (_12486_, _12485_, _12482_);
  and (_12487_, _07578_, _06356_);
  and (_12488_, _09421_, _06212_);
  nor (_12489_, _12488_, _12487_);
  and (_12490_, _07760_, _06647_);
  and (_12491_, _08662_, _06646_);
  nor (_12492_, _12491_, _12490_);
  and (_12493_, _12492_, _12489_);
  and (_12494_, _07135_, _06250_);
  not (_12495_, _12494_);
  and (_12496_, _09422_, _06995_);
  and (_12497_, _07334_, _06996_);
  nor (_12498_, _12497_, _12496_);
  and (_12499_, _12498_, _12495_);
  and (_12500_, _12499_, _12493_);
  and (_12501_, _07157_, _06248_);
  not (_12502_, _12501_);
  not (_12503_, _08024_);
  and (_12504_, _08023_, _06181_);
  nor (_12505_, _12504_, _12503_);
  and (_12506_, _09418_, _06325_);
  and (_12507_, _08125_, _07589_);
  nor (_12508_, _12507_, _12506_);
  and (_12509_, _12508_, _12505_);
  and (_12510_, _08228_, _07873_);
  and (_12511_, _09419_, _06604_);
  nor (_12512_, _12511_, _12510_);
  and (_12513_, _08525_, _07889_);
  and (_12514_, _09420_, _06961_);
  nor (_12515_, _12514_, _12513_);
  and (_12516_, _12515_, _12512_);
  and (_12517_, _12516_, _12509_);
  and (_12518_, _12517_, _12502_);
  and (_12519_, _12518_, _12500_);
  and (_12520_, _12519_, _09465_);
  nor (_12521_, _12519_, _12368_);
  or (_12522_, _12521_, _12520_);
  or (_12523_, _12522_, _12484_);
  and (_12524_, _12523_, _06424_);
  and (_12525_, _12524_, _12486_);
  or (_12526_, _12525_, _06347_);
  or (_12527_, _12526_, _12403_);
  not (_12528_, _06419_);
  nor (_12529_, _11246_, _11247_);
  nor (_12530_, _12529_, _11250_);
  not (_12531_, _11253_);
  nor (_12532_, _08374_, \oc8051_golden_model_1.ACC [0]);
  or (_12533_, _12532_, _11254_);
  and (_12534_, _12533_, _12531_);
  and (_12535_, _12534_, _12530_);
  nor (_12536_, _11241_, _11240_);
  nor (_12537_, _12536_, _11245_);
  nor (_12538_, _11239_, _09042_);
  and (_12539_, _12538_, _12537_);
  and (_12540_, _12539_, _12535_);
  nand (_12541_, _12540_, _09465_);
  or (_12542_, _12540_, _12368_);
  and (_12543_, _12542_, _06347_);
  nand (_12544_, _12543_, _12541_);
  and (_12545_, _12544_, _12528_);
  and (_12546_, _12545_, _12527_);
  nor (_12547_, _06212_, \oc8051_golden_model_1.ACC [3]);
  and (_12548_, _06212_, \oc8051_golden_model_1.ACC [3]);
  nor (_12549_, _12548_, _12547_);
  and (_12550_, _12549_, _11289_);
  nor (_12551_, _06248_, \oc8051_golden_model_1.ACC [0]);
  nor (_12552_, _12551_, _11293_);
  nor (_12553_, _12552_, _11292_);
  and (_12554_, _12553_, _12550_);
  nor (_12555_, _11277_, _11278_);
  nor (_12556_, _12555_, _11283_);
  nor (_12557_, _11276_, _10934_);
  and (_12558_, _12557_, _12556_);
  and (_12559_, _12558_, _12554_);
  not (_12560_, _12559_);
  nand (_12561_, _12560_, _12368_);
  nand (_12562_, _12559_, _12362_);
  and (_12563_, _12562_, _06419_);
  and (_12564_, _12563_, _12561_);
  or (_12565_, _12564_, _12546_);
  and (_12566_, _12565_, _12255_);
  nand (_12567_, _12254_, _12128_);
  not (_12568_, _07373_);
  and (_12569_, _06702_, _06336_);
  nor (_12570_, _12569_, _06368_);
  and (_12571_, _12570_, _08650_);
  and (_12572_, _12571_, _12568_);
  nor (_12573_, _07374_, _07458_);
  not (_12574_, _07435_);
  and (_12575_, _06407_, _06336_);
  nor (_12576_, _12575_, _06270_);
  and (_12577_, _12576_, _12574_);
  and (_12578_, _12577_, _12573_);
  and (_12579_, _12578_, _12572_);
  nand (_12580_, _12579_, _12567_);
  or (_12581_, _12580_, _12566_);
  and (_12582_, _05970_, _06336_);
  not (_12583_, _12582_);
  nor (_12584_, _11535_, _09520_);
  and (_12585_, _12584_, _12583_);
  or (_12586_, _12579_, _09472_);
  and (_12587_, _12586_, _12585_);
  and (_12588_, _12587_, _12581_);
  not (_12589_, _12585_);
  and (_12590_, _12589_, _12128_);
  and (_12591_, _06372_, _05953_);
  not (_12592_, _12591_);
  or (_12593_, _12592_, _12590_);
  or (_12594_, _12593_, _12588_);
  and (_12595_, _10724_, _10555_);
  or (_12596_, _12591_, _09472_);
  and (_12597_, _12596_, _12595_);
  and (_12598_, _12597_, _12594_);
  nor (_12599_, _10486_, _06380_);
  not (_12600_, _12599_);
  not (_12601_, _12595_);
  and (_12602_, _12601_, _12128_);
  or (_12603_, _12602_, _12600_);
  or (_12604_, _12603_, _12598_);
  or (_12605_, _12599_, _09472_);
  and (_12606_, _12605_, _05940_);
  and (_12607_, _12606_, _12604_);
  and (_12608_, _12128_, _05976_);
  nor (_12609_, _06266_, _05974_);
  not (_12610_, _12609_);
  or (_12611_, _12610_, _12608_);
  or (_12612_, _12611_, _12607_);
  or (_12613_, _12609_, _09472_);
  and (_12614_, _12613_, _06396_);
  and (_12615_, _12614_, _12612_);
  nand (_12616_, _09465_, _06395_);
  nand (_12617_, _12616_, _06261_);
  or (_12618_, _12617_, _12615_);
  or (_12619_, _09472_, _06261_);
  and (_12620_, _12619_, _06251_);
  and (_12621_, _12620_, _12618_);
  or (_12622_, _12621_, _12253_);
  and (_12623_, _12622_, _12252_);
  nor (_12624_, _06330_, _05997_);
  not (_12625_, _12624_);
  not (_12626_, _12252_);
  and (_12627_, _12626_, _12128_);
  or (_12628_, _12627_, _12625_);
  or (_12629_, _12628_, _12623_);
  and (_12630_, _05971_, _05931_);
  not (_12631_, _12630_);
  or (_12632_, _12624_, _09472_);
  and (_12633_, _12632_, _12631_);
  and (_12634_, _12633_, _12629_);
  and (_12635_, _12630_, _12237_);
  or (_12636_, _12635_, _09016_);
  or (_12637_, _12636_, _12634_);
  or (_12638_, _09472_, _09015_);
  and (_12639_, _12638_, _06216_);
  and (_12640_, _12639_, _12637_);
  and (_12641_, _09465_, _06215_);
  or (_12642_, _12641_, _10891_);
  or (_12643_, _12642_, _12640_);
  and (_12644_, _06003_, _06397_);
  and (_12645_, _10891_, _09473_);
  nor (_12646_, _12645_, _12644_);
  and (_12647_, _12646_, _12643_);
  and (_12648_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_12649_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nand (_12650_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  or (_12651_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  and (_12652_, _12651_, _12650_);
  and (_12653_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12654_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_12655_, _12654_, _12653_);
  nand (_12656_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  or (_12657_, _06113_, _06109_);
  or (_12658_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  and (_12659_, _12658_, _12656_);
  nand (_12660_, _12659_, _12657_);
  and (_12661_, _12660_, _12656_);
  not (_12662_, _12661_);
  and (_12663_, _12662_, _12655_);
  or (_12664_, _12663_, _12653_);
  nand (_12665_, _12664_, _12652_);
  and (_12666_, _12665_, _12650_);
  nor (_12667_, _12666_, _12649_);
  or (_12668_, _12667_, _12648_);
  and (_12669_, _12668_, \oc8051_golden_model_1.DPH [0]);
  and (_12670_, _12669_, \oc8051_golden_model_1.DPH [1]);
  and (_12671_, _12670_, \oc8051_golden_model_1.DPH [2]);
  and (_12672_, _12671_, \oc8051_golden_model_1.DPH [3]);
  and (_12673_, _12672_, \oc8051_golden_model_1.DPH [4]);
  and (_12674_, _12673_, \oc8051_golden_model_1.DPH [5]);
  and (_12675_, _12674_, \oc8051_golden_model_1.DPH [6]);
  nand (_12676_, _12675_, \oc8051_golden_model_1.DPH [7]);
  or (_12677_, _12675_, \oc8051_golden_model_1.DPH [7]);
  and (_12678_, _12677_, _12644_);
  and (_12679_, _12678_, _12676_);
  nor (_12680_, _06329_, _06004_);
  not (_12681_, _12680_);
  or (_12683_, _12681_, _12679_);
  or (_12684_, _12683_, _12647_);
  not (_12685_, _12247_);
  or (_12686_, _12680_, _09472_);
  and (_12687_, _12686_, _12685_);
  and (_12688_, _12687_, _12684_);
  or (_12689_, _12688_, _12251_);
  nor (_12690_, _09012_, _10907_);
  not (_12691_, _12690_);
  and (_12692_, _09006_, _06000_);
  nor (_12693_, _12692_, _10908_);
  and (_12694_, _12693_, _10905_);
  and (_12695_, _12694_, _12691_);
  and (_12696_, _12695_, _12689_);
  not (_12697_, _12695_);
  and (_12698_, _12697_, _12128_);
  nor (_12699_, _10481_, _06526_);
  not (_12700_, _12699_);
  or (_12701_, _12700_, _12698_);
  or (_12702_, _12701_, _12696_);
  or (_12704_, _12699_, _09472_);
  and (_12705_, _12704_, _09025_);
  and (_12706_, _12705_, _12702_);
  nand (_12707_, _09465_, _06398_);
  nor (_12708_, _06524_, _06001_);
  nand (_12709_, _12708_, _12707_);
  or (_12710_, _12709_, _12706_);
  and (_12711_, _06000_, _05931_);
  not (_12712_, _12711_);
  or (_12713_, _12708_, _09472_);
  and (_12714_, _12713_, _12712_);
  and (_12715_, _12714_, _12710_);
  or (_12716_, _12237_, _12248_);
  or (_12717_, _11327_, _09472_);
  and (_12718_, _12717_, _12711_);
  and (_12719_, _12718_, _12716_);
  not (_12720_, _12244_);
  or (_12721_, _12720_, _12719_);
  or (_12722_, _12721_, _12715_);
  and (_12723_, _12722_, _12245_);
  or (_12724_, _12723_, _10970_);
  or (_12725_, _10969_, _09472_);
  and (_12726_, _12725_, _07219_);
  and (_12727_, _12726_, _12724_);
  nand (_12728_, _09465_, _06426_);
  nor (_12729_, _06532_, _06013_);
  nand (_12730_, _12729_, _12728_);
  or (_12731_, _12730_, _12727_);
  and (_12732_, _06012_, _05931_);
  not (_12733_, _12732_);
  or (_12734_, _12729_, _09472_);
  and (_12735_, _12734_, _12733_);
  and (_12736_, _12735_, _12731_);
  or (_12737_, _12237_, \oc8051_golden_model_1.PSW [7]);
  or (_12738_, _09472_, _10774_);
  and (_12739_, _12738_, _12732_);
  and (_12740_, _12739_, _12737_);
  or (_12741_, _12740_, _12736_);
  nor (_12742_, _06256_, _06801_);
  nor (_12743_, _12742_, _07059_);
  nor (_12744_, _12743_, _06884_);
  and (_12745_, _07466_, _06007_);
  not (_12746_, _12745_);
  nor (_12747_, _10989_, _10984_);
  and (_12748_, _12747_, _12746_);
  and (_12749_, _12748_, _12744_);
  and (_12750_, _12749_, _12741_);
  not (_12751_, _12749_);
  and (_12752_, _12751_, _12128_);
  or (_12753_, _12752_, _11008_);
  or (_12754_, _12753_, _12750_);
  or (_12755_, _11007_, _09472_);
  and (_12756_, _12755_, _07229_);
  and (_12757_, _12756_, _12754_);
  nand (_12758_, _09465_, _06437_);
  nor (_12759_, _06535_, _06008_);
  nand (_12760_, _12759_, _12758_);
  or (_12761_, _12760_, _12757_);
  not (_12762_, _12239_);
  or (_12763_, _12759_, _09472_);
  and (_12764_, _12763_, _12762_);
  and (_12765_, _12764_, _12761_);
  or (_12766_, _12765_, _12242_);
  and (_12767_, _11027_, _11023_);
  and (_12768_, _12767_, _12766_);
  nor (_12769_, _11082_, _06522_);
  not (_12770_, _12769_);
  not (_12771_, _12767_);
  and (_12772_, _12771_, _12128_);
  or (_12773_, _12772_, _12770_);
  or (_12774_, _12773_, _12768_);
  not (_12775_, _11111_);
  or (_12776_, _12769_, _09472_);
  and (_12777_, _12776_, _12775_);
  and (_12778_, _12777_, _12774_);
  and (_12779_, _12128_, _11111_);
  or (_12780_, _12779_, _06543_);
  or (_12781_, _12780_, _12778_);
  not (_12782_, _06543_);
  or (_12783_, _08536_, _12782_);
  and (_12784_, _12783_, _12781_);
  or (_12785_, _12784_, _06011_);
  not (_12786_, _06436_);
  nand (_12787_, _09473_, _06011_);
  and (_12788_, _12787_, _12786_);
  and (_12789_, _12788_, _12785_);
  not (_12790_, _12129_);
  not (_12791_, _07949_);
  and (_12792_, _08607_, \oc8051_golden_model_1.P3 [2]);
  and (_12793_, _08609_, \oc8051_golden_model_1.IE [2]);
  nor (_12794_, _12793_, _12792_);
  and (_12795_, _08612_, \oc8051_golden_model_1.SCON [2]);
  and (_12796_, _08614_, \oc8051_golden_model_1.P2 [2]);
  nor (_12797_, _12796_, _12795_);
  and (_12798_, _12797_, _12794_);
  and (_12799_, _08589_, \oc8051_golden_model_1.IP [2]);
  and (_12800_, _08592_, \oc8051_golden_model_1.PSW [2]);
  and (_12801_, _08596_, \oc8051_golden_model_1.ACC [2]);
  and (_12802_, _08594_, \oc8051_golden_model_1.B [2]);
  or (_12803_, _12802_, _12801_);
  or (_12804_, _12803_, _12800_);
  nor (_12805_, _12804_, _12799_);
  and (_12806_, _08600_, \oc8051_golden_model_1.TCON [2]);
  and (_12807_, _07939_, \oc8051_golden_model_1.P0 [2]);
  and (_12808_, _08603_, \oc8051_golden_model_1.P1 [2]);
  or (_12809_, _12808_, _12807_);
  nor (_12810_, _12809_, _12806_);
  and (_12811_, _12810_, _12805_);
  and (_12812_, _12811_, _12798_);
  and (_12813_, _12812_, _08422_);
  nor (_12814_, _12813_, _12791_);
  not (_12815_, _08255_);
  and (_12816_, _07939_, \oc8051_golden_model_1.P0 [1]);
  and (_12817_, _08600_, \oc8051_golden_model_1.TCON [1]);
  and (_12818_, _08603_, \oc8051_golden_model_1.P1 [1]);
  and (_12819_, _08612_, \oc8051_golden_model_1.SCON [1]);
  and (_12820_, _08614_, \oc8051_golden_model_1.P2 [1]);
  and (_12821_, _08609_, \oc8051_golden_model_1.IE [1]);
  and (_12822_, _08607_, \oc8051_golden_model_1.P3 [1]);
  and (_12823_, _08589_, \oc8051_golden_model_1.IP [1]);
  and (_12824_, _08592_, \oc8051_golden_model_1.PSW [1]);
  and (_12825_, _08594_, \oc8051_golden_model_1.B [1]);
  and (_12826_, _08596_, \oc8051_golden_model_1.ACC [1]);
  or (_12827_, _12826_, _12825_);
  or (_12828_, _12827_, _12824_);
  or (_12829_, _12828_, _12823_);
  or (_12830_, _12829_, _12822_);
  or (_12831_, _12830_, _12821_);
  or (_12832_, _12831_, _12820_);
  or (_12833_, _12832_, _12819_);
  or (_12834_, _12833_, _12818_);
  or (_12835_, _12834_, _12817_);
  nor (_12836_, _12835_, _12816_);
  and (_12837_, _12836_, _08323_);
  nor (_12838_, _12837_, _12815_);
  nor (_12839_, _12838_, _12814_);
  and (_12840_, _08589_, \oc8051_golden_model_1.IP [4]);
  and (_12841_, _08614_, \oc8051_golden_model_1.P2 [4]);
  nor (_12842_, _12841_, _12840_);
  and (_12843_, _08592_, \oc8051_golden_model_1.PSW [4]);
  and (_12844_, _08596_, \oc8051_golden_model_1.ACC [4]);
  and (_12845_, _08594_, \oc8051_golden_model_1.B [4]);
  or (_12846_, _12845_, _12844_);
  nor (_12847_, _12846_, _12843_);
  and (_12848_, _08600_, \oc8051_golden_model_1.TCON [4]);
  and (_12849_, _07939_, \oc8051_golden_model_1.P0 [4]);
  and (_12850_, _08603_, \oc8051_golden_model_1.P1 [4]);
  or (_12851_, _12850_, _12849_);
  nor (_12852_, _12851_, _12848_);
  and (_12853_, _08612_, \oc8051_golden_model_1.SCON [4]);
  and (_12854_, _08609_, \oc8051_golden_model_1.IE [4]);
  and (_12855_, _08607_, \oc8051_golden_model_1.P3 [4]);
  or (_12856_, _12855_, _12854_);
  nor (_12857_, _12856_, _12853_);
  and (_12858_, _12857_, _12852_);
  and (_12859_, _12858_, _12847_);
  and (_12860_, _12859_, _12842_);
  and (_12861_, _12860_, _08526_);
  and (_12862_, _07869_, _06647_);
  not (_12863_, _12862_);
  nor (_12864_, _12863_, _12861_);
  nor (_12865_, _12864_, _08767_);
  and (_12866_, _12865_, _12839_);
  and (_12867_, _07869_, _06646_);
  not (_12868_, _12867_);
  and (_12869_, _08589_, \oc8051_golden_model_1.IP [0]);
  and (_12870_, _08612_, \oc8051_golden_model_1.SCON [0]);
  nor (_12871_, _12870_, _12869_);
  and (_12872_, _08592_, \oc8051_golden_model_1.PSW [0]);
  and (_12873_, _08596_, \oc8051_golden_model_1.ACC [0]);
  and (_12874_, _08594_, \oc8051_golden_model_1.B [0]);
  or (_12875_, _12874_, _12873_);
  nor (_12876_, _12875_, _12872_);
  and (_12877_, _08600_, \oc8051_golden_model_1.TCON [0]);
  and (_12878_, _07939_, \oc8051_golden_model_1.P0 [0]);
  and (_12879_, _08603_, \oc8051_golden_model_1.P1 [0]);
  or (_12880_, _12879_, _12878_);
  nor (_12881_, _12880_, _12877_);
  and (_12882_, _08614_, \oc8051_golden_model_1.P2 [0]);
  and (_12883_, _08609_, \oc8051_golden_model_1.IE [0]);
  and (_12884_, _08607_, \oc8051_golden_model_1.P3 [0]);
  or (_12885_, _12884_, _12883_);
  nor (_12886_, _12885_, _12882_);
  and (_12887_, _12886_, _12881_);
  and (_12888_, _12887_, _12876_);
  and (_12889_, _12888_, _12871_);
  not (_12890_, _12889_);
  nor (_12891_, _12890_, _08373_);
  nor (_12892_, _12891_, _12868_);
  and (_12893_, _08592_, \oc8051_golden_model_1.PSW [6]);
  and (_12894_, _08614_, \oc8051_golden_model_1.P2 [6]);
  nor (_12895_, _12894_, _12893_);
  and (_12896_, _08589_, \oc8051_golden_model_1.IP [6]);
  and (_12897_, _08596_, \oc8051_golden_model_1.ACC [6]);
  and (_12898_, _08594_, \oc8051_golden_model_1.B [6]);
  or (_12899_, _12898_, _12897_);
  nor (_12900_, _12899_, _12896_);
  and (_12901_, _08600_, \oc8051_golden_model_1.TCON [6]);
  and (_12902_, _08603_, \oc8051_golden_model_1.P1 [6]);
  and (_12903_, _07939_, \oc8051_golden_model_1.P0 [6]);
  or (_12904_, _12903_, _12902_);
  nor (_12905_, _12904_, _12901_);
  and (_12906_, _08612_, \oc8051_golden_model_1.SCON [6]);
  and (_12907_, _08609_, \oc8051_golden_model_1.IE [6]);
  and (_12908_, _08607_, \oc8051_golden_model_1.P3 [6]);
  or (_12909_, _12908_, _12907_);
  nor (_12910_, _12909_, _12906_);
  and (_12911_, _12910_, _12905_);
  and (_12912_, _12911_, _12900_);
  and (_12913_, _12912_, _12895_);
  and (_12914_, _12913_, _08126_);
  and (_12915_, _07910_, _06647_);
  not (_12916_, _12915_);
  nor (_12917_, _12916_, _12914_);
  nor (_12918_, _12917_, _12892_);
  not (_12919_, _08260_);
  and (_12920_, _07939_, \oc8051_golden_model_1.P0 [3]);
  and (_12921_, _08600_, \oc8051_golden_model_1.TCON [3]);
  and (_12922_, _08603_, \oc8051_golden_model_1.P1 [3]);
  and (_12923_, _08612_, \oc8051_golden_model_1.SCON [3]);
  and (_12924_, _08614_, \oc8051_golden_model_1.P2 [3]);
  and (_12925_, _08609_, \oc8051_golden_model_1.IE [3]);
  and (_12926_, _08607_, \oc8051_golden_model_1.P3 [3]);
  and (_12927_, _08589_, \oc8051_golden_model_1.IP [3]);
  and (_12928_, _08592_, \oc8051_golden_model_1.PSW [3]);
  and (_12929_, _08596_, \oc8051_golden_model_1.ACC [3]);
  and (_12930_, _08594_, \oc8051_golden_model_1.B [3]);
  or (_12931_, _12930_, _12929_);
  or (_12932_, _12931_, _12928_);
  or (_12933_, _12932_, _12927_);
  or (_12934_, _12933_, _12926_);
  or (_12935_, _12934_, _12925_);
  or (_12936_, _12935_, _12924_);
  or (_12937_, _12936_, _12923_);
  or (_12938_, _12937_, _12922_);
  or (_12939_, _12938_, _12921_);
  nor (_12940_, _12939_, _12920_);
  and (_12941_, _12940_, _08278_);
  nor (_12942_, _12941_, _12919_);
  and (_12943_, _08589_, \oc8051_golden_model_1.IP [5]);
  and (_12944_, _08592_, \oc8051_golden_model_1.PSW [5]);
  and (_12945_, _08596_, \oc8051_golden_model_1.ACC [5]);
  and (_12946_, _08594_, \oc8051_golden_model_1.B [5]);
  or (_12947_, _12946_, _12945_);
  or (_12948_, _12947_, _12944_);
  and (_12949_, _08600_, \oc8051_golden_model_1.TCON [5]);
  and (_12950_, _07939_, \oc8051_golden_model_1.P0 [5]);
  and (_12951_, _08603_, \oc8051_golden_model_1.P1 [5]);
  or (_12952_, _12951_, _12950_);
  or (_12953_, _12952_, _12949_);
  and (_12954_, _08607_, \oc8051_golden_model_1.P3 [5]);
  and (_12955_, _08609_, \oc8051_golden_model_1.IE [5]);
  or (_12956_, _12955_, _12954_);
  and (_12957_, _08612_, \oc8051_golden_model_1.SCON [5]);
  and (_12958_, _08614_, \oc8051_golden_model_1.P2 [5]);
  or (_12959_, _12958_, _12957_);
  or (_12960_, _12959_, _12956_);
  or (_12961_, _12960_, _12953_);
  or (_12962_, _12961_, _12948_);
  nor (_12963_, _12962_, _12943_);
  and (_12964_, _12963_, _08229_);
  and (_12965_, _07892_, _06647_);
  not (_12966_, _12965_);
  nor (_12967_, _12966_, _12964_);
  nor (_12968_, _12967_, _12942_);
  and (_12969_, _12968_, _12918_);
  and (_12970_, _12969_, _12866_);
  nand (_12971_, _12368_, _12970_);
  or (_12972_, _09465_, _12970_);
  and (_12973_, _12972_, _06436_);
  and (_12974_, _12973_, _12971_);
  or (_12975_, _12974_, _12790_);
  or (_12976_, _12975_, _12789_);
  and (_12977_, _12976_, _12130_);
  nor (_12978_, _10474_, _06292_);
  not (_12979_, _12978_);
  or (_12980_, _12979_, _12977_);
  not (_12981_, _10472_);
  or (_12982_, _12978_, _09472_);
  and (_12983_, _12982_, _12981_);
  and (_12984_, _12983_, _12980_);
  and (_12985_, _12128_, _10472_);
  or (_12986_, _12985_, _06290_);
  or (_12987_, _12986_, _12984_);
  or (_12988_, _08536_, _06291_);
  and (_12989_, _12988_, _12987_);
  or (_12990_, _12989_, _05994_);
  nand (_12991_, _09473_, _05994_);
  and (_12992_, _12991_, _06435_);
  and (_12993_, _12992_, _12990_);
  or (_12994_, _12413_, _12970_);
  nand (_12995_, _12362_, _12970_);
  and (_12996_, _12995_, _12994_);
  and (_12997_, _12996_, _06434_);
  and (_12998_, _08547_, _07244_);
  not (_12999_, _12998_);
  or (_13000_, _12999_, _12997_);
  or (_13001_, _13000_, _12993_);
  or (_13002_, _12998_, _12128_);
  and (_13003_, _13002_, _07240_);
  and (_13004_, _13003_, _13001_);
  nor (_13005_, _11320_, _11315_);
  nand (_13006_, _09472_, _06559_);
  nand (_13007_, _13006_, _13005_);
  or (_13008_, _13007_, _13004_);
  or (_13009_, _12128_, _13005_);
  and (_13010_, _13009_, _06433_);
  and (_13011_, _13010_, _13008_);
  and (_13012_, _06432_, _06181_);
  or (_13013_, _13012_, _05991_);
  or (_13014_, _13013_, _13011_);
  nand (_13015_, _09473_, _05991_);
  and (_13016_, _13015_, _05933_);
  and (_13017_, _13016_, _13014_);
  and (_13018_, _12996_, _05932_);
  nor (_13019_, _09413_, _07261_);
  not (_13020_, _13019_);
  or (_13021_, _13020_, _13018_);
  or (_13022_, _13021_, _13017_);
  or (_13023_, _13019_, _12128_);
  and (_13024_, _13023_, _06570_);
  and (_13025_, _13024_, _13022_);
  nand (_13026_, _09472_, _06566_);
  nor (_13027_, _11345_, _11338_);
  nand (_13028_, _13027_, _13026_);
  or (_13029_, _13028_, _13025_);
  not (_13030_, _06393_);
  or (_13031_, _13027_, _12128_);
  and (_13032_, _13031_, _13030_);
  and (_13033_, _13032_, _13029_);
  nand (_13034_, _06393_, _06181_);
  and (_13035_, _05766_, _05931_);
  nor (_13036_, _13035_, _05989_);
  nand (_13037_, _13036_, _13034_);
  or (_13038_, _13037_, _13033_);
  not (_13039_, _13035_);
  or (_13040_, _13039_, _12128_);
  nand (_13041_, _09473_, _05989_);
  and (_13042_, _13041_, _01320_);
  and (_13043_, _13042_, _13040_);
  and (_13044_, _13043_, _13038_);
  or (_13045_, _13044_, _12115_);
  and (_40325_, _13045_, _42355_);
  not (_13046_, _07876_);
  and (_13047_, _13046_, \oc8051_golden_model_1.P2 [7]);
  and (_13048_, _08536_, _07876_);
  or (_13049_, _13048_, _13047_);
  or (_13050_, _13049_, _06260_);
  not (_13051_, _08614_);
  and (_13052_, _13051_, \oc8051_golden_model_1.P2 [7]);
  and (_13053_, _08622_, _08614_);
  or (_13054_, _13053_, _13052_);
  and (_13055_, _13054_, _06277_);
  and (_13056_, _08637_, _07876_);
  or (_13057_, _13056_, _13047_);
  or (_13058_, _13057_, _06286_);
  and (_13059_, _07876_, \oc8051_golden_model_1.ACC [7]);
  or (_13060_, _13059_, _13047_);
  and (_13061_, _13060_, _07143_);
  and (_13062_, _07144_, \oc8051_golden_model_1.P2 [7]);
  or (_13063_, _13062_, _06285_);
  or (_13064_, _13063_, _13061_);
  and (_13065_, _13064_, _06282_);
  and (_13066_, _13065_, _13058_);
  and (_13067_, _08626_, _08614_);
  or (_13068_, _13067_, _13052_);
  and (_13069_, _13068_, _06281_);
  or (_13070_, _13069_, _06354_);
  or (_13071_, _13070_, _13066_);
  or (_13072_, _13049_, _07169_);
  and (_13073_, _13072_, _13071_);
  or (_13074_, _13073_, _06345_);
  or (_13075_, _13060_, _06346_);
  and (_13076_, _13075_, _06278_);
  and (_13077_, _13076_, _13074_);
  or (_13078_, _13077_, _13055_);
  and (_13079_, _13078_, _06271_);
  or (_13080_, _13052_, _08768_);
  and (_13081_, _13080_, _06270_);
  and (_13082_, _13081_, _13068_);
  or (_13083_, _13082_, _13079_);
  and (_13084_, _13083_, _06267_);
  and (_13085_, _08789_, _08614_);
  or (_13086_, _13085_, _13052_);
  and (_13087_, _13086_, _06266_);
  or (_13088_, _13087_, _06259_);
  or (_13089_, _13088_, _13084_);
  and (_13090_, _13089_, _13050_);
  or (_13091_, _13090_, _09486_);
  and (_13092_, _08731_, _07876_);
  or (_13093_, _13047_, _06258_);
  or (_13094_, _13093_, _13092_);
  and (_13095_, _13094_, _06251_);
  and (_13096_, _13095_, _13091_);
  and (_13097_, _09004_, _07876_);
  or (_13098_, _13097_, _13047_);
  and (_13099_, _13098_, _05972_);
  or (_13100_, _13099_, _10080_);
  or (_13101_, _13100_, _13096_);
  and (_13102_, _09034_, _07876_);
  or (_13103_, _13047_, _09025_);
  or (_13104_, _13103_, _13102_);
  and (_13105_, _08806_, _07876_);
  or (_13106_, _13105_, _13047_);
  or (_13107_, _13106_, _06216_);
  and (_13108_, _13107_, _09030_);
  and (_13109_, _13108_, _13104_);
  and (_13110_, _13109_, _13101_);
  and (_13111_, _09042_, _07876_);
  or (_13112_, _13111_, _13047_);
  and (_13113_, _13112_, _06524_);
  or (_13114_, _13113_, _13110_);
  and (_13115_, _13114_, _07219_);
  or (_13116_, _13047_, _08026_);
  and (_13117_, _13106_, _06426_);
  and (_13118_, _13117_, _13116_);
  or (_13119_, _13118_, _13115_);
  and (_13120_, _13119_, _07217_);
  and (_13121_, _13060_, _06532_);
  and (_13122_, _13121_, _13116_);
  or (_13123_, _13122_, _06437_);
  or (_13124_, _13123_, _13120_);
  and (_13125_, _09033_, _07876_);
  or (_13126_, _13047_, _07229_);
  or (_13127_, _13126_, _13125_);
  and (_13128_, _13127_, _07231_);
  and (_13129_, _13128_, _13124_);
  nor (_13130_, _09041_, _13046_);
  or (_13131_, _13130_, _13047_);
  and (_13132_, _13131_, _06535_);
  or (_13133_, _13132_, _06559_);
  or (_13134_, _13133_, _13129_);
  or (_13135_, _13057_, _07240_);
  and (_13136_, _13135_, _05933_);
  and (_13137_, _13136_, _13134_);
  and (_13138_, _13054_, _05932_);
  or (_13139_, _13138_, _06566_);
  or (_13140_, _13139_, _13137_);
  and (_13141_, _08534_, _07876_);
  or (_13142_, _13047_, _06570_);
  or (_13143_, _13142_, _13141_);
  and (_13144_, _13143_, _01320_);
  and (_13145_, _13144_, _13140_);
  nor (_13146_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_13147_, _13146_, _00000_);
  or (_40326_, _13147_, _13145_);
  not (_13148_, _07885_);
  and (_13149_, _13148_, \oc8051_golden_model_1.P3 [7]);
  and (_13150_, _08536_, _07885_);
  or (_13151_, _13150_, _13149_);
  or (_13152_, _13151_, _06260_);
  not (_13153_, _08607_);
  and (_13154_, _13153_, \oc8051_golden_model_1.P3 [7]);
  and (_13155_, _08622_, _08607_);
  or (_13156_, _13155_, _13154_);
  and (_13157_, _13156_, _06277_);
  and (_13158_, _08637_, _07885_);
  or (_13159_, _13158_, _13149_);
  or (_13160_, _13159_, _06286_);
  and (_13161_, _07885_, \oc8051_golden_model_1.ACC [7]);
  or (_13162_, _13161_, _13149_);
  and (_13163_, _13162_, _07143_);
  and (_13164_, _07144_, \oc8051_golden_model_1.P3 [7]);
  or (_13165_, _13164_, _06285_);
  or (_13166_, _13165_, _13163_);
  and (_13167_, _13166_, _06282_);
  and (_13168_, _13167_, _13160_);
  and (_13169_, _08626_, _08607_);
  or (_13170_, _13169_, _13154_);
  and (_13171_, _13170_, _06281_);
  or (_13172_, _13171_, _06354_);
  or (_13173_, _13172_, _13168_);
  or (_13174_, _13151_, _07169_);
  and (_13175_, _13174_, _13173_);
  or (_13176_, _13175_, _06345_);
  or (_13177_, _13162_, _06346_);
  and (_13178_, _13177_, _06278_);
  and (_13179_, _13178_, _13176_);
  or (_13180_, _13179_, _13157_);
  and (_13181_, _13180_, _06271_);
  and (_13182_, _08769_, _08607_);
  or (_13183_, _13182_, _13154_);
  and (_13184_, _13183_, _06270_);
  or (_13185_, _13184_, _13181_);
  and (_13186_, _13185_, _06267_);
  and (_13187_, _08789_, _08607_);
  or (_13188_, _13187_, _13154_);
  and (_13189_, _13188_, _06266_);
  or (_13190_, _13189_, _06259_);
  or (_13191_, _13190_, _13186_);
  and (_13192_, _13191_, _13152_);
  or (_13193_, _13192_, _09486_);
  and (_13194_, _08731_, _07885_);
  or (_13195_, _13149_, _06258_);
  or (_13196_, _13195_, _13194_);
  and (_13197_, _13196_, _06251_);
  and (_13198_, _13197_, _13193_);
  and (_13199_, _09004_, _07885_);
  or (_13200_, _13199_, _13149_);
  and (_13201_, _13200_, _05972_);
  or (_13202_, _13201_, _10080_);
  or (_13203_, _13202_, _13198_);
  and (_13204_, _09034_, _07885_);
  or (_13205_, _13149_, _09025_);
  or (_13206_, _13205_, _13204_);
  and (_13207_, _08806_, _07885_);
  or (_13208_, _13207_, _13149_);
  or (_13209_, _13208_, _06216_);
  and (_13210_, _13209_, _09030_);
  and (_13211_, _13210_, _13206_);
  and (_13212_, _13211_, _13203_);
  and (_13213_, _09042_, _07885_);
  or (_13214_, _13213_, _13149_);
  and (_13215_, _13214_, _06524_);
  or (_13216_, _13215_, _13212_);
  and (_13217_, _13216_, _07219_);
  or (_13218_, _13149_, _08026_);
  and (_13219_, _13208_, _06426_);
  and (_13220_, _13219_, _13218_);
  or (_13221_, _13220_, _13217_);
  and (_13222_, _13221_, _07217_);
  and (_13223_, _13162_, _06532_);
  and (_13224_, _13223_, _13218_);
  or (_13225_, _13224_, _06437_);
  or (_13226_, _13225_, _13222_);
  and (_13227_, _09033_, _07885_);
  or (_13228_, _13149_, _07229_);
  or (_13229_, _13228_, _13227_);
  and (_13230_, _13229_, _07231_);
  and (_13231_, _13230_, _13226_);
  nor (_13232_, _09041_, _13148_);
  or (_13233_, _13232_, _13149_);
  and (_13234_, _13233_, _06535_);
  or (_13235_, _13234_, _06559_);
  or (_13236_, _13235_, _13231_);
  or (_13237_, _13159_, _07240_);
  and (_13238_, _13237_, _05933_);
  and (_13239_, _13238_, _13236_);
  and (_13240_, _13156_, _05932_);
  or (_13241_, _13240_, _06566_);
  or (_13242_, _13241_, _13239_);
  and (_13243_, _08534_, _07885_);
  or (_13244_, _13149_, _06570_);
  or (_13245_, _13244_, _13243_);
  and (_13246_, _13245_, _01320_);
  and (_13247_, _13246_, _13242_);
  nor (_13248_, \oc8051_golden_model_1.P3 [7], rst);
  nor (_13249_, _13248_, _00000_);
  or (_40327_, _13249_, _13247_);
  not (_13250_, _07946_);
  and (_13251_, _13250_, \oc8051_golden_model_1.P0 [7]);
  and (_13252_, _08536_, _07946_);
  or (_13253_, _13252_, _13251_);
  or (_13254_, _13253_, _06260_);
  not (_13255_, _07939_);
  and (_13256_, _13255_, \oc8051_golden_model_1.P0 [7]);
  and (_13257_, _08622_, _07939_);
  or (_13258_, _13257_, _13256_);
  and (_13259_, _13258_, _06277_);
  and (_13260_, _08637_, _07946_);
  or (_13261_, _13260_, _13251_);
  or (_13262_, _13261_, _06286_);
  and (_13263_, _07946_, \oc8051_golden_model_1.ACC [7]);
  or (_13264_, _13263_, _13251_);
  and (_13265_, _13264_, _07143_);
  and (_13266_, _07144_, \oc8051_golden_model_1.P0 [7]);
  or (_13267_, _13266_, _06285_);
  or (_13268_, _13267_, _13265_);
  and (_13269_, _13268_, _06282_);
  and (_13270_, _13269_, _13262_);
  and (_13271_, _08626_, _07939_);
  or (_13272_, _13271_, _13256_);
  and (_13273_, _13272_, _06281_);
  or (_13274_, _13273_, _06354_);
  or (_13275_, _13274_, _13270_);
  or (_13276_, _13253_, _07169_);
  and (_13277_, _13276_, _13275_);
  or (_13278_, _13277_, _06345_);
  or (_13279_, _13264_, _06346_);
  and (_13280_, _13279_, _06278_);
  and (_13281_, _13280_, _13278_);
  or (_13282_, _13281_, _13259_);
  and (_13283_, _13282_, _06271_);
  and (_13284_, _08769_, _07939_);
  or (_13285_, _13284_, _13256_);
  and (_13286_, _13285_, _06270_);
  or (_13287_, _13286_, _13283_);
  and (_13288_, _13287_, _06267_);
  and (_13289_, _08789_, _07939_);
  or (_13290_, _13289_, _13256_);
  and (_13291_, _13290_, _06266_);
  or (_13292_, _13291_, _06259_);
  or (_13293_, _13292_, _13288_);
  and (_13294_, _13293_, _13254_);
  or (_13295_, _13294_, _09486_);
  and (_13296_, _08731_, _07946_);
  or (_13297_, _13251_, _06258_);
  or (_13298_, _13297_, _13296_);
  and (_13299_, _13298_, _06251_);
  and (_13300_, _13299_, _13295_);
  and (_13301_, _09004_, _07946_);
  or (_13302_, _13301_, _13251_);
  and (_13303_, _13302_, _05972_);
  or (_13304_, _13303_, _10080_);
  or (_13305_, _13304_, _13300_);
  and (_13306_, _09034_, _07946_);
  or (_13307_, _13251_, _09025_);
  or (_13308_, _13307_, _13306_);
  and (_13309_, _08806_, _07946_);
  or (_13310_, _13309_, _13251_);
  or (_13311_, _13310_, _06216_);
  and (_13312_, _13311_, _09030_);
  and (_13313_, _13312_, _13308_);
  and (_13314_, _13313_, _13305_);
  and (_13315_, _09042_, _07946_);
  or (_13316_, _13315_, _13251_);
  and (_13317_, _13316_, _06524_);
  or (_13318_, _13317_, _13314_);
  and (_13319_, _13318_, _07219_);
  or (_13320_, _13251_, _08026_);
  and (_13321_, _13310_, _06426_);
  and (_13322_, _13321_, _13320_);
  or (_13323_, _13322_, _13319_);
  and (_13324_, _13323_, _07217_);
  and (_13325_, _13264_, _06532_);
  and (_13326_, _13325_, _13320_);
  or (_13327_, _13326_, _06437_);
  or (_13328_, _13327_, _13324_);
  and (_13329_, _09033_, _07946_);
  or (_13330_, _13251_, _07229_);
  or (_13331_, _13330_, _13329_);
  and (_13332_, _13331_, _07231_);
  and (_13333_, _13332_, _13328_);
  nor (_13334_, _09041_, _13250_);
  or (_13335_, _13334_, _13251_);
  and (_13336_, _13335_, _06535_);
  or (_13337_, _13336_, _06559_);
  or (_13338_, _13337_, _13333_);
  or (_13339_, _13261_, _07240_);
  and (_13340_, _13339_, _05933_);
  and (_13341_, _13340_, _13338_);
  and (_13342_, _13258_, _05932_);
  or (_13343_, _13342_, _06566_);
  or (_13344_, _13343_, _13341_);
  and (_13345_, _08534_, _07946_);
  or (_13346_, _13251_, _06570_);
  or (_13347_, _13346_, _13345_);
  and (_13348_, _13347_, _01320_);
  and (_13349_, _13348_, _13344_);
  nor (_13350_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_13351_, _13350_, _00000_);
  or (_40328_, _13351_, _13349_);
  nor (_13352_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_13353_, _13352_, _00000_);
  not (_13354_, _07961_);
  and (_13355_, _13354_, \oc8051_golden_model_1.P1 [7]);
  and (_13356_, _08536_, _07961_);
  or (_13357_, _13356_, _13355_);
  or (_13358_, _13357_, _06260_);
  not (_13359_, _08603_);
  and (_13360_, _13359_, \oc8051_golden_model_1.P1 [7]);
  and (_13361_, _08622_, _08603_);
  or (_13362_, _13361_, _13360_);
  and (_13363_, _13362_, _06277_);
  and (_13364_, _08637_, _07961_);
  or (_13365_, _13364_, _13355_);
  or (_13366_, _13365_, _06286_);
  and (_13367_, _07961_, \oc8051_golden_model_1.ACC [7]);
  or (_13368_, _13367_, _13355_);
  and (_13369_, _13368_, _07143_);
  and (_13370_, _07144_, \oc8051_golden_model_1.P1 [7]);
  or (_13371_, _13370_, _06285_);
  or (_13372_, _13371_, _13369_);
  and (_13373_, _13372_, _06282_);
  and (_13374_, _13373_, _13366_);
  and (_13375_, _08626_, _08603_);
  or (_13376_, _13375_, _13360_);
  and (_13377_, _13376_, _06281_);
  or (_13378_, _13377_, _06354_);
  or (_13379_, _13378_, _13374_);
  or (_13380_, _13357_, _07169_);
  and (_13381_, _13380_, _13379_);
  or (_13382_, _13381_, _06345_);
  or (_13383_, _13368_, _06346_);
  and (_13384_, _13383_, _06278_);
  and (_13385_, _13384_, _13382_);
  or (_13386_, _13385_, _13363_);
  and (_13387_, _13386_, _06271_);
  or (_13388_, _13360_, _08768_);
  and (_13389_, _13388_, _06270_);
  and (_13390_, _13389_, _13376_);
  or (_13391_, _13390_, _13387_);
  and (_13392_, _13391_, _06267_);
  and (_13393_, _08789_, _08603_);
  or (_13394_, _13393_, _13360_);
  and (_13395_, _13394_, _06266_);
  or (_13396_, _13395_, _06259_);
  or (_13397_, _13396_, _13392_);
  and (_13398_, _13397_, _13358_);
  or (_13399_, _13398_, _09486_);
  and (_13400_, _08731_, _07961_);
  or (_13401_, _13355_, _06258_);
  or (_13402_, _13401_, _13400_);
  and (_13403_, _13402_, _06251_);
  and (_13404_, _13403_, _13399_);
  and (_13405_, _09004_, _07961_);
  or (_13406_, _13405_, _13355_);
  and (_13407_, _13406_, _05972_);
  or (_13408_, _13407_, _10080_);
  or (_13409_, _13408_, _13404_);
  and (_13410_, _09034_, _07961_);
  or (_13411_, _13355_, _09025_);
  or (_13412_, _13411_, _13410_);
  and (_13413_, _08806_, _07961_);
  or (_13414_, _13413_, _13355_);
  or (_13415_, _13414_, _06216_);
  and (_13416_, _13415_, _09030_);
  and (_13417_, _13416_, _13412_);
  and (_13418_, _13417_, _13409_);
  and (_13419_, _09042_, _07961_);
  or (_13420_, _13419_, _13355_);
  and (_13421_, _13420_, _06524_);
  or (_13422_, _13421_, _13418_);
  and (_13423_, _13422_, _07219_);
  or (_13424_, _13355_, _08026_);
  and (_13425_, _13414_, _06426_);
  and (_13426_, _13425_, _13424_);
  or (_13427_, _13426_, _13423_);
  and (_13428_, _13427_, _07217_);
  and (_13429_, _13368_, _06532_);
  and (_13430_, _13429_, _13424_);
  or (_13431_, _13430_, _06437_);
  or (_13432_, _13431_, _13428_);
  and (_13433_, _09033_, _07961_);
  or (_13434_, _13355_, _07229_);
  or (_13435_, _13434_, _13433_);
  and (_13436_, _13435_, _07231_);
  and (_13437_, _13436_, _13432_);
  nor (_13438_, _09041_, _13354_);
  or (_13439_, _13438_, _13355_);
  and (_13440_, _13439_, _06535_);
  or (_13441_, _13440_, _06559_);
  or (_13442_, _13441_, _13437_);
  or (_13443_, _13365_, _07240_);
  and (_13444_, _13443_, _05933_);
  and (_13445_, _13444_, _13442_);
  and (_13446_, _13362_, _05932_);
  or (_13447_, _13446_, _06566_);
  or (_13448_, _13447_, _13445_);
  and (_13449_, _08534_, _07961_);
  or (_13450_, _13355_, _06570_);
  or (_13451_, _13450_, _13449_);
  and (_13452_, _13451_, _01320_);
  and (_13453_, _13452_, _13448_);
  or (_40330_, _13453_, _13353_);
  and (_13454_, _01324_, \oc8051_golden_model_1.IP [7]);
  not (_13455_, _07937_);
  and (_13456_, _13455_, \oc8051_golden_model_1.IP [7]);
  and (_13457_, _08536_, _07937_);
  or (_13458_, _13457_, _13456_);
  or (_13459_, _13458_, _06260_);
  not (_13460_, _08589_);
  and (_13461_, _13460_, \oc8051_golden_model_1.IP [7]);
  and (_13462_, _08622_, _08589_);
  or (_13463_, _13462_, _13461_);
  and (_13464_, _13463_, _06277_);
  and (_13465_, _08637_, _07937_);
  or (_13466_, _13465_, _13456_);
  or (_13467_, _13466_, _06286_);
  and (_13468_, _07937_, \oc8051_golden_model_1.ACC [7]);
  or (_13469_, _13468_, _13456_);
  and (_13470_, _13469_, _07143_);
  and (_13471_, _07144_, \oc8051_golden_model_1.IP [7]);
  or (_13472_, _13471_, _06285_);
  or (_13473_, _13472_, _13470_);
  and (_13474_, _13473_, _06282_);
  and (_13475_, _13474_, _13467_);
  and (_13476_, _08626_, _08589_);
  or (_13477_, _13476_, _13461_);
  and (_13478_, _13477_, _06281_);
  or (_13479_, _13478_, _06354_);
  or (_13480_, _13479_, _13475_);
  or (_13481_, _13458_, _07169_);
  and (_13482_, _13481_, _13480_);
  or (_13483_, _13482_, _06345_);
  or (_13484_, _13469_, _06346_);
  and (_13485_, _13484_, _06278_);
  and (_13486_, _13485_, _13483_);
  or (_13487_, _13486_, _13464_);
  and (_13488_, _13487_, _06271_);
  and (_13489_, _08769_, _08589_);
  or (_13490_, _13489_, _13461_);
  and (_13491_, _13490_, _06270_);
  or (_13492_, _13491_, _13488_);
  and (_13493_, _13492_, _06267_);
  and (_13494_, _08789_, _08589_);
  or (_13495_, _13494_, _13461_);
  and (_13496_, _13495_, _06266_);
  or (_13497_, _13496_, _06259_);
  or (_13498_, _13497_, _13493_);
  and (_13499_, _13498_, _13459_);
  or (_13500_, _13499_, _09486_);
  and (_13501_, _08731_, _07937_);
  or (_13502_, _13456_, _06258_);
  or (_13503_, _13502_, _13501_);
  and (_13504_, _13503_, _06251_);
  and (_13505_, _13504_, _13500_);
  and (_13506_, _09004_, _07937_);
  or (_13507_, _13506_, _13456_);
  and (_13508_, _13507_, _05972_);
  or (_13509_, _13508_, _10080_);
  or (_13510_, _13509_, _13505_);
  and (_13511_, _09034_, _07937_);
  or (_13512_, _13456_, _09025_);
  or (_13513_, _13512_, _13511_);
  and (_13514_, _08806_, _07937_);
  or (_13515_, _13514_, _13456_);
  or (_13516_, _13515_, _06216_);
  and (_13517_, _13516_, _09030_);
  and (_13518_, _13517_, _13513_);
  and (_13519_, _13518_, _13510_);
  and (_13520_, _09042_, _07937_);
  or (_13521_, _13520_, _13456_);
  and (_13522_, _13521_, _06524_);
  or (_13523_, _13522_, _13519_);
  and (_13524_, _13523_, _07219_);
  or (_13525_, _13456_, _08026_);
  and (_13526_, _13515_, _06426_);
  and (_13527_, _13526_, _13525_);
  or (_13528_, _13527_, _13524_);
  and (_13529_, _13528_, _07217_);
  and (_13530_, _13469_, _06532_);
  and (_13531_, _13530_, _13525_);
  or (_13532_, _13531_, _06437_);
  or (_13533_, _13532_, _13529_);
  and (_13534_, _09033_, _07937_);
  or (_13535_, _13456_, _07229_);
  or (_13536_, _13535_, _13534_);
  and (_13537_, _13536_, _07231_);
  and (_13538_, _13537_, _13533_);
  nor (_13539_, _09041_, _13455_);
  or (_13540_, _13539_, _13456_);
  and (_13541_, _13540_, _06535_);
  or (_13542_, _13541_, _06559_);
  or (_13543_, _13542_, _13538_);
  or (_13544_, _13466_, _07240_);
  and (_13545_, _13544_, _05933_);
  and (_13546_, _13545_, _13543_);
  and (_13547_, _13463_, _05932_);
  or (_13548_, _13547_, _06566_);
  or (_13549_, _13548_, _13546_);
  and (_13550_, _08534_, _07937_);
  or (_13551_, _13456_, _06570_);
  or (_13552_, _13551_, _13550_);
  and (_13553_, _13552_, _01320_);
  and (_13554_, _13553_, _13549_);
  or (_13555_, _13554_, _13454_);
  and (_40331_, _13555_, _42355_);
  and (_13556_, _01324_, \oc8051_golden_model_1.IE [7]);
  not (_13557_, _07881_);
  and (_13558_, _13557_, \oc8051_golden_model_1.IE [7]);
  and (_13559_, _08536_, _07881_);
  or (_13560_, _13559_, _13558_);
  or (_13561_, _13560_, _06260_);
  not (_13562_, _08609_);
  and (_13563_, _13562_, \oc8051_golden_model_1.IE [7]);
  and (_13564_, _08622_, _08609_);
  or (_13565_, _13564_, _13563_);
  and (_13566_, _13565_, _06277_);
  and (_13567_, _08637_, _07881_);
  or (_13568_, _13567_, _13558_);
  or (_13569_, _13568_, _06286_);
  and (_13570_, _07881_, \oc8051_golden_model_1.ACC [7]);
  or (_13571_, _13570_, _13558_);
  and (_13572_, _13571_, _07143_);
  and (_13573_, _07144_, \oc8051_golden_model_1.IE [7]);
  or (_13574_, _13573_, _06285_);
  or (_13575_, _13574_, _13572_);
  and (_13576_, _13575_, _06282_);
  and (_13577_, _13576_, _13569_);
  and (_13578_, _08626_, _08609_);
  or (_13579_, _13578_, _13563_);
  and (_13580_, _13579_, _06281_);
  or (_13581_, _13580_, _06354_);
  or (_13582_, _13581_, _13577_);
  or (_13583_, _13560_, _07169_);
  and (_13584_, _13583_, _13582_);
  or (_13585_, _13584_, _06345_);
  or (_13586_, _13571_, _06346_);
  and (_13587_, _13586_, _06278_);
  and (_13588_, _13587_, _13585_);
  or (_13589_, _13588_, _13566_);
  and (_13590_, _13589_, _06271_);
  and (_13591_, _08769_, _08609_);
  or (_13592_, _13591_, _13563_);
  and (_13593_, _13592_, _06270_);
  or (_13594_, _13593_, _13590_);
  and (_13595_, _13594_, _06267_);
  and (_13596_, _08789_, _08609_);
  or (_13597_, _13596_, _13563_);
  and (_13598_, _13597_, _06266_);
  or (_13599_, _13598_, _06259_);
  or (_13600_, _13599_, _13595_);
  and (_13601_, _13600_, _13561_);
  or (_13602_, _13601_, _09486_);
  and (_13603_, _08731_, _07881_);
  or (_13604_, _13558_, _06258_);
  or (_13605_, _13604_, _13603_);
  and (_13606_, _13605_, _06251_);
  and (_13607_, _13606_, _13602_);
  and (_13608_, _09004_, _07881_);
  or (_13609_, _13608_, _13558_);
  and (_13610_, _13609_, _05972_);
  or (_13611_, _13610_, _10080_);
  or (_13612_, _13611_, _13607_);
  and (_13613_, _09034_, _07881_);
  or (_13614_, _13558_, _09025_);
  or (_13615_, _13614_, _13613_);
  and (_13616_, _08806_, _07881_);
  or (_13617_, _13616_, _13558_);
  or (_13619_, _13617_, _06216_);
  and (_13620_, _13619_, _09030_);
  and (_13621_, _13620_, _13615_);
  and (_13622_, _13621_, _13612_);
  and (_13623_, _09042_, _07881_);
  or (_13624_, _13623_, _13558_);
  and (_13625_, _13624_, _06524_);
  or (_13626_, _13625_, _13622_);
  and (_13627_, _13626_, _07219_);
  or (_13628_, _13558_, _08026_);
  and (_13630_, _13617_, _06426_);
  and (_13631_, _13630_, _13628_);
  or (_13632_, _13631_, _13627_);
  and (_13633_, _13632_, _07217_);
  and (_13634_, _13571_, _06532_);
  and (_13635_, _13634_, _13628_);
  or (_13636_, _13635_, _06437_);
  or (_13637_, _13636_, _13633_);
  and (_13638_, _09033_, _07881_);
  or (_13639_, _13558_, _07229_);
  or (_13641_, _13639_, _13638_);
  and (_13642_, _13641_, _07231_);
  and (_13643_, _13642_, _13637_);
  nor (_13644_, _09041_, _13557_);
  or (_13645_, _13644_, _13558_);
  and (_13646_, _13645_, _06535_);
  or (_13647_, _13646_, _06559_);
  or (_13648_, _13647_, _13643_);
  or (_13649_, _13568_, _07240_);
  and (_13650_, _13649_, _05933_);
  and (_13652_, _13650_, _13648_);
  and (_13653_, _13565_, _05932_);
  or (_13654_, _13653_, _06566_);
  or (_13655_, _13654_, _13652_);
  and (_13656_, _08534_, _07881_);
  or (_13657_, _13558_, _06570_);
  or (_13658_, _13657_, _13656_);
  and (_13659_, _13658_, _01320_);
  and (_13660_, _13659_, _13655_);
  or (_13661_, _13660_, _13556_);
  and (_40332_, _13661_, _42355_);
  and (_13663_, _01324_, \oc8051_golden_model_1.SCON [7]);
  not (_13664_, _07963_);
  and (_13665_, _13664_, \oc8051_golden_model_1.SCON [7]);
  and (_13666_, _08536_, _07963_);
  or (_13667_, _13666_, _13665_);
  or (_13668_, _13667_, _06260_);
  not (_13669_, _08612_);
  and (_13670_, _13669_, \oc8051_golden_model_1.SCON [7]);
  and (_13671_, _08622_, _08612_);
  or (_13673_, _13671_, _13670_);
  and (_13674_, _13673_, _06277_);
  and (_13675_, _08637_, _07963_);
  or (_13676_, _13675_, _13665_);
  or (_13677_, _13676_, _06286_);
  and (_13678_, _07963_, \oc8051_golden_model_1.ACC [7]);
  or (_13679_, _13678_, _13665_);
  and (_13680_, _13679_, _07143_);
  and (_13681_, _07144_, \oc8051_golden_model_1.SCON [7]);
  or (_13682_, _13681_, _06285_);
  or (_13684_, _13682_, _13680_);
  and (_13685_, _13684_, _06282_);
  and (_13686_, _13685_, _13677_);
  and (_13687_, _08626_, _08612_);
  or (_13688_, _13687_, _13670_);
  and (_13689_, _13688_, _06281_);
  or (_13690_, _13689_, _06354_);
  or (_13691_, _13690_, _13686_);
  or (_13692_, _13667_, _07169_);
  and (_13693_, _13692_, _13691_);
  or (_13695_, _13693_, _06345_);
  or (_13696_, _13679_, _06346_);
  and (_13697_, _13696_, _06278_);
  and (_13698_, _13697_, _13695_);
  or (_13699_, _13698_, _13674_);
  and (_13700_, _13699_, _06271_);
  and (_13701_, _08769_, _08612_);
  or (_13702_, _13701_, _13670_);
  and (_13703_, _13702_, _06270_);
  or (_13704_, _13703_, _13700_);
  and (_13706_, _13704_, _06267_);
  and (_13707_, _08789_, _08612_);
  or (_13708_, _13707_, _13670_);
  and (_13709_, _13708_, _06266_);
  or (_13710_, _13709_, _06259_);
  or (_13711_, _13710_, _13706_);
  and (_13712_, _13711_, _13668_);
  or (_13713_, _13712_, _09486_);
  and (_13714_, _08731_, _07963_);
  or (_13715_, _13665_, _06258_);
  or (_13717_, _13715_, _13714_);
  and (_13718_, _13717_, _06251_);
  and (_13719_, _13718_, _13713_);
  and (_13720_, _09004_, _07963_);
  or (_13721_, _13720_, _13665_);
  and (_13722_, _13721_, _05972_);
  or (_13723_, _13722_, _10080_);
  or (_13724_, _13723_, _13719_);
  and (_13725_, _09034_, _07963_);
  or (_13726_, _13665_, _09025_);
  or (_13728_, _13726_, _13725_);
  and (_13729_, _08806_, _07963_);
  or (_13730_, _13729_, _13665_);
  or (_13731_, _13730_, _06216_);
  and (_13732_, _13731_, _09030_);
  and (_13733_, _13732_, _13728_);
  and (_13734_, _13733_, _13724_);
  and (_13735_, _09042_, _07963_);
  or (_13736_, _13735_, _13665_);
  and (_13737_, _13736_, _06524_);
  or (_13739_, _13737_, _13734_);
  and (_13740_, _13739_, _07219_);
  or (_13741_, _13665_, _08026_);
  and (_13742_, _13730_, _06426_);
  and (_13743_, _13742_, _13741_);
  or (_13744_, _13743_, _13740_);
  and (_13745_, _13744_, _07217_);
  and (_13746_, _13679_, _06532_);
  and (_13747_, _13746_, _13741_);
  or (_13748_, _13747_, _06437_);
  or (_13750_, _13748_, _13745_);
  and (_13751_, _09033_, _07963_);
  or (_13752_, _13665_, _07229_);
  or (_13753_, _13752_, _13751_);
  and (_13754_, _13753_, _07231_);
  and (_13755_, _13754_, _13750_);
  nor (_13756_, _09041_, _13664_);
  or (_13757_, _13756_, _13665_);
  and (_13758_, _13757_, _06535_);
  or (_13759_, _13758_, _06559_);
  or (_13761_, _13759_, _13755_);
  or (_13762_, _13676_, _07240_);
  and (_13763_, _13762_, _05933_);
  and (_13764_, _13763_, _13761_);
  and (_13765_, _13673_, _05932_);
  or (_13766_, _13765_, _06566_);
  or (_13767_, _13766_, _13764_);
  and (_13768_, _08534_, _07963_);
  or (_13769_, _13665_, _06570_);
  or (_13770_, _13769_, _13768_);
  and (_13771_, _13770_, _01320_);
  and (_13772_, _13771_, _13767_);
  or (_13773_, _13772_, _13663_);
  and (_40333_, _13773_, _42355_);
  not (_13774_, \oc8051_golden_model_1.SP [7]);
  nor (_13775_, _01320_, _13774_);
  and (_13776_, _07585_, \oc8051_golden_model_1.SP [4]);
  and (_13777_, _13776_, \oc8051_golden_model_1.SP [5]);
  and (_13778_, _13777_, \oc8051_golden_model_1.SP [6]);
  or (_13779_, _13778_, \oc8051_golden_model_1.SP [7]);
  nand (_13780_, _13778_, \oc8051_golden_model_1.SP [7]);
  and (_13781_, _13780_, _13779_);
  or (_13782_, _13781_, _07252_);
  nor (_13783_, _07919_, _13774_);
  and (_13784_, _09042_, _08256_);
  or (_13785_, _13784_, _13783_);
  and (_13786_, _13785_, _06524_);
  not (_13787_, _06261_);
  and (_13788_, _08536_, _08256_);
  or (_13789_, _13783_, _09486_);
  or (_13790_, _13789_, _13788_);
  and (_13791_, _13790_, _13787_);
  and (_13792_, _08637_, _08256_);
  or (_13793_, _13792_, _13783_);
  or (_13794_, _13793_, _06286_);
  and (_13795_, _07919_, \oc8051_golden_model_1.ACC [7]);
  or (_13796_, _13795_, _13783_);
  or (_13797_, _13796_, _07144_);
  or (_13798_, _07143_, \oc8051_golden_model_1.SP [7]);
  and (_13799_, _13798_, _07858_);
  and (_13800_, _13799_, _13797_);
  and (_13801_, _13781_, _07152_);
  or (_13802_, _13801_, _06285_);
  or (_13803_, _13802_, _13800_);
  and (_13804_, _13803_, _05949_);
  and (_13805_, _13804_, _13794_);
  and (_13806_, _13781_, _07460_);
  or (_13807_, _13806_, _06354_);
  or (_13808_, _13807_, _13805_);
  not (_13809_, \oc8051_golden_model_1.SP [6]);
  not (_13810_, \oc8051_golden_model_1.SP [5]);
  not (_13811_, \oc8051_golden_model_1.SP [4]);
  and (_13812_, _08645_, _13811_);
  and (_13813_, _13812_, _13810_);
  and (_13814_, _13813_, _13809_);
  and (_13815_, _13814_, _06766_);
  nor (_13816_, _13815_, _13774_);
  and (_13817_, _13815_, _13774_);
  nor (_13818_, _13817_, _13816_);
  nand (_13819_, _13818_, _06354_);
  and (_13820_, _13819_, _13808_);
  or (_13821_, _13820_, _06345_);
  or (_13822_, _13796_, _06346_);
  and (_13823_, _13822_, _06778_);
  and (_13824_, _13823_, _13821_);
  and (_13825_, _13777_, \oc8051_golden_model_1.SP [0]);
  and (_13826_, _13825_, \oc8051_golden_model_1.SP [6]);
  or (_13827_, _13826_, \oc8051_golden_model_1.SP [7]);
  nand (_13828_, _13826_, \oc8051_golden_model_1.SP [7]);
  and (_13829_, _13828_, _13827_);
  nand (_13830_, _13829_, _06276_);
  nand (_13831_, _13830_, _07459_);
  or (_13832_, _13831_, _13824_);
  or (_13833_, _13781_, _07459_);
  and (_13834_, _13833_, _06260_);
  and (_13835_, _13834_, _13832_);
  or (_13836_, _13835_, _13791_);
  or (_13837_, _13783_, _06258_);
  and (_13838_, _08731_, _07919_);
  or (_13839_, _13838_, _13837_);
  and (_13840_, _13839_, _06251_);
  and (_13841_, _13840_, _13836_);
  and (_13842_, _09004_, _08256_);
  or (_13843_, _13842_, _13783_);
  and (_13844_, _13843_, _05972_);
  or (_13845_, _13844_, _06215_);
  or (_13846_, _13845_, _13841_);
  and (_13847_, _08806_, _07919_);
  or (_13848_, _13847_, _13783_);
  or (_13849_, _13848_, _06216_);
  and (_13850_, _13849_, _13846_);
  or (_13851_, _13850_, _06004_);
  not (_13852_, _06004_);
  or (_13853_, _13781_, _13852_);
  and (_13854_, _13853_, _13851_);
  or (_13855_, _13854_, _06398_);
  and (_13856_, _09034_, _07919_);
  or (_13857_, _13856_, _13783_);
  or (_13858_, _13857_, _09025_);
  and (_13859_, _13858_, _09030_);
  and (_13860_, _13859_, _13855_);
  or (_13861_, _13860_, _13786_);
  and (_13862_, _13861_, _07219_);
  or (_13863_, _13783_, _08026_);
  and (_13864_, _13848_, _06426_);
  and (_13865_, _13864_, _13863_);
  or (_13866_, _13865_, _13862_);
  and (_13867_, _13866_, _12729_);
  and (_13868_, _13796_, _06532_);
  and (_13869_, _13868_, _13863_);
  and (_13870_, _13781_, _06013_);
  or (_13871_, _13870_, _06437_);
  or (_13872_, _13871_, _13869_);
  or (_13873_, _13872_, _13867_);
  and (_13874_, _09033_, _07919_);
  or (_13875_, _13874_, _13783_);
  or (_13876_, _13875_, _07229_);
  and (_13877_, _13876_, _13873_);
  or (_13878_, _13877_, _06535_);
  not (_13879_, _08256_);
  nor (_13880_, _09041_, _13879_);
  or (_13881_, _13783_, _07231_);
  or (_13882_, _13881_, _13880_);
  and (_13883_, _13882_, _12782_);
  and (_13884_, _13883_, _13878_);
  or (_13885_, _13814_, \oc8051_golden_model_1.SP [7]);
  nand (_13886_, _13814_, \oc8051_golden_model_1.SP [7]);
  and (_13887_, _13886_, _13885_);
  and (_13888_, _13887_, _06543_);
  or (_13889_, _13888_, _06011_);
  or (_13890_, _13889_, _13884_);
  or (_13891_, _13781_, _09057_);
  and (_13892_, _13891_, _13890_);
  or (_13893_, _13892_, _06290_);
  or (_13894_, _13887_, _06291_);
  and (_13895_, _13894_, _07240_);
  and (_13896_, _13895_, _13893_);
  and (_13897_, _13793_, _06559_);
  or (_13898_, _13897_, _07678_);
  or (_13899_, _13898_, _13896_);
  and (_13900_, _13899_, _13782_);
  or (_13901_, _13900_, _06566_);
  and (_13902_, _08534_, _08256_);
  or (_13903_, _13783_, _06570_);
  or (_13904_, _13903_, _13902_);
  and (_13905_, _13904_, _01320_);
  and (_13906_, _13905_, _13901_);
  or (_13907_, _13906_, _13775_);
  and (_40334_, _13907_, _42355_);
  not (_13908_, _07894_);
  and (_13909_, _13908_, \oc8051_golden_model_1.SBUF [7]);
  and (_13910_, _08536_, _07894_);
  or (_13911_, _13910_, _13909_);
  or (_13912_, _13911_, _06260_);
  and (_13913_, _08637_, _07894_);
  or (_13914_, _13913_, _13909_);
  or (_13915_, _13914_, _06286_);
  and (_13916_, _07894_, \oc8051_golden_model_1.ACC [7]);
  or (_13917_, _13916_, _13909_);
  and (_13918_, _13917_, _07143_);
  and (_13919_, _07144_, \oc8051_golden_model_1.SBUF [7]);
  or (_13920_, _13919_, _06285_);
  or (_13921_, _13920_, _13918_);
  and (_13922_, _13921_, _07169_);
  and (_13923_, _13922_, _13915_);
  and (_13924_, _13911_, _06354_);
  or (_13925_, _13924_, _13923_);
  and (_13926_, _13925_, _06346_);
  and (_13927_, _13917_, _06345_);
  or (_13928_, _13927_, _06259_);
  or (_13929_, _13928_, _13926_);
  and (_13930_, _13929_, _13912_);
  or (_13931_, _13930_, _09486_);
  and (_13932_, _08731_, _07894_);
  or (_13933_, _13909_, _06258_);
  or (_13934_, _13933_, _13932_);
  and (_13935_, _13934_, _06251_);
  and (_13936_, _13935_, _13931_);
  and (_13937_, _09004_, _07894_);
  or (_13938_, _13937_, _13909_);
  and (_13939_, _13938_, _05972_);
  or (_13940_, _13939_, _13936_);
  or (_13941_, _13940_, _10080_);
  and (_13942_, _09034_, _07894_);
  or (_13943_, _13909_, _09025_);
  or (_13944_, _13943_, _13942_);
  and (_13945_, _08806_, _07894_);
  or (_13946_, _13945_, _13909_);
  or (_13947_, _13946_, _06216_);
  and (_13948_, _13947_, _09030_);
  and (_13949_, _13948_, _13944_);
  and (_13950_, _13949_, _13941_);
  and (_13951_, _09042_, _07894_);
  or (_13952_, _13951_, _13909_);
  and (_13953_, _13952_, _06524_);
  or (_13954_, _13953_, _13950_);
  and (_13955_, _13954_, _07219_);
  or (_13956_, _13909_, _08026_);
  and (_13957_, _13946_, _06426_);
  and (_13958_, _13957_, _13956_);
  or (_13959_, _13958_, _13955_);
  and (_13960_, _13959_, _07217_);
  and (_13961_, _13917_, _06532_);
  and (_13962_, _13961_, _13956_);
  or (_13963_, _13962_, _06437_);
  or (_13964_, _13963_, _13960_);
  and (_13965_, _09033_, _07894_);
  or (_13966_, _13909_, _07229_);
  or (_13967_, _13966_, _13965_);
  and (_13968_, _13967_, _07231_);
  and (_13969_, _13968_, _13964_);
  nor (_13970_, _09041_, _13908_);
  or (_13971_, _13970_, _13909_);
  and (_13972_, _13971_, _06535_);
  or (_13973_, _13972_, _06559_);
  or (_13974_, _13973_, _13969_);
  or (_13975_, _13914_, _07240_);
  and (_13976_, _13975_, _06570_);
  and (_13977_, _13976_, _13974_);
  and (_13978_, _08534_, _07894_);
  or (_13979_, _13978_, _13909_);
  and (_13980_, _13979_, _06566_);
  or (_13981_, _13980_, _01324_);
  or (_13982_, _13981_, _13977_);
  or (_13983_, _01320_, \oc8051_golden_model_1.SBUF [7]);
  and (_13984_, _13983_, _42355_);
  and (_40336_, _13984_, _13982_);
  nor (_13985_, _01320_, _10774_);
  nor (_13986_, _08592_, _10774_);
  and (_13987_, _08622_, _08592_);
  or (_13988_, _13987_, _13986_);
  or (_13989_, _13988_, _05933_);
  not (_13990_, _11027_);
  nor (_13991_, _10732_, _08737_);
  or (_13992_, _13991_, _11049_);
  or (_13993_, _11023_, _10729_);
  or (_13994_, _13993_, _13992_);
  nor (_13995_, _07926_, _10774_);
  and (_13996_, _09042_, _07926_);
  or (_13997_, _13996_, _13995_);
  and (_13998_, _13997_, _06524_);
  and (_13999_, _09004_, _07926_);
  or (_14000_, _13999_, _13995_);
  and (_14001_, _14000_, _05972_);
  and (_14002_, _08536_, _07926_);
  or (_14003_, _14002_, _13995_);
  or (_14004_, _14003_, _06260_);
  and (_14005_, _10572_, _10568_);
  nor (_14006_, _14005_, _10566_);
  nand (_14007_, _10614_, _10568_);
  or (_14008_, _14007_, _10612_);
  and (_14009_, _14008_, _14006_);
  and (_14010_, _10562_, _08731_);
  or (_14011_, _14010_, _10555_);
  or (_14012_, _14011_, _14009_);
  not (_14013_, _06370_);
  not (_14014_, _06371_);
  nor (_14015_, _12970_, _14014_);
  nor (_14016_, _09520_, _06371_);
  and (_14017_, _12489_, _12490_);
  or (_14018_, _14017_, _12487_);
  or (_14019_, _12499_, _12497_);
  and (_14020_, _14019_, _12493_);
  or (_14021_, _14020_, _14018_);
  and (_14022_, _14021_, _12517_);
  and (_14023_, _12512_, _12513_);
  or (_14024_, _14023_, _12510_);
  and (_14025_, _14024_, _12509_);
  and (_14026_, _12507_, _12505_);
  or (_14027_, _14026_, _12504_);
  or (_14028_, _14027_, _14025_);
  or (_14029_, _14028_, _14022_);
  nor (_14030_, _12519_, _12484_);
  and (_14031_, _14030_, _14029_);
  and (_14032_, _13988_, _06277_);
  and (_14033_, _08637_, _07926_);
  or (_14034_, _14033_, _13995_);
  or (_14035_, _14034_, _06286_);
  and (_14036_, _07926_, \oc8051_golden_model_1.ACC [7]);
  or (_14037_, _14036_, _13995_);
  and (_14038_, _14037_, _07143_);
  nor (_14039_, _07143_, _10774_);
  or (_14040_, _14039_, _06285_);
  or (_14041_, _14040_, _14038_);
  and (_14042_, _14041_, _10657_);
  and (_14043_, _14042_, _14035_);
  nor (_14044_, _10678_, _10657_);
  not (_14045_, _12408_);
  nand (_14046_, _14045_, _06361_);
  or (_14047_, _14046_, _14044_);
  or (_14048_, _14047_, _14043_);
  and (_14049_, _08626_, _08592_);
  or (_14050_, _14049_, _13986_);
  or (_14051_, _14050_, _06282_);
  or (_14052_, _14003_, _07169_);
  and (_14053_, _14052_, _14051_);
  and (_14054_, _14053_, _14048_);
  or (_14055_, _14054_, _06345_);
  or (_14056_, _14037_, _06346_);
  nor (_14057_, _12467_, _06277_);
  and (_14058_, _14057_, _14056_);
  and (_14059_, _14058_, _14055_);
  or (_14060_, _14059_, _14032_);
  and (_14061_, _14060_, _12484_);
  or (_14062_, _14061_, _14031_);
  and (_14063_, _14062_, _06424_);
  nand (_14064_, _12373_, _12370_);
  nand (_14065_, _14064_, _12369_);
  or (_14066_, _12380_, _12377_);
  and (_14067_, _14066_, _12375_);
  or (_14068_, _14067_, _14065_);
  and (_14069_, _14068_, _12396_);
  nor (_14070_, _12385_, _08781_);
  or (_14071_, _14070_, _12383_);
  nand (_14072_, _12393_, _12390_);
  and (_14073_, _12388_, _14072_);
  and (_14074_, _14073_, _12389_);
  or (_14075_, _14074_, _14071_);
  or (_14076_, _14075_, _14069_);
  and (_14077_, _12398_, _06423_);
  and (_14078_, _14077_, _14076_);
  or (_14079_, _14078_, _14063_);
  and (_14080_, _14079_, _06420_);
  nand (_14081_, _08230_, \oc8051_golden_model_1.ACC [5]);
  nor (_14082_, _08230_, \oc8051_golden_model_1.ACC [5]);
  nor (_14083_, _08527_, \oc8051_golden_model_1.ACC [4]);
  or (_14084_, _14083_, _14082_);
  and (_14085_, _14084_, _14081_);
  and (_14086_, _14085_, _12538_);
  nor (_14087_, _08025_, \oc8051_golden_model_1.ACC [7]);
  or (_14088_, _08127_, \oc8051_golden_model_1.ACC [6]);
  nor (_14089_, _14088_, _09042_);
  or (_14090_, _14089_, _14087_);
  or (_14091_, _14090_, _14086_);
  nand (_14092_, _08279_, \oc8051_golden_model_1.ACC [3]);
  nor (_14093_, _08279_, \oc8051_golden_model_1.ACC [3]);
  nor (_14094_, _08423_, \oc8051_golden_model_1.ACC [2]);
  or (_14095_, _14094_, _14093_);
  and (_14096_, _14095_, _14092_);
  nor (_14097_, _08324_, \oc8051_golden_model_1.ACC [1]);
  nor (_14098_, _08374_, _06018_);
  nor (_14099_, _14098_, _11253_);
  or (_14100_, _14099_, _14097_);
  and (_14101_, _14100_, _12530_);
  or (_14102_, _14101_, _14096_);
  and (_14103_, _14102_, _12539_);
  or (_14104_, _14103_, _14091_);
  not (_14105_, _06347_);
  nor (_14106_, _12540_, _14105_);
  and (_14107_, _14106_, _14104_);
  nor (_14108_, _06995_, \oc8051_golden_model_1.ACC [1]);
  and (_14109_, _06995_, \oc8051_golden_model_1.ACC [1]);
  nor (_14110_, _06248_, _06018_);
  nor (_14111_, _14110_, _14109_);
  or (_14112_, _14111_, _14108_);
  and (_14113_, _14112_, _12550_);
  and (_14114_, _12549_, _11288_);
  or (_14115_, _14114_, _12547_);
  or (_14116_, _14115_, _14113_);
  and (_14117_, _14116_, _12558_);
  nand (_14118_, _06604_, \oc8051_golden_model_1.ACC [5]);
  nor (_14119_, _06604_, \oc8051_golden_model_1.ACC [5]);
  nor (_14120_, _06961_, \oc8051_golden_model_1.ACC [4]);
  or (_14121_, _14120_, _14119_);
  and (_14122_, _14121_, _14118_);
  and (_14123_, _14122_, _12557_);
  and (_14124_, _06181_, _08737_);
  or (_14125_, _06325_, \oc8051_golden_model_1.ACC [6]);
  nor (_14126_, _14125_, _10934_);
  or (_14127_, _14126_, _14124_);
  or (_14128_, _14127_, _14123_);
  or (_14129_, _14128_, _14117_);
  nor (_14130_, _12559_, _12528_);
  and (_14131_, _14130_, _14129_);
  or (_14132_, _14131_, _12254_);
  or (_14133_, _14132_, _14107_);
  or (_14134_, _14133_, _14080_);
  nand (_14135_, _12254_, \oc8051_golden_model_1.PSW [7]);
  and (_14136_, _14135_, _06271_);
  and (_14137_, _14136_, _14134_);
  or (_14138_, _13986_, _08768_);
  and (_14139_, _14138_, _06270_);
  and (_14140_, _14139_, _14050_);
  nor (_14141_, _14140_, _14137_);
  nor (_14142_, _14141_, _06368_);
  and (_14143_, _12970_, \oc8051_golden_model_1.PSW [7]);
  and (_14144_, _14143_, _06368_);
  or (_14145_, _14144_, _14142_);
  and (_14146_, _14145_, _14016_);
  or (_14147_, _14146_, _14015_);
  and (_14148_, _14147_, _14013_);
  and (_14149_, _09006_, _05938_);
  not (_14150_, _14149_);
  and (_14151_, _10722_, _14150_);
  and (_14152_, _14151_, _10719_);
  or (_14153_, _12970_, \oc8051_golden_model_1.PSW [7]);
  nand (_14154_, _14153_, _06370_);
  nand (_14155_, _14154_, _14152_);
  or (_14156_, _14155_, _14148_);
  and (_14157_, _10739_, _10735_);
  nor (_14158_, _14157_, _10733_);
  nand (_14159_, _10787_, _10735_);
  or (_14160_, _14159_, _10785_);
  and (_14161_, _14160_, _14158_);
  or (_14162_, _14161_, _10729_);
  and (_14163_, _14162_, _06803_);
  or (_14164_, _14163_, _10724_);
  and (_14165_, _14164_, _14156_);
  and (_14166_, _14162_, _06802_);
  or (_14167_, _14166_, _10727_);
  or (_14168_, _14167_, _14165_);
  and (_14169_, _14168_, _14012_);
  or (_14170_, _14169_, _06380_);
  and (_14171_, _10504_, _10500_);
  nor (_14172_, _14171_, _10498_);
  nand (_14173_, _10546_, _10500_);
  or (_14174_, _14173_, _10544_);
  and (_14175_, _14174_, _14172_);
  and (_14176_, _10494_, _08026_);
  or (_14177_, _14176_, _06386_);
  or (_14178_, _14177_, _14175_);
  and (_14179_, _14178_, _10487_);
  and (_14180_, _14179_, _14170_);
  and (_14181_, _10812_, _10809_);
  nor (_14182_, _14181_, _10807_);
  nand (_14183_, _10856_, _10809_);
  or (_14184_, _14183_, _10854_);
  and (_14185_, _14184_, _14182_);
  or (_14186_, _14185_, _10802_);
  and (_14187_, _14186_, _10486_);
  or (_14188_, _14187_, _06259_);
  or (_14189_, _14188_, _14180_);
  and (_14190_, _14189_, _14004_);
  or (_14191_, _14190_, _09486_);
  and (_14192_, _08731_, _07926_);
  or (_14193_, _13995_, _06258_);
  or (_14194_, _14193_, _14192_);
  and (_14195_, _14194_, _06251_);
  and (_14196_, _14195_, _14191_);
  or (_14197_, _14196_, _14001_);
  nor (_14198_, _09480_, _06330_);
  and (_14199_, _14198_, _14197_);
  nor (_14200_, _12970_, _10774_);
  and (_14201_, _14200_, _06330_);
  or (_14202_, _14201_, _06215_);
  or (_14203_, _14202_, _14199_);
  and (_14204_, _08806_, _07926_);
  or (_14205_, _14204_, _13995_);
  or (_14206_, _14205_, _06216_);
  and (_14207_, _14206_, _14203_);
  or (_14208_, _14207_, _06329_);
  nand (_14209_, _12970_, _10774_);
  or (_14210_, _14209_, _06860_);
  and (_14211_, _14210_, _14208_);
  or (_14212_, _14211_, _06398_);
  and (_14213_, _09034_, _07926_);
  or (_14214_, _14213_, _13995_);
  or (_14215_, _14214_, _09025_);
  and (_14216_, _14215_, _09030_);
  and (_14217_, _14216_, _14212_);
  or (_14218_, _14217_, _13998_);
  and (_14219_, _14218_, _07219_);
  or (_14220_, _13995_, _08026_);
  and (_14221_, _14205_, _06426_);
  and (_14222_, _14221_, _14220_);
  or (_14223_, _14222_, _14219_);
  and (_14224_, _14223_, _07217_);
  and (_14225_, _14037_, _06532_);
  and (_14226_, _14225_, _14220_);
  or (_14227_, _14226_, _06437_);
  or (_14228_, _14227_, _14224_);
  and (_14229_, _09033_, _07926_);
  or (_14230_, _13995_, _07229_);
  or (_14231_, _14230_, _14229_);
  and (_14232_, _14231_, _07231_);
  and (_14233_, _14232_, _14228_);
  not (_14234_, _07926_);
  nor (_14235_, _09041_, _14234_);
  or (_14236_, _14235_, _13995_);
  and (_14237_, _14236_, _06535_);
  or (_14238_, _14237_, _11024_);
  or (_14239_, _14238_, _14233_);
  and (_14240_, _14239_, _13994_);
  or (_14241_, _14240_, _13990_);
  or (_14242_, _11027_, _14010_);
  nor (_14243_, _10565_, _08737_);
  or (_14244_, _14243_, _11076_);
  or (_14245_, _14244_, _14242_);
  and (_14246_, _14245_, _06523_);
  and (_14247_, _14246_, _14241_);
  nor (_14248_, _10497_, _08737_);
  or (_14249_, _14248_, _11105_);
  or (_14250_, _11082_, _14176_);
  or (_14251_, _14250_, _14249_);
  and (_14252_, _14251_, _12770_);
  or (_14253_, _14252_, _14247_);
  and (_14254_, _10806_, \oc8051_golden_model_1.ACC [7]);
  or (_14255_, _14254_, _11133_);
  or (_14256_, _11083_, _10802_);
  or (_14257_, _14256_, _14255_);
  and (_14258_, _14257_, _12775_);
  and (_14259_, _14258_, _14253_);
  and (_14260_, _11111_, \oc8051_golden_model_1.ACC [7]);
  or (_14261_, _14260_, _11184_);
  or (_14262_, _14261_, _14259_);
  and (_14263_, _11177_, _10904_);
  nor (_14264_, _11145_, _10903_);
  nor (_14265_, _14264_, _10902_);
  or (_14266_, _14265_, _11185_);
  or (_14267_, _14266_, _14263_);
  and (_14268_, _14267_, _14262_);
  or (_14269_, _14268_, _11191_);
  and (_14270_, _11228_, _10925_);
  nor (_14271_, _11195_, _10924_);
  nor (_14272_, _14271_, _10923_);
  or (_14273_, _14272_, _11190_);
  or (_14274_, _14273_, _14270_);
  and (_14275_, _14274_, _06293_);
  and (_14276_, _14275_, _14269_);
  not (_14277_, _09041_);
  not (_14278_, _09040_);
  nand (_14279_, _11267_, _14278_);
  and (_14280_, _14279_, _06292_);
  and (_14281_, _14280_, _14277_);
  or (_14282_, _14281_, _10474_);
  or (_14283_, _14282_, _14276_);
  nor (_14284_, _11306_, _10932_);
  or (_14285_, _14284_, _10475_);
  or (_14286_, _14285_, _10933_);
  and (_14287_, _14286_, _14283_);
  or (_14288_, _14287_, _06559_);
  not (_14289_, _11320_);
  or (_14290_, _14034_, _07240_);
  and (_14291_, _14290_, _14289_);
  and (_14292_, _14291_, _14288_);
  and (_14293_, _11320_, \oc8051_golden_model_1.ACC [0]);
  or (_14294_, _14293_, _05932_);
  or (_14295_, _14294_, _14292_);
  and (_14296_, _14295_, _13989_);
  or (_14297_, _14296_, _06566_);
  and (_14298_, _08534_, _07926_);
  or (_14299_, _13995_, _06570_);
  or (_14300_, _14299_, _14298_);
  and (_14301_, _14300_, _01320_);
  and (_14302_, _14301_, _14297_);
  or (_14303_, _14302_, _13985_);
  and (_40337_, _14303_, _42355_);
  nand (_14304_, _09384_, _07261_);
  nand (_14305_, _05991_, _05619_);
  not (_14306_, _07232_);
  or (_14307_, _08374_, _08929_);
  and (_14308_, _14307_, _07230_);
  and (_14309_, _08374_, _08929_);
  not (_14310_, _14309_);
  and (_14311_, _14310_, _14307_);
  and (_14312_, _14311_, _09026_);
  or (_14313_, _08374_, _06778_);
  nor (_14314_, _12891_, _12867_);
  or (_14315_, _14314_, _08585_);
  or (_14316_, _08736_, _07157_);
  nand (_14317_, _07152_, _05619_);
  or (_14318_, _07152_, \oc8051_golden_model_1.ACC [0]);
  and (_14319_, _14318_, _14317_);
  nor (_14320_, _14319_, _08734_);
  nor (_14321_, _14320_, _06287_);
  and (_14322_, _14321_, _14316_);
  nor (_14323_, _08374_, _08733_);
  or (_14324_, _14323_, _14322_);
  and (_14325_, _14324_, _08624_);
  nand (_14326_, _12891_, _12868_);
  and (_14327_, _14326_, _06284_);
  or (_14328_, _14327_, _07460_);
  or (_14329_, _14328_, _14325_);
  nor (_14330_, _05949_, \oc8051_golden_model_1.PC [0]);
  nor (_14331_, _14330_, _07170_);
  and (_14332_, _14331_, _14329_);
  and (_14333_, _07170_, _07135_);
  or (_14334_, _14333_, _07178_);
  or (_14335_, _14334_, _14332_);
  and (_14336_, _14335_, _14315_);
  or (_14337_, _14336_, _06276_);
  and (_14338_, _14337_, _14313_);
  or (_14339_, _14338_, _06273_);
  not (_14340_, _12892_);
  and (_14341_, _14326_, _14340_);
  or (_14342_, _14341_, _06274_);
  and (_14343_, _14342_, _05946_);
  and (_14344_, _14343_, _14339_);
  or (_14345_, _05946_, _05619_);
  nand (_14346_, _06343_, _14345_);
  or (_14347_, _14346_, _14344_);
  or (_14348_, _08374_, _06343_);
  and (_14349_, _14348_, _14347_);
  or (_14350_, _14349_, _07197_);
  and (_14351_, _09384_, _06294_);
  or (_14352_, _14351_, _08372_);
  or (_14353_, _14352_, _08650_);
  and (_14354_, _14353_, _08780_);
  and (_14355_, _14354_, _14350_);
  and (_14356_, _07869_, \oc8051_golden_model_1.PSW [7]);
  and (_14357_, _14356_, _06646_);
  or (_14358_, _14357_, _14314_);
  and (_14359_, _14358_, _07196_);
  or (_14360_, _14359_, _05974_);
  or (_14361_, _14360_, _14355_);
  and (_14362_, _05974_, _05619_);
  nor (_14363_, _14362_, _08793_);
  and (_14364_, _14363_, _14361_);
  and (_14365_, _08793_, _07135_);
  or (_14366_, _14365_, _08797_);
  or (_14367_, _14366_, _14364_);
  or (_14368_, _09384_, _08802_);
  and (_14369_, _14368_, _08801_);
  and (_14370_, _14369_, _14367_);
  nor (_14371_, _08806_, _07157_);
  and (_14372_, _08968_, \oc8051_golden_model_1.TMOD [0]);
  and (_14373_, _08917_, \oc8051_golden_model_1.SCON [0]);
  or (_14374_, _14373_, _14372_);
  and (_14375_, _08942_, \oc8051_golden_model_1.TCON [0]);
  and (_14376_, _08944_, \oc8051_golden_model_1.P1 [0]);
  or (_14377_, _14376_, _14375_);
  or (_14378_, _14377_, _14374_);
  and (_14379_, _08935_, \oc8051_golden_model_1.ACC [0]);
  and (_14380_, _08925_, \oc8051_golden_model_1.B [0]);
  or (_14381_, _14380_, _14379_);
  and (_14382_, _08947_, \oc8051_golden_model_1.P0 [0]);
  and (_14383_, _08932_, \oc8051_golden_model_1.SBUF [0]);
  or (_14384_, _14383_, _14382_);
  or (_14385_, _14384_, _14381_);
  and (_14386_, _08956_, \oc8051_golden_model_1.P2 [0]);
  and (_14387_, _08962_, \oc8051_golden_model_1.IE [0]);
  or (_14388_, _14387_, _14386_);
  and (_14389_, _08959_, \oc8051_golden_model_1.P3 [0]);
  and (_14390_, _08964_, \oc8051_golden_model_1.IP [0]);
  or (_14391_, _14390_, _14389_);
  or (_14392_, _14391_, _14388_);
  and (_14393_, _08951_, \oc8051_golden_model_1.TL0 [0]);
  and (_14394_, _08970_, \oc8051_golden_model_1.PSW [0]);
  or (_14395_, _14394_, _14393_);
  or (_14396_, _14395_, _14392_);
  or (_14397_, _14396_, _14385_);
  or (_14398_, _14397_, _14378_);
  and (_14399_, _08990_, \oc8051_golden_model_1.TL1 [0]);
  and (_14400_, _08982_, \oc8051_golden_model_1.PCON [0]);
  and (_14401_, _08993_, \oc8051_golden_model_1.SP [0]);
  or (_14402_, _14401_, _14400_);
  or (_14403_, _14402_, _14399_);
  and (_14404_, _08996_, \oc8051_golden_model_1.DPL [0]);
  and (_14405_, _08986_, \oc8051_golden_model_1.TH0 [0]);
  or (_14406_, _14405_, _14404_);
  and (_14407_, _08998_, \oc8051_golden_model_1.TH1 [0]);
  and (_14408_, _08978_, \oc8051_golden_model_1.DPH [0]);
  or (_14409_, _14408_, _14407_);
  or (_14410_, _14409_, _14406_);
  or (_14411_, _14410_, _14403_);
  or (_14412_, _14411_, _14398_);
  or (_14413_, _14412_, _14371_);
  and (_14414_, _14413_, _07506_);
  or (_14415_, _14414_, _09016_);
  or (_14416_, _14415_, _14370_);
  nor (_14417_, _09015_, _06248_);
  nor (_14418_, _14417_, _06217_);
  and (_14419_, _14418_, _14416_);
  and (_14420_, _08929_, _06217_);
  or (_14421_, _14420_, _06004_);
  or (_14422_, _14421_, _14419_);
  and (_14423_, _06004_, _05619_);
  nor (_14424_, _14423_, _09026_);
  and (_14425_, _14424_, _14422_);
  or (_14426_, _14425_, _14312_);
  and (_14427_, _14426_, _09039_);
  nor (_14428_, _12533_, _09039_);
  or (_14429_, _14428_, _14427_);
  and (_14430_, _14429_, _09038_);
  and (_14431_, _14309_, _08550_);
  or (_14432_, _14431_, _14430_);
  and (_14433_, _14432_, _08549_);
  and (_14434_, _11254_, _07218_);
  or (_14435_, _14434_, _06013_);
  or (_14436_, _14435_, _14433_);
  and (_14437_, _06013_, _05619_);
  nor (_14438_, _14437_, _07230_);
  and (_14439_, _14438_, _14436_);
  or (_14440_, _14439_, _14308_);
  and (_14441_, _14440_, _14306_);
  nor (_14442_, _12532_, _14306_);
  or (_14443_, _14442_, _06011_);
  or (_14444_, _14443_, _14441_);
  nand (_14445_, _06011_, _05619_);
  and (_14446_, _14445_, _08547_);
  and (_14447_, _14446_, _14444_);
  not (_14448_, _08547_);
  and (_14449_, _14448_, _07157_);
  or (_14450_, _14449_, _07245_);
  or (_14451_, _14450_, _14447_);
  nand (_14452_, _09384_, _07245_);
  and (_14453_, _14452_, _14451_);
  or (_14454_, _14453_, _07241_);
  nand (_14455_, _08374_, _07241_);
  and (_14456_, _14455_, _06433_);
  and (_14457_, _14456_, _14454_);
  and (_14458_, _06432_, _05619_);
  or (_14459_, _14458_, _05991_);
  or (_14460_, _14459_, _14457_);
  and (_14461_, _14460_, _14305_);
  or (_14462_, _14461_, _07251_);
  not (_14463_, _07251_);
  or (_14464_, _14314_, _14463_);
  and (_14465_, _14464_, _09417_);
  and (_14466_, _14465_, _14462_);
  nor (_14467_, _09417_, _07135_);
  or (_14468_, _14467_, _07261_);
  or (_14469_, _14468_, _14466_);
  and (_14470_, _14469_, _14304_);
  or (_14471_, _14470_, _07265_);
  nand (_14472_, _08374_, _07265_);
  and (_14473_, _14472_, _07522_);
  and (_14474_, _14473_, _14471_);
  and (_14475_, _07522_, _07268_);
  nor (_14476_, _14475_, _07524_);
  nor (_14477_, _07694_, _07523_);
  nor (_14478_, _14477_, _07847_);
  and (_14479_, _14478_, _07522_);
  and (_14480_, _14479_, _14476_);
  not (_14481_, _14480_);
  or (_14482_, _14481_, _14474_);
  or (_14483_, _14480_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_14484_, _08645_, _07585_);
  not (_14485_, _14484_);
  and (_14486_, _14485_, _07862_);
  and (_14487_, _14486_, _07273_);
  not (_14488_, _14487_);
  and (_14489_, _14488_, _14483_);
  and (_14490_, _14489_, _14482_);
  and (_14491_, _12342_, _06432_);
  and (_14492_, _12212_, _06433_);
  or (_14493_, _14492_, _14491_);
  and (_14494_, _14493_, _14487_);
  or (_40350_, _14494_, _14490_);
  and (_14495_, _12287_, _06432_);
  and (_14496_, _12162_, _06433_);
  or (_14497_, _14496_, _14495_);
  or (_14498_, _14497_, _14488_);
  or (_14499_, _09423_, _08537_);
  nor (_14500_, _14499_, _09417_);
  and (_14501_, _06011_, _05585_);
  nand (_14502_, _08324_, _07031_);
  nor (_14503_, _08324_, _07031_);
  not (_14504_, _14503_);
  and (_14505_, _14504_, _14502_);
  and (_14506_, _14505_, _09026_);
  not (_14507_, _12838_);
  nand (_14508_, _12837_, _12815_);
  and (_14509_, _14508_, _06273_);
  and (_14510_, _14509_, _14507_);
  nor (_14511_, _12837_, _08255_);
  or (_14512_, _14511_, _08585_);
  or (_14513_, _14499_, _08736_);
  and (_14514_, _07152_, _05585_);
  nor (_14515_, _07152_, _06044_);
  or (_14516_, _14515_, _14514_);
  or (_14517_, _14516_, _08734_);
  and (_14518_, _14517_, _14513_);
  or (_14519_, _14518_, _06287_);
  nor (_14520_, _08630_, _08375_);
  nand (_14521_, _14520_, _06287_);
  and (_14522_, _14521_, _14519_);
  or (_14523_, _14522_, _06284_);
  or (_14524_, _14508_, _08624_);
  and (_14525_, _14524_, _14523_);
  or (_14526_, _14525_, _07460_);
  nor (_14527_, _05949_, _05585_);
  nor (_14528_, _14527_, _07170_);
  and (_14529_, _14528_, _14526_);
  and (_14530_, _09422_, _07170_);
  or (_14531_, _14530_, _07178_);
  or (_14532_, _14531_, _14529_);
  and (_14533_, _14532_, _14512_);
  or (_14534_, _14533_, _06276_);
  nand (_14535_, _08324_, _06276_);
  and (_14536_, _14535_, _06274_);
  and (_14537_, _14536_, _14534_);
  or (_14538_, _14537_, _14510_);
  and (_14539_, _14538_, _05946_);
  or (_14540_, _05946_, \oc8051_golden_model_1.PC [1]);
  nand (_14541_, _06343_, _14540_);
  or (_14542_, _14541_, _14539_);
  nand (_14543_, _08324_, _06344_);
  and (_14544_, _14543_, _14542_);
  or (_14545_, _14544_, _07197_);
  nand (_14546_, _09339_, _06294_);
  nand (_14547_, _14546_, _08322_);
  or (_14548_, _14547_, _08650_);
  and (_14549_, _14548_, _08780_);
  and (_14550_, _14549_, _14545_);
  nand (_14551_, _08255_, _10774_);
  and (_14552_, _14551_, _07196_);
  and (_14553_, _14552_, _14508_);
  or (_14554_, _14553_, _05974_);
  or (_14555_, _14554_, _14550_);
  and (_14556_, _05974_, \oc8051_golden_model_1.PC [1]);
  nor (_14557_, _14556_, _08793_);
  and (_14558_, _14557_, _14555_);
  and (_14559_, _09422_, _08793_);
  or (_14560_, _14559_, _08797_);
  or (_14561_, _14560_, _14558_);
  or (_14562_, _09339_, _08802_);
  and (_14563_, _14562_, _08801_);
  and (_14564_, _14563_, _14561_);
  nor (_14565_, _08806_, _07334_);
  and (_14566_, _08942_, \oc8051_golden_model_1.TCON [1]);
  and (_14567_, _08935_, \oc8051_golden_model_1.ACC [1]);
  or (_14568_, _14567_, _14566_);
  and (_14569_, _08968_, \oc8051_golden_model_1.TMOD [1]);
  and (_14570_, _08951_, \oc8051_golden_model_1.TL0 [1]);
  or (_14571_, _14570_, _14569_);
  or (_14572_, _14571_, _14568_);
  and (_14573_, _08947_, \oc8051_golden_model_1.P0 [1]);
  and (_14574_, _08944_, \oc8051_golden_model_1.P1 [1]);
  or (_14575_, _14574_, _14573_);
  and (_14576_, _08925_, \oc8051_golden_model_1.B [1]);
  and (_14577_, _08970_, \oc8051_golden_model_1.PSW [1]);
  or (_14578_, _14577_, _14576_);
  or (_14579_, _14578_, _14575_);
  and (_14580_, _08962_, \oc8051_golden_model_1.IE [1]);
  and (_14581_, _08964_, \oc8051_golden_model_1.IP [1]);
  or (_14582_, _14581_, _14580_);
  and (_14583_, _08956_, \oc8051_golden_model_1.P2 [1]);
  and (_14584_, _08959_, \oc8051_golden_model_1.P3 [1]);
  or (_14585_, _14584_, _14583_);
  or (_14586_, _14585_, _14582_);
  and (_14587_, _08917_, \oc8051_golden_model_1.SCON [1]);
  and (_14588_, _08932_, \oc8051_golden_model_1.SBUF [1]);
  or (_14589_, _14588_, _14587_);
  or (_14590_, _14589_, _14586_);
  or (_14591_, _14590_, _14579_);
  or (_14592_, _14591_, _14572_);
  and (_14593_, _08998_, \oc8051_golden_model_1.TH1 [1]);
  and (_14594_, _08996_, \oc8051_golden_model_1.DPL [1]);
  and (_14595_, _08978_, \oc8051_golden_model_1.DPH [1]);
  or (_14596_, _14595_, _14594_);
  or (_14597_, _14596_, _14593_);
  and (_14598_, _08990_, \oc8051_golden_model_1.TL1 [1]);
  and (_14599_, _08993_, \oc8051_golden_model_1.SP [1]);
  or (_14600_, _14599_, _14598_);
  and (_14601_, _08982_, \oc8051_golden_model_1.PCON [1]);
  and (_14602_, _08986_, \oc8051_golden_model_1.TH0 [1]);
  or (_14603_, _14602_, _14601_);
  or (_14604_, _14603_, _14600_);
  or (_14605_, _14604_, _14597_);
  or (_14606_, _14605_, _14592_);
  or (_14607_, _14606_, _14565_);
  and (_14608_, _14607_, _07506_);
  or (_14609_, _14608_, _09016_);
  or (_14610_, _14609_, _14564_);
  and (_14611_, _09016_, _06995_);
  nor (_14612_, _14611_, _06217_);
  and (_14613_, _14612_, _14610_);
  not (_14614_, _07031_);
  and (_14615_, _14614_, _06217_);
  or (_14616_, _14615_, _06004_);
  or (_14617_, _14616_, _14613_);
  and (_14618_, _06004_, \oc8051_golden_model_1.PC [1]);
  nor (_14619_, _14618_, _09026_);
  and (_14620_, _14619_, _14617_);
  or (_14621_, _14620_, _14506_);
  and (_14622_, _14621_, _09039_);
  and (_14623_, _11253_, _09031_);
  or (_14624_, _14623_, _14622_);
  and (_14625_, _14624_, _09038_);
  and (_14626_, _14503_, _08550_);
  or (_14627_, _14626_, _14625_);
  and (_14628_, _14627_, _08549_);
  and (_14629_, _11251_, _07218_);
  or (_14630_, _14629_, _06013_);
  or (_14631_, _14630_, _14628_);
  and (_14632_, _06013_, \oc8051_golden_model_1.PC [1]);
  nor (_14633_, _14632_, _07230_);
  and (_14634_, _14633_, _14631_);
  and (_14635_, _14502_, _07230_);
  or (_14636_, _14635_, _07232_);
  or (_14637_, _14636_, _14634_);
  nand (_14638_, _11252_, _07232_);
  and (_14639_, _14638_, _09057_);
  and (_14640_, _14639_, _14637_);
  or (_14641_, _14640_, _14501_);
  and (_14642_, _14641_, _07062_);
  or (_14643_, _14499_, _05927_);
  and (_14644_, _14643_, _07465_);
  or (_14645_, _14644_, _14642_);
  nor (_14646_, _14499_, _07412_);
  nor (_14647_, _14646_, _07486_);
  and (_14648_, _14647_, _14645_);
  and (_14649_, _14643_, _07827_);
  or (_14650_, _14649_, _14648_);
  not (_14651_, _07243_);
  or (_14652_, _14499_, _07411_);
  and (_14653_, _14652_, _14651_);
  and (_14654_, _14653_, _14650_);
  not (_14655_, _07242_);
  nor (_14656_, _09438_, _09385_);
  nand (_14657_, _14656_, _14655_);
  and (_14658_, _14657_, _07245_);
  or (_14659_, _14658_, _14654_);
  nand (_14660_, _14656_, _07242_);
  and (_14661_, _14660_, _09066_);
  and (_14662_, _14661_, _14659_);
  nor (_14663_, _14520_, _09066_);
  or (_14664_, _14663_, _06432_);
  or (_14665_, _14664_, _14662_);
  not (_14666_, _05991_);
  nand (_14667_, _06432_, _06035_);
  and (_14668_, _14667_, _14666_);
  and (_14669_, _14668_, _14665_);
  and (_14670_, _05991_, _05585_);
  or (_14671_, _07251_, _14670_);
  or (_14672_, _14671_, _14669_);
  or (_14673_, _14511_, _14463_);
  and (_14674_, _14673_, _09417_);
  and (_14675_, _14674_, _14672_);
  or (_14676_, _14675_, _14500_);
  and (_14677_, _14676_, _07439_);
  and (_14678_, _14656_, _07261_);
  or (_14679_, _14678_, _07265_);
  or (_14680_, _14679_, _14677_);
  not (_14681_, _07265_);
  or (_14682_, _14520_, _14681_);
  and (_14683_, _14682_, _07522_);
  and (_14684_, _14683_, _14680_);
  and (_14685_, _14684_, _14480_);
  nor (_14686_, _14480_, _07282_);
  or (_14687_, _14686_, _14487_);
  or (_14688_, _14687_, _14685_);
  and (_40351_, _14688_, _14498_);
  not (_14689_, _07260_);
  or (_14690_, _09423_, _08662_);
  nor (_14691_, _09424_, _09417_);
  and (_14692_, _14691_, _14690_);
  and (_14693_, _06060_, _06011_);
  nand (_14694_, _08423_, _06689_);
  nor (_14695_, _08423_, _06689_);
  not (_14696_, _14695_);
  and (_14697_, _14696_, _14694_);
  and (_14698_, _14697_, _09026_);
  nor (_14699_, _12813_, _07949_);
  or (_14700_, _14699_, _08585_);
  and (_14701_, _08630_, _08423_);
  nor (_14702_, _08630_, _08423_);
  or (_14703_, _14702_, _14701_);
  or (_14704_, _14703_, _08733_);
  nor (_14705_, _08537_, _07760_);
  or (_14706_, _14705_, _08538_);
  and (_14707_, _14706_, _08734_);
  and (_14708_, _07152_, _06060_);
  nor (_14709_, _07152_, _10198_);
  or (_14710_, _14709_, _14708_);
  and (_14711_, _14710_, _08736_);
  or (_14712_, _14711_, _06287_);
  or (_14713_, _14712_, _14707_);
  and (_14714_, _14713_, _08624_);
  and (_14715_, _14714_, _14704_);
  nand (_14716_, _12813_, _12791_);
  and (_14717_, _14716_, _06284_);
  or (_14718_, _14717_, _07460_);
  or (_14719_, _14718_, _14715_);
  nor (_14720_, _06060_, _05949_);
  nor (_14721_, _14720_, _07170_);
  and (_14722_, _14721_, _14719_);
  and (_14723_, _08662_, _07170_);
  or (_14724_, _14723_, _07178_);
  or (_14725_, _14724_, _14722_);
  and (_14726_, _14725_, _14700_);
  or (_14727_, _14726_, _06276_);
  nand (_14728_, _08423_, _06276_);
  and (_14729_, _14728_, _06274_);
  and (_14730_, _14729_, _14727_);
  not (_14731_, _12814_);
  and (_14732_, _14716_, _14731_);
  and (_14733_, _14732_, _06273_);
  or (_14734_, _14733_, _14730_);
  and (_14735_, _14734_, _05946_);
  or (_14736_, _06451_, _05946_);
  nand (_14737_, _06343_, _14736_);
  or (_14738_, _14737_, _14735_);
  nand (_14739_, _08423_, _06344_);
  and (_14740_, _14739_, _14738_);
  or (_14741_, _14740_, _07197_);
  nand (_14742_, _09293_, _06294_);
  nand (_14743_, _14742_, _08421_);
  or (_14744_, _14743_, _08650_);
  and (_14745_, _14744_, _08780_);
  and (_14746_, _14745_, _14741_);
  and (_14747_, _07910_, \oc8051_golden_model_1.PSW [7]);
  and (_14748_, _14747_, _06646_);
  or (_14749_, _14748_, _14699_);
  and (_14750_, _14749_, _07196_);
  or (_14751_, _14750_, _05974_);
  or (_14752_, _14751_, _14746_);
  and (_14753_, _06451_, _05974_);
  nor (_14754_, _14753_, _08793_);
  and (_14755_, _14754_, _14752_);
  and (_14756_, _08662_, _08793_);
  or (_14757_, _14756_, _08797_);
  or (_14758_, _14757_, _14755_);
  or (_14759_, _09293_, _08802_);
  and (_14760_, _14759_, _08801_);
  and (_14761_, _14760_, _14758_);
  nor (_14762_, _08806_, _07760_);
  and (_14763_, _08925_, \oc8051_golden_model_1.B [2]);
  and (_14764_, _08935_, \oc8051_golden_model_1.ACC [2]);
  or (_14765_, _14764_, _14763_);
  and (_14766_, _08947_, \oc8051_golden_model_1.P0 [2]);
  and (_14767_, _08944_, \oc8051_golden_model_1.P1 [2]);
  or (_14768_, _14767_, _14766_);
  or (_14769_, _14768_, _14765_);
  and (_14770_, _08968_, \oc8051_golden_model_1.TMOD [2]);
  and (_14771_, _08932_, \oc8051_golden_model_1.SBUF [2]);
  or (_14772_, _14771_, _14770_);
  and (_14773_, _08942_, \oc8051_golden_model_1.TCON [2]);
  and (_14774_, _08917_, \oc8051_golden_model_1.SCON [2]);
  or (_14775_, _14774_, _14773_);
  or (_14776_, _14775_, _14772_);
  and (_14777_, _08956_, \oc8051_golden_model_1.P2 [2]);
  and (_14778_, _08964_, \oc8051_golden_model_1.IP [2]);
  or (_14779_, _14778_, _14777_);
  and (_14780_, _08962_, \oc8051_golden_model_1.IE [2]);
  and (_14781_, _08959_, \oc8051_golden_model_1.P3 [2]);
  or (_14782_, _14781_, _14780_);
  or (_14783_, _14782_, _14779_);
  and (_14784_, _08951_, \oc8051_golden_model_1.TL0 [2]);
  and (_14785_, _08970_, \oc8051_golden_model_1.PSW [2]);
  or (_14786_, _14785_, _14784_);
  or (_14787_, _14786_, _14783_);
  or (_14788_, _14787_, _14776_);
  or (_14789_, _14788_, _14769_);
  and (_14790_, _08986_, \oc8051_golden_model_1.TH0 [2]);
  and (_14791_, _08990_, \oc8051_golden_model_1.TL1 [2]);
  and (_14792_, _08978_, \oc8051_golden_model_1.DPH [2]);
  or (_14793_, _14792_, _14791_);
  or (_14794_, _14793_, _14790_);
  and (_14795_, _08982_, \oc8051_golden_model_1.PCON [2]);
  and (_14796_, _08998_, \oc8051_golden_model_1.TH1 [2]);
  or (_14797_, _14796_, _14795_);
  and (_14798_, _08996_, \oc8051_golden_model_1.DPL [2]);
  and (_14799_, _08993_, \oc8051_golden_model_1.SP [2]);
  or (_14800_, _14799_, _14798_);
  or (_14801_, _14800_, _14797_);
  or (_14802_, _14801_, _14794_);
  or (_14803_, _14802_, _14789_);
  or (_14804_, _14803_, _14762_);
  and (_14805_, _14804_, _07506_);
  or (_14806_, _14805_, _09016_);
  or (_14807_, _14806_, _14761_);
  and (_14808_, _09016_, _06646_);
  nor (_14809_, _14808_, _06217_);
  and (_14810_, _14809_, _14807_);
  and (_14811_, _08980_, _06217_);
  or (_14812_, _14811_, _06004_);
  or (_14813_, _14812_, _14810_);
  and (_14814_, _06451_, _06004_);
  nor (_14815_, _14814_, _09026_);
  and (_14816_, _14815_, _14813_);
  or (_14817_, _14816_, _14698_);
  and (_14818_, _14817_, _09039_);
  and (_14819_, _11250_, _09031_);
  or (_14820_, _14819_, _14818_);
  and (_14821_, _14820_, _09038_);
  and (_14822_, _14695_, _08550_);
  or (_14823_, _14822_, _14821_);
  and (_14824_, _14823_, _08549_);
  and (_14825_, _11248_, _07218_);
  or (_14826_, _14825_, _06013_);
  or (_14827_, _14826_, _14824_);
  and (_14828_, _06451_, _06013_);
  nor (_14829_, _14828_, _07230_);
  and (_14830_, _14829_, _14827_);
  and (_14831_, _14694_, _07230_);
  or (_14832_, _14831_, _07232_);
  or (_14833_, _14832_, _14830_);
  nand (_14834_, _11249_, _07232_);
  and (_14835_, _14834_, _09057_);
  and (_14836_, _14835_, _14833_);
  or (_14837_, _14836_, _14693_);
  and (_14838_, _14837_, _08547_);
  and (_14839_, _14706_, _14448_);
  or (_14840_, _14839_, _14838_);
  and (_14841_, _14840_, _14651_);
  nor (_14842_, _09385_, _09294_);
  or (_14843_, _14842_, _09386_);
  and (_14844_, _14843_, _07243_);
  or (_14845_, _14844_, _14841_);
  and (_14846_, _14845_, _14655_);
  and (_14847_, _14843_, _07242_);
  or (_14848_, _14847_, _14846_);
  and (_14849_, _14848_, _09066_);
  and (_14850_, _14703_, _07241_);
  or (_14851_, _14850_, _06432_);
  or (_14852_, _14851_, _14849_);
  or (_14853_, _12314_, _06433_);
  and (_14854_, _14853_, _14666_);
  and (_14855_, _14854_, _14852_);
  and (_14856_, _06060_, _05991_);
  or (_14857_, _07251_, _14856_);
  or (_14858_, _14857_, _14855_);
  or (_14859_, _14699_, _14463_);
  and (_14860_, _14859_, _09417_);
  and (_14861_, _14860_, _14858_);
  or (_14862_, _14861_, _14692_);
  and (_14863_, _14862_, _14689_);
  nor (_14864_, _09438_, _09293_);
  nor (_14865_, _14864_, _09439_);
  and (_14866_, _14865_, _07260_);
  or (_14867_, _14866_, _14863_);
  and (_14868_, _14867_, _06924_);
  and (_14869_, _14865_, _06923_);
  or (_14870_, _14869_, _07265_);
  or (_14871_, _14870_, _14868_);
  nor (_14872_, _08424_, _08375_);
  nor (_14873_, _14872_, _08425_);
  or (_14874_, _14873_, _14681_);
  and (_14875_, _14874_, _07522_);
  and (_14876_, _14875_, _14871_);
  or (_14877_, _14876_, _14481_);
  or (_14878_, _14480_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_14879_, _14878_, _14488_);
  and (_14880_, _14879_, _14877_);
  not (_14881_, _12156_);
  nor (_14882_, _14881_, _06432_);
  and (_14883_, _12281_, _06432_);
  or (_14884_, _14883_, _14882_);
  and (_14885_, _14884_, _14487_);
  or (_40352_, _14885_, _14880_);
  nor (_14886_, _09424_, _09421_);
  nor (_14887_, _14886_, _09425_);
  and (_14888_, _14887_, _09413_);
  and (_14889_, _06095_, _06011_);
  nand (_14890_, _08279_, _06517_);
  nor (_14891_, _08279_, _06517_);
  not (_14892_, _14891_);
  and (_14893_, _14892_, _14890_);
  and (_14894_, _14893_, _09026_);
  nor (_14895_, _12941_, _08260_);
  or (_14896_, _14895_, _08585_);
  nand (_14897_, _12941_, _12919_);
  or (_14898_, _14897_, _08624_);
  nor (_14899_, _14701_, _08279_);
  or (_14900_, _14899_, _08632_);
  and (_14901_, _14900_, _06287_);
  nor (_14902_, _08538_, _07578_);
  or (_14903_, _14902_, _08539_);
  or (_14904_, _14903_, _08736_);
  and (_14905_, _07152_, _06095_);
  nor (_14906_, _07152_, _10248_);
  or (_14907_, _14906_, _14905_);
  nor (_14908_, _14907_, _08734_);
  nor (_14909_, _14908_, _06287_);
  and (_14910_, _14909_, _14904_);
  or (_14911_, _14910_, _06284_);
  or (_14912_, _14911_, _14901_);
  and (_14913_, _14912_, _14898_);
  or (_14914_, _14913_, _07460_);
  nor (_14915_, _06095_, _05949_);
  nor (_14916_, _14915_, _07170_);
  and (_14917_, _14916_, _14914_);
  and (_14918_, _09421_, _07170_);
  or (_14919_, _14918_, _07178_);
  or (_14920_, _14919_, _14917_);
  and (_14921_, _14920_, _14896_);
  or (_14922_, _14921_, _06276_);
  nand (_14923_, _08279_, _06276_);
  and (_14924_, _14923_, _06274_);
  and (_14925_, _14924_, _14922_);
  not (_14926_, _12942_);
  and (_14927_, _14897_, _14926_);
  and (_14928_, _14927_, _06273_);
  or (_14929_, _14928_, _14925_);
  and (_14930_, _14929_, _05946_);
  or (_14931_, _06456_, _05946_);
  nand (_14932_, _06343_, _14931_);
  or (_14933_, _14932_, _14930_);
  nand (_14934_, _08279_, _06344_);
  and (_14935_, _14934_, _14933_);
  or (_14936_, _14935_, _07197_);
  nand (_14937_, _09247_, _06294_);
  nand (_14938_, _14937_, _08277_);
  or (_14939_, _14938_, _08650_);
  and (_14940_, _14939_, _08780_);
  and (_14941_, _14940_, _14936_);
  and (_14942_, _08787_, _06646_);
  or (_14943_, _14895_, _14942_);
  and (_14944_, _14943_, _07196_);
  or (_14945_, _14944_, _05974_);
  or (_14946_, _14945_, _14941_);
  and (_14947_, _06456_, _05974_);
  nor (_14948_, _14947_, _08793_);
  and (_14949_, _14948_, _14946_);
  and (_14950_, _09421_, _08793_);
  or (_14951_, _14950_, _08797_);
  or (_14952_, _14951_, _14949_);
  or (_14953_, _09247_, _08802_);
  and (_14954_, _14953_, _08801_);
  and (_14955_, _14954_, _14952_);
  nor (_14956_, _08806_, _07578_);
  and (_14957_, _08944_, \oc8051_golden_model_1.P1 [3]);
  and (_14958_, _08970_, \oc8051_golden_model_1.PSW [3]);
  or (_14959_, _14958_, _14957_);
  and (_14960_, _08951_, \oc8051_golden_model_1.TL0 [3]);
  and (_14961_, _08917_, \oc8051_golden_model_1.SCON [3]);
  or (_14962_, _14961_, _14960_);
  or (_14963_, _14962_, _14959_);
  and (_14964_, _08968_, \oc8051_golden_model_1.TMOD [3]);
  and (_14965_, _08925_, \oc8051_golden_model_1.B [3]);
  or (_14966_, _14965_, _14964_);
  and (_14967_, _08947_, \oc8051_golden_model_1.P0 [3]);
  and (_14968_, _08932_, \oc8051_golden_model_1.SBUF [3]);
  or (_14969_, _14968_, _14967_);
  or (_14970_, _14969_, _14966_);
  and (_14971_, _08956_, \oc8051_golden_model_1.P2 [3]);
  and (_14972_, _08962_, \oc8051_golden_model_1.IE [3]);
  or (_14973_, _14972_, _14971_);
  and (_14974_, _08959_, \oc8051_golden_model_1.P3 [3]);
  and (_14975_, _08964_, \oc8051_golden_model_1.IP [3]);
  or (_14976_, _14975_, _14974_);
  or (_14977_, _14976_, _14973_);
  and (_14978_, _08942_, \oc8051_golden_model_1.TCON [3]);
  and (_14979_, _08935_, \oc8051_golden_model_1.ACC [3]);
  or (_14980_, _14979_, _14978_);
  or (_14981_, _14980_, _14977_);
  or (_14982_, _14981_, _14970_);
  or (_14983_, _14982_, _14963_);
  and (_14984_, _08996_, \oc8051_golden_model_1.DPL [3]);
  and (_14985_, _08990_, \oc8051_golden_model_1.TL1 [3]);
  and (_14986_, _08993_, \oc8051_golden_model_1.SP [3]);
  or (_14987_, _14986_, _14985_);
  or (_14988_, _14987_, _14984_);
  and (_14989_, _08982_, \oc8051_golden_model_1.PCON [3]);
  and (_14990_, _08978_, \oc8051_golden_model_1.DPH [3]);
  or (_14991_, _14990_, _14989_);
  and (_14992_, _08986_, \oc8051_golden_model_1.TH0 [3]);
  and (_14993_, _08998_, \oc8051_golden_model_1.TH1 [3]);
  or (_14994_, _14993_, _14992_);
  or (_14995_, _14994_, _14991_);
  or (_14996_, _14995_, _14988_);
  or (_14997_, _14996_, _14983_);
  or (_14998_, _14997_, _14956_);
  and (_14999_, _14998_, _07506_);
  or (_15000_, _14999_, _09016_);
  or (_15001_, _15000_, _14955_);
  and (_15002_, _09016_, _06212_);
  nor (_15003_, _15002_, _06217_);
  and (_15004_, _15003_, _15001_);
  and (_15005_, _08809_, _06217_);
  or (_15006_, _15005_, _06004_);
  or (_15007_, _15006_, _15004_);
  and (_15008_, _06456_, _06004_);
  nor (_15009_, _15008_, _09026_);
  and (_15010_, _15009_, _15007_);
  or (_15011_, _15010_, _14894_);
  and (_15012_, _15011_, _09039_);
  and (_15013_, _12529_, _09031_);
  or (_15014_, _15013_, _15012_);
  and (_15015_, _15014_, _09038_);
  and (_15016_, _14891_, _08550_);
  or (_15017_, _15016_, _15015_);
  and (_15018_, _15017_, _08549_);
  and (_15019_, _11246_, _07218_);
  or (_15020_, _15019_, _06013_);
  or (_15021_, _15020_, _15018_);
  and (_15022_, _06456_, _06013_);
  nor (_15023_, _15022_, _07230_);
  and (_15024_, _15023_, _15021_);
  and (_15025_, _14890_, _07230_);
  or (_15026_, _15025_, _07232_);
  or (_15027_, _15026_, _15024_);
  nand (_15028_, _11247_, _07232_);
  and (_15029_, _15028_, _09057_);
  and (_15030_, _15029_, _15027_);
  or (_15031_, _15030_, _14889_);
  and (_15032_, _15031_, _08546_);
  not (_15033_, _08546_);
  and (_15034_, _14903_, _15033_);
  or (_15035_, _15034_, _07410_);
  or (_15036_, _15035_, _15032_);
  or (_15037_, _14903_, _07411_);
  and (_15038_, _15037_, _14651_);
  and (_15039_, _15038_, _15036_);
  nor (_15040_, _09386_, _09248_);
  or (_15041_, _15040_, _09387_);
  or (_15042_, _15041_, _07242_);
  and (_15043_, _15042_, _07245_);
  or (_15044_, _15043_, _15039_);
  or (_15045_, _15041_, _14655_);
  and (_15046_, _15045_, _09066_);
  and (_15047_, _15046_, _15044_);
  and (_15048_, _14900_, _07241_);
  or (_15049_, _15048_, _06432_);
  or (_15050_, _15049_, _15047_);
  or (_15051_, _12310_, _06433_);
  and (_15052_, _15051_, _14666_);
  and (_15053_, _15052_, _15050_);
  and (_15054_, _06095_, _05991_);
  or (_15055_, _07251_, _15054_);
  or (_15056_, _15055_, _15053_);
  or (_15057_, _14895_, _14463_);
  and (_15058_, _15057_, _09417_);
  and (_15059_, _15058_, _15056_);
  or (_15060_, _15059_, _14888_);
  and (_15061_, _15060_, _07439_);
  or (_15062_, _09439_, _09247_);
  nor (_15063_, _09440_, _07439_);
  and (_15064_, _15063_, _15062_);
  or (_15065_, _15064_, _07265_);
  or (_15066_, _15065_, _15061_);
  nor (_15067_, _08425_, _08280_);
  nor (_15068_, _15067_, _08426_);
  or (_15069_, _15068_, _14681_);
  and (_15070_, _15069_, _07522_);
  and (_15071_, _15070_, _15066_);
  or (_15072_, _15071_, _14481_);
  or (_15073_, _14480_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_15074_, _15073_, _14488_);
  and (_15075_, _15074_, _15072_);
  nor (_15076_, _07861_, _01324_);
  and (_15077_, _15076_, _42355_);
  nor (_15078_, _07861_, _06766_);
  and (_15079_, _15078_, _01320_);
  and (_15080_, _15079_, _42355_);
  nor (_15081_, _07861_, \oc8051_golden_model_1.SP [1]);
  and (_15082_, _15081_, _01320_);
  and (_15083_, _15082_, _42355_);
  nor (_15084_, _15083_, _15080_);
  not (_15085_, _07854_);
  or (_15086_, _07861_, _15085_);
  or (_15087_, _15086_, _01324_);
  or (_15088_, _15087_, rst);
  not (_15089_, _07857_);
  nor (_15090_, _07861_, _15089_);
  and (_15091_, _15090_, _01320_);
  and (_15092_, _15091_, _42355_);
  not (_15093_, _15092_);
  and (_15094_, _15093_, _15088_);
  and (_15095_, _15094_, _15084_);
  and (_15096_, _15095_, _15077_);
  not (_15097_, _07861_);
  and (_15098_, _12276_, _06432_);
  and (_15099_, _12151_, _06433_);
  or (_15100_, _15099_, _15098_);
  and (_15101_, _15100_, _15097_);
  and (_15102_, _15101_, _01320_);
  and (_15103_, _15102_, _42355_);
  and (_15104_, _15103_, _15096_);
  or (_40353_, _15104_, _15075_);
  nor (_15105_, _09440_, _09437_);
  nor (_15106_, _15105_, _09441_);
  or (_15107_, _15106_, _07439_);
  nor (_15108_, _08539_, _08525_);
  or (_15109_, _15108_, _08540_);
  or (_15110_, _15109_, _08546_);
  nand (_15111_, _08879_, _08527_);
  nor (_15112_, _08879_, _08527_);
  not (_15113_, _15112_);
  and (_15114_, _15113_, _15111_);
  and (_15115_, _15114_, _09026_);
  nand (_15116_, _12863_, _12861_);
  or (_15117_, _15116_, _08624_);
  or (_15118_, _15109_, _08736_);
  and (_15119_, _05887_, _06280_);
  or (_15120_, _15119_, _07044_);
  and (_15121_, _12183_, _07152_);
  nor (_15122_, _07152_, _10123_);
  or (_15123_, _15122_, _07341_);
  or (_15124_, _15123_, _15121_);
  or (_15125_, _15124_, _15120_);
  and (_15126_, _15125_, _15118_);
  or (_15127_, _15126_, _07159_);
  or (_15128_, _09437_, _08639_);
  and (_15129_, _15128_, _15127_);
  or (_15130_, _15129_, _06287_);
  and (_15131_, _08632_, _08527_);
  nor (_15132_, _08632_, _08527_);
  or (_15133_, _15132_, _15131_);
  or (_15134_, _15133_, _08733_);
  and (_15135_, _15134_, _15130_);
  or (_15136_, _15135_, _06284_);
  and (_15137_, _15136_, _15117_);
  or (_15138_, _15137_, _07460_);
  nor (_15139_, _12183_, _05949_);
  nor (_15140_, _15139_, _07170_);
  and (_15141_, _15140_, _15138_);
  and (_15142_, _09420_, _07170_);
  or (_15143_, _15142_, _07178_);
  or (_15144_, _15143_, _15141_);
  nor (_15145_, _12862_, _12861_);
  or (_15146_, _15145_, _08585_);
  and (_15147_, _15146_, _15144_);
  or (_15148_, _15147_, _06276_);
  nand (_15149_, _08527_, _06276_);
  and (_15150_, _15149_, _06274_);
  and (_15151_, _15150_, _15148_);
  not (_15152_, _12864_);
  and (_15153_, _15116_, _15152_);
  and (_15154_, _15153_, _06273_);
  or (_15155_, _15154_, _15151_);
  and (_15156_, _15155_, _05946_);
  nand (_15157_, _12183_, _07458_);
  nand (_15158_, _15157_, _06343_);
  or (_15159_, _15158_, _15156_);
  nand (_15160_, _08527_, _06344_);
  and (_15161_, _15160_, _15159_);
  or (_15162_, _15161_, _07197_);
  and (_15164_, _09437_, _06294_);
  nand (_15165_, _08472_, _07197_);
  or (_15166_, _15165_, _15164_);
  and (_15167_, _15166_, _08780_);
  and (_15168_, _15167_, _15162_);
  and (_15169_, _14356_, _06647_);
  or (_15170_, _15169_, _15145_);
  and (_15171_, _15170_, _07196_);
  or (_15172_, _15171_, _05974_);
  or (_15173_, _15172_, _15168_);
  not (_15174_, _05974_);
  nor (_15175_, _12183_, _15174_);
  nor (_15176_, _15175_, _08793_);
  and (_15177_, _15176_, _15173_);
  and (_15178_, _09420_, _08793_);
  or (_15179_, _15178_, _08797_);
  or (_15180_, _15179_, _15177_);
  or (_15181_, _09437_, _08802_);
  and (_15182_, _15181_, _08801_);
  and (_15183_, _15182_, _15180_);
  and (_15184_, _08582_, _09420_);
  and (_15185_, _08942_, \oc8051_golden_model_1.TCON [4]);
  and (_15186_, _08968_, \oc8051_golden_model_1.TMOD [4]);
  or (_15187_, _15186_, _15185_);
  and (_15188_, _08944_, \oc8051_golden_model_1.P1 [4]);
  and (_15189_, _08917_, \oc8051_golden_model_1.SCON [4]);
  or (_15190_, _15189_, _15188_);
  or (_15191_, _15190_, _15187_);
  and (_15192_, _08947_, \oc8051_golden_model_1.P0 [4]);
  and (_15193_, _08951_, \oc8051_golden_model_1.TL0 [4]);
  or (_15194_, _15193_, _15192_);
  and (_15195_, _08932_, \oc8051_golden_model_1.SBUF [4]);
  and (_15196_, _08970_, \oc8051_golden_model_1.PSW [4]);
  or (_15197_, _15196_, _15195_);
  or (_15198_, _15197_, _15194_);
  and (_15199_, _08935_, \oc8051_golden_model_1.ACC [4]);
  and (_15200_, _08925_, \oc8051_golden_model_1.B [4]);
  or (_15201_, _15200_, _15199_);
  and (_15202_, _08962_, \oc8051_golden_model_1.IE [4]);
  and (_15203_, _08964_, \oc8051_golden_model_1.IP [4]);
  or (_15204_, _15203_, _15202_);
  and (_15205_, _08956_, \oc8051_golden_model_1.P2 [4]);
  and (_15206_, _08959_, \oc8051_golden_model_1.P3 [4]);
  or (_15207_, _15206_, _15205_);
  or (_15208_, _15207_, _15204_);
  or (_15209_, _15208_, _15201_);
  or (_15210_, _15209_, _15198_);
  or (_15211_, _15210_, _15191_);
  and (_15212_, _08986_, \oc8051_golden_model_1.TH0 [4]);
  and (_15213_, _08982_, \oc8051_golden_model_1.PCON [4]);
  and (_15214_, _08990_, \oc8051_golden_model_1.TL1 [4]);
  or (_15215_, _15214_, _15213_);
  or (_15216_, _15215_, _15212_);
  and (_15217_, _08996_, \oc8051_golden_model_1.DPL [4]);
  and (_15218_, _08993_, \oc8051_golden_model_1.SP [4]);
  or (_15219_, _15218_, _15217_);
  and (_15220_, _08998_, \oc8051_golden_model_1.TH1 [4]);
  and (_15221_, _08978_, \oc8051_golden_model_1.DPH [4]);
  or (_15222_, _15221_, _15220_);
  or (_15223_, _15222_, _15219_);
  or (_15224_, _15223_, _15216_);
  or (_15225_, _15224_, _15211_);
  or (_15226_, _15225_, _15184_);
  and (_15227_, _15226_, _07506_);
  or (_15228_, _15227_, _09016_);
  or (_15229_, _15228_, _15183_);
  and (_15230_, _09016_, _06961_);
  nor (_15231_, _15230_, _06217_);
  and (_15232_, _15231_, _15229_);
  and (_15233_, _08919_, _06217_);
  or (_15234_, _15233_, _06004_);
  or (_15235_, _15234_, _15232_);
  nor (_15236_, _12183_, _13852_);
  nor (_15237_, _15236_, _09026_);
  and (_15238_, _15237_, _15235_);
  or (_15239_, _15238_, _15115_);
  and (_15240_, _15239_, _09039_);
  and (_15241_, _11245_, _09031_);
  or (_15242_, _15241_, _15240_);
  and (_15243_, _15242_, _09038_);
  and (_15244_, _15112_, _08550_);
  or (_15245_, _15244_, _15243_);
  and (_15246_, _15245_, _08549_);
  and (_15247_, _11242_, _07218_);
  or (_15248_, _15247_, _06013_);
  or (_15249_, _15248_, _15246_);
  not (_15250_, _06013_);
  nor (_15251_, _12183_, _15250_);
  nor (_15252_, _15251_, _07230_);
  and (_15253_, _15252_, _15249_);
  and (_15254_, _15111_, _07230_);
  or (_15255_, _15254_, _07232_);
  or (_15256_, _15255_, _15253_);
  nand (_15257_, _11244_, _07232_);
  and (_15258_, _15257_, _09057_);
  and (_15259_, _15258_, _15256_);
  nand (_15260_, _12183_, _06011_);
  nand (_15261_, _15260_, _08546_);
  or (_15262_, _15261_, _15259_);
  and (_15263_, _15262_, _15110_);
  or (_15264_, _15263_, _07410_);
  or (_15265_, _15109_, _07411_);
  and (_15266_, _15265_, _14651_);
  and (_15267_, _15266_, _15264_);
  nor (_15268_, _09387_, _09202_);
  or (_15269_, _15268_, _09388_);
  or (_15270_, _15269_, _07242_);
  and (_15271_, _15270_, _07245_);
  or (_15272_, _15271_, _15267_);
  or (_15273_, _15269_, _14655_);
  and (_15274_, _15273_, _09066_);
  and (_15275_, _15274_, _15272_);
  and (_15276_, _15133_, _07241_);
  or (_15277_, _15276_, _06432_);
  or (_15278_, _15277_, _15275_);
  or (_15279_, _12307_, _06433_);
  and (_15280_, _15279_, _14666_);
  and (_15281_, _15280_, _15278_);
  and (_15282_, _12183_, _05991_);
  or (_15283_, _15282_, _07251_);
  or (_15284_, _15283_, _15281_);
  or (_15285_, _15145_, _14463_);
  and (_15286_, _15285_, _09417_);
  and (_15287_, _15286_, _15284_);
  or (_15288_, _09425_, _09420_);
  nor (_15289_, _09426_, _09417_);
  and (_15290_, _15289_, _15288_);
  or (_15291_, _15290_, _07261_);
  or (_15292_, _15291_, _15287_);
  and (_15293_, _15292_, _15107_);
  or (_15294_, _15293_, _07265_);
  nor (_15295_, _08528_, _08426_);
  nor (_15296_, _15295_, _08529_);
  or (_15297_, _15296_, _14681_);
  and (_15298_, _15297_, _07522_);
  and (_15299_, _15298_, _15294_);
  or (_15300_, _15299_, _14481_);
  or (_15301_, _14480_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_15302_, _15301_, _14488_);
  and (_15303_, _15302_, _15300_);
  not (_15304_, _12148_);
  nor (_15305_, _15304_, _06432_);
  and (_15306_, _12273_, _06432_);
  or (_15307_, _15306_, _15305_);
  and (_15308_, _15307_, _14487_);
  or (_40354_, _15308_, _15303_);
  and (_15309_, _12178_, _06011_);
  or (_15310_, _08913_, _08231_);
  and (_15311_, _08913_, _08231_);
  not (_15312_, _15311_);
  and (_15313_, _15312_, _15310_);
  and (_15314_, _15313_, _09026_);
  nand (_15315_, _12966_, _12964_);
  or (_15316_, _15315_, _08624_);
  or (_15317_, _09436_, _08639_);
  nor (_15318_, _08540_, _08228_);
  or (_15319_, _15318_, _08541_);
  and (_15320_, _15319_, _08734_);
  nor (_15321_, _07152_, _10152_);
  and (_15322_, _12178_, _07152_);
  or (_15323_, _15322_, _15321_);
  and (_15324_, _15323_, _08736_);
  or (_15325_, _15324_, _07159_);
  or (_15326_, _15325_, _15320_);
  and (_15327_, _15326_, _15317_);
  or (_15328_, _15327_, _06287_);
  nor (_15329_, _15131_, _08230_);
  or (_15330_, _15329_, _08633_);
  or (_15331_, _15330_, _08733_);
  and (_15332_, _15331_, _15328_);
  or (_15333_, _15332_, _06284_);
  and (_15334_, _15333_, _15316_);
  or (_15335_, _15334_, _07460_);
  nor (_15336_, _12178_, _05949_);
  nor (_15337_, _15336_, _07170_);
  and (_15338_, _15337_, _15335_);
  and (_15339_, _09419_, _07170_);
  or (_15340_, _15339_, _07178_);
  or (_15341_, _15340_, _15338_);
  nor (_15342_, _12965_, _12964_);
  or (_15343_, _15342_, _08585_);
  and (_15344_, _15343_, _15341_);
  or (_15345_, _15344_, _06276_);
  nand (_15346_, _08230_, _06276_);
  and (_15347_, _15346_, _06274_);
  and (_15348_, _15347_, _15345_);
  not (_15349_, _12967_);
  and (_15350_, _15315_, _06273_);
  and (_15351_, _15350_, _15349_);
  or (_15352_, _15351_, _15348_);
  and (_15353_, _15352_, _05946_);
  or (_15354_, _12179_, _05946_);
  nand (_15355_, _15354_, _06343_);
  or (_15356_, _15355_, _15353_);
  nand (_15357_, _08230_, _06344_);
  and (_15358_, _15357_, _15356_);
  or (_15359_, _15358_, _07197_);
  and (_15360_, _09436_, _06294_);
  nand (_15361_, _08174_, _07197_);
  or (_15362_, _15361_, _15360_);
  and (_15363_, _15362_, _08780_);
  and (_15364_, _15363_, _15359_);
  nand (_15365_, _12965_, _10774_);
  and (_15366_, _15365_, _07196_);
  and (_15367_, _15366_, _15315_);
  or (_15368_, _15367_, _05974_);
  or (_15369_, _15368_, _15364_);
  and (_15370_, _12179_, _05974_);
  nor (_15371_, _15370_, _08793_);
  and (_15372_, _15371_, _15369_);
  and (_15373_, _09419_, _08793_);
  or (_15374_, _15373_, _08797_);
  or (_15375_, _15374_, _15372_);
  or (_15376_, _09436_, _08802_);
  and (_15377_, _15376_, _08801_);
  and (_15378_, _15377_, _15375_);
  and (_15379_, _08582_, _09419_);
  and (_15380_, _08944_, \oc8051_golden_model_1.P1 [5]);
  and (_15381_, _08917_, \oc8051_golden_model_1.SCON [5]);
  or (_15382_, _15381_, _15380_);
  and (_15383_, _08942_, \oc8051_golden_model_1.TCON [5]);
  and (_15384_, _08951_, \oc8051_golden_model_1.TL0 [5]);
  or (_15385_, _15384_, _15383_);
  or (_15386_, _15385_, _15382_);
  and (_15387_, _08947_, \oc8051_golden_model_1.P0 [5]);
  and (_15388_, _08935_, \oc8051_golden_model_1.ACC [5]);
  or (_15389_, _15388_, _15387_);
  and (_15390_, _08968_, \oc8051_golden_model_1.TMOD [5]);
  and (_15391_, _08925_, \oc8051_golden_model_1.B [5]);
  or (_15392_, _15391_, _15390_);
  or (_15393_, _15392_, _15389_);
  and (_15394_, _08962_, \oc8051_golden_model_1.IE [5]);
  and (_15395_, _08964_, \oc8051_golden_model_1.IP [5]);
  or (_15396_, _15395_, _15394_);
  and (_15397_, _08956_, \oc8051_golden_model_1.P2 [5]);
  and (_15398_, _08959_, \oc8051_golden_model_1.P3 [5]);
  or (_15399_, _15398_, _15397_);
  or (_15400_, _15399_, _15396_);
  and (_15401_, _08932_, \oc8051_golden_model_1.SBUF [5]);
  and (_15402_, _08970_, \oc8051_golden_model_1.PSW [5]);
  or (_15403_, _15402_, _15401_);
  or (_15404_, _15403_, _15400_);
  or (_15405_, _15404_, _15393_);
  or (_15406_, _15405_, _15386_);
  and (_15407_, _08990_, \oc8051_golden_model_1.TL1 [5]);
  and (_15408_, _08986_, \oc8051_golden_model_1.TH0 [5]);
  and (_15409_, _08993_, \oc8051_golden_model_1.SP [5]);
  or (_15410_, _15409_, _15408_);
  or (_15411_, _15410_, _15407_);
  and (_15412_, _08996_, \oc8051_golden_model_1.DPL [5]);
  and (_15413_, _08978_, \oc8051_golden_model_1.DPH [5]);
  or (_15414_, _15413_, _15412_);
  and (_15415_, _08982_, \oc8051_golden_model_1.PCON [5]);
  and (_15416_, _08998_, \oc8051_golden_model_1.TH1 [5]);
  or (_15417_, _15416_, _15415_);
  or (_15418_, _15417_, _15414_);
  or (_15419_, _15418_, _15411_);
  or (_15420_, _15419_, _15406_);
  or (_15421_, _15420_, _15379_);
  and (_15422_, _15421_, _07506_);
  or (_15423_, _15422_, _09016_);
  or (_15424_, _15423_, _15378_);
  and (_15425_, _09016_, _06604_);
  nor (_15426_, _15425_, _06217_);
  and (_15427_, _15426_, _15424_);
  and (_15428_, _08913_, _06217_);
  or (_15429_, _15428_, _06004_);
  or (_15430_, _15429_, _15427_);
  and (_15431_, _12179_, _06004_);
  nor (_15432_, _15431_, _09026_);
  and (_15433_, _15432_, _15430_);
  or (_15434_, _15433_, _15314_);
  and (_15435_, _15434_, _09039_);
  and (_15436_, _12536_, _09031_);
  or (_15437_, _15436_, _15435_);
  and (_15438_, _15437_, _09038_);
  and (_15439_, _15311_, _08550_);
  or (_15440_, _15439_, _15438_);
  and (_15441_, _15440_, _08549_);
  and (_15442_, _11240_, _07218_);
  or (_15443_, _15442_, _06013_);
  or (_15444_, _15443_, _15441_);
  and (_15445_, _12179_, _06013_);
  nor (_15446_, _15445_, _07230_);
  and (_15447_, _15446_, _15444_);
  and (_15448_, _15310_, _07230_);
  or (_15449_, _15448_, _07232_);
  or (_15450_, _15449_, _15447_);
  nand (_15451_, _11241_, _07232_);
  and (_15452_, _15451_, _09057_);
  and (_15453_, _15452_, _15450_);
  or (_15454_, _15453_, _15309_);
  and (_15455_, _15454_, _08546_);
  and (_15456_, _15319_, _15033_);
  or (_15457_, _15456_, _07410_);
  or (_15458_, _15457_, _15455_);
  or (_15459_, _15319_, _07411_);
  and (_15460_, _15459_, _14651_);
  and (_15461_, _15460_, _15458_);
  nor (_15462_, _09388_, _09157_);
  or (_15463_, _15462_, _09389_);
  or (_15464_, _15463_, _07242_);
  and (_15465_, _15464_, _07245_);
  or (_15466_, _15465_, _15461_);
  or (_15467_, _15463_, _14655_);
  and (_15468_, _15467_, _09066_);
  and (_15469_, _15468_, _15466_);
  and (_15470_, _15330_, _07241_);
  or (_15471_, _15470_, _06432_);
  or (_15472_, _15471_, _15469_);
  or (_15473_, _12303_, _06433_);
  and (_15474_, _15473_, _14666_);
  and (_15475_, _15474_, _15472_);
  and (_15476_, _12178_, _05991_);
  or (_15477_, _15476_, _07251_);
  or (_15478_, _15477_, _15475_);
  or (_15479_, _15342_, _14463_);
  and (_15480_, _15479_, _09417_);
  and (_15481_, _15480_, _15478_);
  or (_15482_, _09426_, _09419_);
  nor (_15483_, _09427_, _09417_);
  and (_15484_, _15483_, _15482_);
  or (_15485_, _15484_, _15481_);
  and (_15486_, _15485_, _07439_);
  or (_15487_, _09441_, _09436_);
  nor (_15488_, _09442_, _07439_);
  and (_15489_, _15488_, _15487_);
  or (_15490_, _15489_, _07265_);
  or (_15491_, _15490_, _15486_);
  nor (_15492_, _08529_, _08231_);
  nor (_15493_, _15492_, _08530_);
  or (_15494_, _15493_, _14681_);
  and (_15495_, _15494_, _07522_);
  and (_15496_, _15495_, _15491_);
  or (_15497_, _15496_, _14481_);
  or (_15498_, _14480_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_15499_, _15498_, _14488_);
  and (_15500_, _15499_, _15497_);
  and (_15501_, _12144_, _06433_);
  and (_15502_, _12269_, _06432_);
  or (_15503_, _15502_, _15501_);
  and (_15504_, _15503_, _15097_);
  and (_15505_, _15504_, _01320_);
  and (_15506_, _15505_, _42355_);
  and (_15507_, _15506_, _15096_);
  or (_40357_, _15507_, _15500_);
  or (_15508_, _09427_, _09418_);
  nor (_15509_, _09428_, _09417_);
  and (_15510_, _15509_, _15508_);
  nor (_15511_, _08541_, _08125_);
  or (_15512_, _15511_, _08542_);
  or (_15513_, _15512_, _08546_);
  nand (_15514_, _08844_, _08127_);
  nor (_15515_, _08844_, _08127_);
  not (_15516_, _15515_);
  and (_15517_, _15516_, _15514_);
  and (_15518_, _15517_, _09026_);
  and (_15519_, _09418_, _07170_);
  nor (_15520_, _08633_, _08127_);
  or (_15521_, _15520_, _08634_);
  and (_15522_, _15521_, _06287_);
  or (_15523_, _09435_, _08639_);
  and (_15524_, _15512_, _08734_);
  nor (_15525_, _07152_, _10105_);
  and (_15526_, _12171_, _07152_);
  or (_15527_, _15526_, _15525_);
  and (_15528_, _15527_, _08736_);
  or (_15529_, _15528_, _07159_);
  or (_15530_, _15529_, _15524_);
  and (_15531_, _15530_, _08733_);
  and (_15532_, _15531_, _15523_);
  or (_15533_, _15532_, _15522_);
  and (_15534_, _15533_, _08624_);
  nand (_15535_, _12916_, _12914_);
  and (_15536_, _15535_, _06284_);
  or (_15537_, _15536_, _07460_);
  or (_15538_, _15537_, _15534_);
  nor (_15539_, _12171_, _05949_);
  nor (_15540_, _15539_, _07170_);
  and (_15541_, _15540_, _15538_);
  or (_15542_, _15541_, _15519_);
  and (_15543_, _15542_, _08585_);
  nor (_15544_, _12915_, _12914_);
  and (_15545_, _15544_, _07178_);
  or (_15546_, _15545_, _06276_);
  or (_15547_, _15546_, _15543_);
  nand (_15548_, _08127_, _06276_);
  and (_15549_, _15548_, _06274_);
  and (_15550_, _15549_, _15547_);
  not (_15551_, _12917_);
  and (_15552_, _15535_, _15551_);
  and (_15553_, _15552_, _06273_);
  or (_15554_, _15553_, _15550_);
  and (_15555_, _15554_, _05946_);
  or (_15556_, _12172_, _05946_);
  nand (_15557_, _15556_, _06343_);
  or (_15558_, _15557_, _15555_);
  nand (_15559_, _08127_, _06344_);
  and (_15560_, _15559_, _15558_);
  or (_15561_, _15560_, _07197_);
  and (_15562_, _09435_, _06294_);
  nand (_15563_, _08072_, _07197_);
  or (_15564_, _15563_, _15562_);
  and (_15565_, _15564_, _08780_);
  and (_15566_, _15565_, _15561_);
  and (_15567_, _14747_, _06647_);
  or (_15568_, _15567_, _15544_);
  and (_15569_, _15568_, _07196_);
  or (_15570_, _15569_, _05974_);
  or (_15571_, _15570_, _15566_);
  and (_15572_, _12172_, _05974_);
  nor (_15573_, _15572_, _08793_);
  and (_15574_, _15573_, _15571_);
  and (_15575_, _09418_, _08793_);
  or (_15576_, _15575_, _08797_);
  or (_15577_, _15576_, _15574_);
  or (_15578_, _09435_, _08802_);
  and (_15579_, _15578_, _08801_);
  and (_15580_, _15579_, _15577_);
  and (_15581_, _08582_, _09418_);
  and (_15582_, _08947_, \oc8051_golden_model_1.P0 [6]);
  and (_15583_, _08917_, \oc8051_golden_model_1.SCON [6]);
  or (_15584_, _15583_, _15582_);
  and (_15585_, _08951_, \oc8051_golden_model_1.TL0 [6]);
  and (_15586_, _08932_, \oc8051_golden_model_1.SBUF [6]);
  or (_15587_, _15586_, _15585_);
  or (_15588_, _15587_, _15584_);
  and (_15589_, _08942_, \oc8051_golden_model_1.TCON [6]);
  and (_15590_, _08970_, \oc8051_golden_model_1.PSW [6]);
  or (_15591_, _15590_, _15589_);
  and (_15592_, _08968_, \oc8051_golden_model_1.TMOD [6]);
  and (_15593_, _08925_, \oc8051_golden_model_1.B [6]);
  or (_15594_, _15593_, _15592_);
  or (_15595_, _15594_, _15591_);
  and (_15596_, _08962_, \oc8051_golden_model_1.IE [6]);
  and (_15597_, _08959_, \oc8051_golden_model_1.P3 [6]);
  or (_15598_, _15597_, _15596_);
  and (_15599_, _08956_, \oc8051_golden_model_1.P2 [6]);
  and (_15600_, _08964_, \oc8051_golden_model_1.IP [6]);
  or (_15601_, _15600_, _15599_);
  or (_15602_, _15601_, _15598_);
  and (_15603_, _08944_, \oc8051_golden_model_1.P1 [6]);
  and (_15604_, _08935_, \oc8051_golden_model_1.ACC [6]);
  or (_15605_, _15604_, _15603_);
  or (_15606_, _15605_, _15602_);
  or (_15607_, _15606_, _15595_);
  or (_15608_, _15607_, _15588_);
  and (_15609_, _08996_, \oc8051_golden_model_1.DPL [6]);
  and (_15610_, _08982_, \oc8051_golden_model_1.PCON [6]);
  and (_15611_, _08990_, \oc8051_golden_model_1.TL1 [6]);
  or (_15612_, _15611_, _15610_);
  or (_15613_, _15612_, _15609_);
  and (_15614_, _08998_, \oc8051_golden_model_1.TH1 [6]);
  and (_15615_, _08993_, \oc8051_golden_model_1.SP [6]);
  or (_15616_, _15615_, _15614_);
  and (_15617_, _08986_, \oc8051_golden_model_1.TH0 [6]);
  and (_15618_, _08978_, \oc8051_golden_model_1.DPH [6]);
  or (_15619_, _15618_, _15617_);
  or (_15620_, _15619_, _15616_);
  or (_15621_, _15620_, _15613_);
  or (_15622_, _15621_, _15608_);
  or (_15623_, _15622_, _15581_);
  and (_15624_, _15623_, _07506_);
  or (_15625_, _15624_, _09016_);
  or (_15626_, _15625_, _15580_);
  and (_15627_, _09016_, _06325_);
  nor (_15628_, _15627_, _06217_);
  and (_15629_, _15628_, _15626_);
  and (_15630_, _08845_, _06217_);
  or (_15631_, _15630_, _06004_);
  or (_15632_, _15631_, _15629_);
  and (_15633_, _12172_, _06004_);
  nor (_15634_, _15633_, _09026_);
  and (_15635_, _15634_, _15632_);
  or (_15636_, _15635_, _15518_);
  and (_15637_, _15636_, _09039_);
  and (_15638_, _11239_, _09031_);
  or (_15639_, _15638_, _15637_);
  and (_15640_, _15639_, _09038_);
  and (_15641_, _15515_, _08550_);
  or (_15642_, _15641_, _15640_);
  and (_15643_, _15642_, _08549_);
  and (_15644_, _11236_, _07218_);
  or (_15645_, _15644_, _06013_);
  or (_15646_, _15645_, _15643_);
  and (_15647_, _12172_, _06013_);
  nor (_15648_, _15647_, _07230_);
  and (_15649_, _15648_, _15646_);
  and (_15650_, _15514_, _07230_);
  or (_15651_, _15650_, _07232_);
  or (_15652_, _15651_, _15649_);
  nand (_15653_, _11238_, _07232_);
  and (_15654_, _15653_, _09057_);
  and (_15655_, _15654_, _15652_);
  nand (_15656_, _12171_, _06011_);
  nand (_15657_, _15656_, _08546_);
  or (_15658_, _15657_, _15655_);
  and (_15659_, _15658_, _15513_);
  or (_15660_, _15659_, _07410_);
  or (_15661_, _15512_, _07411_);
  and (_15662_, _15661_, _14651_);
  and (_15663_, _15662_, _15660_);
  nor (_15664_, _09389_, _09112_);
  or (_15665_, _15664_, _09390_);
  or (_15666_, _15665_, _07242_);
  and (_15667_, _15666_, _07245_);
  or (_15668_, _15667_, _15663_);
  or (_15669_, _15665_, _14655_);
  and (_15670_, _15669_, _09066_);
  and (_15671_, _15670_, _15668_);
  and (_15672_, _15521_, _07241_);
  or (_15673_, _15672_, _06432_);
  or (_15674_, _15673_, _15671_);
  nand (_15675_, _12297_, _06432_);
  and (_15676_, _15675_, _14666_);
  and (_15677_, _15676_, _15674_);
  and (_15678_, _12171_, _05991_);
  or (_15679_, _15678_, _07251_);
  or (_15680_, _15679_, _15677_);
  or (_15681_, _15544_, _14463_);
  and (_15682_, _15681_, _09417_);
  and (_15683_, _15682_, _15680_);
  or (_15684_, _15683_, _15510_);
  and (_15685_, _15684_, _14689_);
  nor (_15686_, _09442_, _09435_);
  nor (_15687_, _15686_, _09443_);
  and (_15688_, _15687_, _07260_);
  or (_15689_, _15688_, _15685_);
  and (_15690_, _15689_, _06924_);
  and (_15691_, _15687_, _06923_);
  or (_15692_, _15691_, _07265_);
  or (_15693_, _15692_, _15690_);
  nor (_15694_, _08530_, _08128_);
  nor (_15695_, _15694_, _08531_);
  or (_15696_, _15695_, _14681_);
  and (_15697_, _15696_, _07522_);
  and (_15698_, _15697_, _15693_);
  or (_15699_, _15698_, _14481_);
  or (_15700_, _14480_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_15701_, _15700_, _14488_);
  and (_15702_, _15701_, _15699_);
  and (_15703_, _12264_, _06432_);
  and (_15704_, _12139_, _06433_);
  or (_15705_, _15704_, _15703_);
  and (_15706_, _15705_, _14487_);
  or (_40358_, _15706_, _15702_);
  nor (_15707_, _14480_, _07970_);
  nor (_15708_, _14481_, _09451_);
  or (_15709_, _15708_, _15707_);
  and (_15710_, _15709_, _14488_);
  and (_15711_, _09475_, _15097_);
  and (_15712_, _15711_, _01320_);
  and (_15713_, _15712_, _42355_);
  and (_15714_, _15096_, _15713_);
  or (_40359_, _15714_, _15710_);
  and (_15715_, _14475_, _07433_);
  and (_15716_, _15715_, _14478_);
  not (_15717_, _15716_);
  or (_15718_, _15717_, _14474_);
  and (_15719_, _07862_, _07854_);
  nor (_15720_, _07863_, _15719_);
  and (_15721_, _15720_, _07862_);
  and (_15722_, _15721_, _07581_);
  not (_15723_, _15722_);
  or (_15724_, _15716_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_15725_, _15724_, _15723_);
  and (_15726_, _15725_, _15718_);
  and (_15727_, _15722_, _14493_);
  or (_40362_, _15727_, _15726_);
  or (_15728_, _15717_, _14684_);
  or (_15729_, _15716_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_15730_, _15729_, _15723_);
  and (_15731_, _15730_, _15728_);
  and (_15732_, _14497_, _15097_);
  and (_15733_, _15732_, _01320_);
  and (_15734_, _15733_, _42355_);
  not (_15735_, _15080_);
  nor (_15736_, _15083_, _15735_);
  and (_15737_, _15736_, _15094_);
  and (_15738_, _15737_, _15734_);
  or (_40365_, _15738_, _15731_);
  or (_15739_, _15717_, _14876_);
  and (_15740_, _14486_, _07581_);
  not (_15741_, _15740_);
  or (_15742_, _15716_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_15743_, _15742_, _15741_);
  and (_15744_, _15743_, _15739_);
  and (_15745_, _15740_, _14884_);
  or (_40366_, _15745_, _15744_);
  or (_15746_, _15717_, _15071_);
  or (_15747_, _15716_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_15748_, _15747_, _15741_);
  and (_15749_, _15748_, _15746_);
  and (_15750_, _15737_, _15103_);
  or (_40367_, _15750_, _15749_);
  or (_15751_, _15717_, _15299_);
  or (_15752_, _15716_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_15753_, _15752_, _15741_);
  and (_15754_, _15753_, _15751_);
  and (_15755_, _15307_, _15097_);
  and (_15756_, _15755_, _01320_);
  and (_15757_, _15756_, _42355_);
  and (_15758_, _15737_, _15757_);
  or (_40368_, _15758_, _15754_);
  or (_15759_, _15717_, _15496_);
  or (_15760_, _15716_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_15761_, _15760_, _15741_);
  and (_15762_, _15761_, _15759_);
  and (_15763_, _15737_, _15506_);
  or (_40369_, _15763_, _15762_);
  or (_15764_, _15717_, _15698_);
  or (_15765_, _15716_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_15766_, _15765_, _15741_);
  and (_15767_, _15766_, _15764_);
  and (_15768_, _15705_, _15097_);
  and (_15769_, _15768_, _01320_);
  and (_15770_, _15769_, _42355_);
  and (_15771_, _15737_, _15770_);
  or (_40371_, _15771_, _15767_);
  or (_15772_, _15717_, _09452_);
  or (_15773_, _15716_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_15774_, _15773_, _15741_);
  and (_15775_, _15774_, _15772_);
  and (_15776_, _15737_, _15713_);
  or (_40372_, _15776_, _15775_);
  and (_15777_, _14486_, _08641_);
  not (_15778_, _15777_);
  or (_15779_, _15778_, _14493_);
  not (_15780_, _07524_);
  nor (_15781_, _15780_, _07268_);
  and (_15782_, _15781_, _14478_);
  and (_15783_, _15782_, _14474_);
  nor (_15784_, _15782_, _07085_);
  or (_15785_, _15784_, _15777_);
  or (_15786_, _15785_, _15783_);
  and (_40376_, _15786_, _15779_);
  not (_15787_, _15782_);
  or (_15788_, _15787_, _14684_);
  or (_15789_, _15782_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_15790_, _15789_, _15778_);
  and (_15791_, _15790_, _15788_);
  and (_15792_, _15083_, _15735_);
  and (_15793_, _15792_, _15094_);
  and (_15794_, _15793_, _15734_);
  or (_40377_, _15794_, _15791_);
  nor (_15795_, _15782_, _07712_);
  and (_15796_, _15782_, _14876_);
  or (_15797_, _15796_, _15795_);
  and (_15798_, _15797_, _15778_);
  and (_15799_, _15777_, _14884_);
  or (_40379_, _15799_, _15798_);
  or (_15800_, _15787_, _15071_);
  or (_15801_, _15782_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_15802_, _15801_, _15778_);
  and (_15803_, _15802_, _15800_);
  and (_15804_, _15100_, _07862_);
  and (_15805_, _15804_, _15777_);
  or (_40380_, _15805_, _15803_);
  or (_15806_, _15787_, _15299_);
  or (_15807_, _15782_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_15808_, _15807_, _15778_);
  and (_15809_, _15808_, _15806_);
  and (_15810_, _15307_, _07862_);
  and (_15811_, _15810_, _15777_);
  or (_40381_, _15811_, _15809_);
  or (_15812_, _15787_, _15496_);
  or (_15813_, _15782_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_15814_, _15813_, _15778_);
  and (_15815_, _15814_, _15812_);
  and (_15816_, _15503_, _07862_);
  and (_15817_, _15816_, _15777_);
  or (_40382_, _15817_, _15815_);
  or (_15818_, _15787_, _15698_);
  or (_15819_, _15782_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_15820_, _15819_, _15778_);
  and (_15821_, _15820_, _15818_);
  and (_15822_, _15793_, _15770_);
  or (_40383_, _15822_, _15821_);
  or (_15823_, _15787_, _09452_);
  or (_15824_, _15782_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_15825_, _15824_, _15778_);
  and (_15826_, _15825_, _15823_);
  and (_15827_, _15777_, _09476_);
  or (_40385_, _15827_, _15826_);
  and (_15828_, _14486_, _07272_);
  not (_15829_, _15828_);
  or (_15830_, _15829_, _14493_);
  and (_15831_, _14478_, _07525_);
  and (_15832_, _15831_, _14474_);
  nor (_15833_, _15831_, _07082_);
  or (_15834_, _15833_, _15828_);
  or (_15835_, _15834_, _15832_);
  and (_40388_, _15835_, _15830_);
  or (_15836_, _15831_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_15837_, _15836_, _15829_);
  not (_15838_, _15831_);
  or (_15839_, _15838_, _14684_);
  and (_15840_, _15839_, _15837_);
  and (_15841_, _15083_, _15080_);
  and (_15842_, _15094_, _15841_);
  and (_15843_, _15842_, _15734_);
  or (_40390_, _15843_, _15840_);
  nor (_15844_, _15831_, _07710_);
  and (_15845_, _15831_, _14876_);
  or (_15846_, _15845_, _15844_);
  and (_15847_, _15846_, _15829_);
  and (_15848_, _15828_, _14884_);
  or (_40391_, _15848_, _15847_);
  or (_15849_, _15831_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_15850_, _15849_, _15829_);
  or (_15851_, _15838_, _15071_);
  and (_15852_, _15851_, _15850_);
  and (_15853_, _15828_, _15804_);
  or (_40392_, _15853_, _15852_);
  or (_15854_, _15831_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_15855_, _15854_, _15829_);
  or (_15856_, _15838_, _15299_);
  and (_15857_, _15856_, _15855_);
  and (_15858_, _15842_, _15757_);
  or (_40393_, _15858_, _15857_);
  or (_15859_, _15831_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_15860_, _15859_, _15829_);
  or (_15861_, _15838_, _15496_);
  and (_15862_, _15861_, _15860_);
  and (_15863_, _15828_, _15816_);
  or (_40394_, _15863_, _15862_);
  or (_15864_, _15831_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_15865_, _15864_, _15829_);
  or (_15866_, _15838_, _15698_);
  and (_15867_, _15866_, _15865_);
  and (_15868_, _15705_, _07862_);
  and (_15869_, _15868_, _15828_);
  or (_40396_, _15869_, _15867_);
  or (_15870_, _15831_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_15871_, _15870_, _15829_);
  or (_15872_, _15838_, _09452_);
  and (_15873_, _15872_, _15871_);
  and (_15874_, _15828_, _09476_);
  or (_40397_, _15874_, _15873_);
  and (_15875_, _07847_, _07694_);
  and (_15876_, _15875_, _14476_);
  not (_15877_, _15876_);
  or (_15878_, _15877_, _14474_);
  and (_15879_, _15719_, _15089_);
  and (_15880_, _15879_, _07273_);
  not (_15881_, _15880_);
  or (_15882_, _15876_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_15883_, _15882_, _15881_);
  and (_15884_, _15883_, _15878_);
  and (_15885_, _14493_, _07862_);
  and (_15886_, _15885_, _15880_);
  or (_40401_, _15886_, _15884_);
  or (_15887_, _15877_, _14684_);
  or (_15888_, _15876_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_15889_, _15888_, _15881_);
  and (_15890_, _15889_, _15887_);
  and (_15891_, _14497_, _07862_);
  and (_15892_, _15891_, _15880_);
  or (_40402_, _15892_, _15890_);
  or (_15893_, _15877_, _14876_);
  or (_15894_, _15876_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_15895_, _15894_, _15881_);
  and (_15896_, _15895_, _15893_);
  and (_15897_, _14884_, _07862_);
  and (_15898_, _15897_, _15880_);
  or (_40404_, _15898_, _15896_);
  or (_15899_, _15877_, _15071_);
  or (_15900_, _15876_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_15901_, _15900_, _15881_);
  and (_15902_, _15901_, _15899_);
  and (_15903_, _15880_, _15804_);
  or (_40405_, _15903_, _15902_);
  or (_15904_, _15877_, _15299_);
  or (_15905_, _15876_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_15906_, _15905_, _15881_);
  and (_15907_, _15906_, _15904_);
  and (_15908_, _15880_, _15810_);
  or (_40406_, _15908_, _15907_);
  or (_15909_, _15877_, _15496_);
  or (_15910_, _15876_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_15911_, _15910_, _15881_);
  and (_15912_, _15911_, _15909_);
  and (_15913_, _15880_, _15816_);
  or (_40407_, _15913_, _15912_);
  or (_15914_, _15877_, _15698_);
  or (_15915_, _15876_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_15916_, _15915_, _15881_);
  and (_15917_, _15916_, _15914_);
  and (_15918_, _15880_, _15868_);
  or (_40408_, _15918_, _15917_);
  or (_15919_, _15877_, _09452_);
  or (_15920_, _15876_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_15921_, _15920_, _15881_);
  and (_15922_, _15921_, _15919_);
  and (_15923_, _15880_, _09476_);
  or (_40410_, _15923_, _15922_);
  and (_15924_, _15875_, _15715_);
  not (_15925_, _15924_);
  or (_15926_, _15925_, _14474_);
  and (_15927_, _15879_, _07581_);
  not (_15928_, _15927_);
  or (_15929_, _15924_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_15930_, _15929_, _15928_);
  and (_15931_, _15930_, _15926_);
  and (_15932_, _15927_, _15885_);
  or (_40412_, _15932_, _15931_);
  or (_15933_, _15925_, _14684_);
  or (_15934_, _15924_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_15935_, _15934_, _15928_);
  and (_15936_, _15935_, _15933_);
  and (_15937_, _15927_, _15891_);
  or (_40413_, _15937_, _15936_);
  or (_15938_, _15925_, _14876_);
  or (_15939_, _15924_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_15940_, _15939_, _15928_);
  and (_15941_, _15940_, _15938_);
  and (_15942_, _15927_, _15897_);
  or (_40416_, _15942_, _15941_);
  or (_15943_, _15925_, _15071_);
  or (_15944_, _15924_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_15945_, _15944_, _15928_);
  and (_15946_, _15945_, _15943_);
  and (_15947_, _15927_, _15804_);
  or (_40417_, _15947_, _15946_);
  or (_15948_, _15925_, _15299_);
  or (_15949_, _15924_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_15950_, _15949_, _15928_);
  and (_15951_, _15950_, _15948_);
  and (_15952_, _15927_, _15810_);
  or (_40418_, _15952_, _15951_);
  or (_15953_, _15925_, _15496_);
  or (_15954_, _15924_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_15955_, _15954_, _15928_);
  and (_15956_, _15955_, _15953_);
  and (_15957_, _15927_, _15816_);
  or (_40419_, _15957_, _15956_);
  or (_15958_, _15925_, _15698_);
  or (_15959_, _15924_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_15960_, _15959_, _15928_);
  and (_15961_, _15960_, _15958_);
  and (_15962_, _15927_, _15868_);
  or (_40420_, _15962_, _15961_);
  or (_15963_, _15925_, _09452_);
  or (_15964_, _15924_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_15965_, _15964_, _15928_);
  and (_15966_, _15965_, _15963_);
  and (_15967_, _15927_, _09476_);
  or (_40422_, _15967_, _15966_);
  and (_15968_, _15875_, _15781_);
  not (_15969_, _15968_);
  or (_15970_, _15969_, _14474_);
  or (_15971_, _15968_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_15972_, _15879_, _08641_);
  not (_15973_, _15972_);
  and (_15974_, _15973_, _15971_);
  and (_15975_, _15974_, _15970_);
  and (_15976_, _15972_, _15885_);
  or (_40424_, _15976_, _15975_);
  or (_15977_, _15969_, _14684_);
  or (_15978_, _15968_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_15979_, _15978_, _15973_);
  and (_15980_, _15979_, _15977_);
  and (_15981_, _15972_, _15891_);
  or (_40427_, _15981_, _15980_);
  or (_15982_, _15969_, _14876_);
  or (_15983_, _15968_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_15984_, _15983_, _15973_);
  and (_15985_, _15984_, _15982_);
  and (_15986_, _15972_, _15897_);
  or (_40428_, _15986_, _15985_);
  or (_15987_, _15969_, _15071_);
  or (_15988_, _15968_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_15989_, _15988_, _15973_);
  and (_15990_, _15989_, _15987_);
  and (_15991_, _15972_, _15804_);
  or (_40429_, _15991_, _15990_);
  or (_15992_, _15969_, _15299_);
  or (_15993_, _15968_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_15994_, _15993_, _15973_);
  and (_15995_, _15994_, _15992_);
  and (_15996_, _15972_, _15810_);
  or (_40430_, _15996_, _15995_);
  or (_15997_, _15969_, _15496_);
  or (_15998_, _15968_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_15999_, _15998_, _15973_);
  and (_16000_, _15999_, _15997_);
  and (_16001_, _15972_, _15816_);
  or (_40431_, _16001_, _16000_);
  or (_16002_, _15969_, _15698_);
  or (_16003_, _15968_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_16004_, _16003_, _15973_);
  and (_16005_, _16004_, _16002_);
  and (_16006_, _15972_, _15868_);
  or (_40433_, _16006_, _16005_);
  or (_16007_, _15969_, _09452_);
  or (_16008_, _15968_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_16009_, _16008_, _15973_);
  and (_16010_, _16009_, _16007_);
  and (_16011_, _15972_, _09476_);
  or (_40434_, _16011_, _16010_);
  and (_16012_, _15879_, _07272_);
  not (_16013_, _16012_);
  or (_16014_, _16013_, _15885_);
  and (_16015_, _15875_, _07525_);
  nor (_16016_, _16015_, _07092_);
  and (_16017_, _16015_, _14474_);
  or (_16018_, _16017_, _16012_);
  or (_16019_, _16018_, _16016_);
  and (_40437_, _16019_, _16014_);
  or (_16020_, _16015_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_16021_, _16020_, _16013_);
  not (_16022_, _16015_);
  or (_16023_, _16022_, _14684_);
  and (_16024_, _16023_, _16021_);
  and (_16025_, _16012_, _15891_);
  or (_40439_, _16025_, _16024_);
  nor (_16026_, _16015_, _07718_);
  and (_16027_, _16015_, _14876_);
  or (_16028_, _16027_, _16026_);
  and (_16029_, _16028_, _16013_);
  and (_16030_, _16012_, _15897_);
  or (_40440_, _16030_, _16029_);
  or (_16031_, _16015_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_16032_, _16031_, _16013_);
  or (_16033_, _16022_, _15071_);
  and (_16034_, _16033_, _16032_);
  and (_16035_, _16012_, _15804_);
  or (_40441_, _16035_, _16034_);
  or (_16036_, _16015_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_16037_, _16036_, _16013_);
  or (_16038_, _16022_, _15299_);
  and (_16039_, _16038_, _16037_);
  and (_16040_, _16012_, _15810_);
  or (_40442_, _16040_, _16039_);
  or (_16041_, _16015_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_16042_, _16041_, _16013_);
  or (_16043_, _16022_, _15496_);
  and (_16044_, _16043_, _16042_);
  and (_16045_, _16012_, _15816_);
  or (_40443_, _16045_, _16044_);
  or (_16046_, _16015_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_16047_, _16046_, _16013_);
  or (_16048_, _16022_, _15698_);
  and (_16049_, _16048_, _16047_);
  and (_16050_, _16012_, _15868_);
  or (_40445_, _16050_, _16049_);
  or (_16051_, _16015_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_16052_, _16051_, _16013_);
  or (_16053_, _16022_, _09452_);
  and (_16054_, _16053_, _16052_);
  and (_16055_, _16012_, _09476_);
  or (_40446_, _16055_, _16054_);
  and (_16056_, _14477_, _07846_);
  and (_16057_, _16056_, _14476_);
  not (_16058_, _16057_);
  or (_16059_, _16058_, _14474_);
  and (_16060_, _07863_, _15085_);
  and (_16061_, _16060_, _07273_);
  not (_16062_, _16061_);
  or (_16063_, _16057_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_16064_, _16063_, _16062_);
  and (_16065_, _16064_, _16059_);
  and (_16066_, _16061_, _15885_);
  or (_40449_, _16066_, _16065_);
  or (_16067_, _16058_, _14684_);
  or (_16068_, _16057_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_16069_, _16068_, _16062_);
  and (_16070_, _16069_, _16067_);
  and (_16071_, _16061_, _15891_);
  or (_40450_, _16071_, _16070_);
  or (_16072_, _16058_, _14876_);
  or (_16073_, _16057_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_16074_, _16073_, _16062_);
  and (_16075_, _16074_, _16072_);
  and (_16076_, _16061_, _15897_);
  or (_40452_, _16076_, _16075_);
  or (_16077_, _16058_, _15071_);
  or (_16078_, _16057_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_16079_, _16078_, _16062_);
  and (_16080_, _16079_, _16077_);
  and (_16081_, _16061_, _15804_);
  or (_40453_, _16081_, _16080_);
  or (_16082_, _16058_, _15299_);
  or (_16083_, _16057_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_16084_, _16083_, _16062_);
  and (_16085_, _16084_, _16082_);
  and (_16086_, _16061_, _15810_);
  or (_40454_, _16086_, _16085_);
  or (_16087_, _16058_, _15496_);
  or (_16088_, _16057_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_16089_, _16088_, _16062_);
  and (_16090_, _16089_, _16087_);
  and (_16091_, _16061_, _15816_);
  or (_40455_, _16091_, _16090_);
  or (_16092_, _16058_, _15698_);
  or (_16093_, _16057_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_16094_, _16093_, _16062_);
  and (_16095_, _16094_, _16092_);
  and (_16096_, _16061_, _15868_);
  or (_40456_, _16096_, _16095_);
  or (_16097_, _16058_, _09452_);
  or (_16098_, _16057_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_16099_, _16098_, _16062_);
  and (_16100_, _16099_, _16097_);
  and (_16101_, _16061_, _09476_);
  or (_40458_, _16101_, _16100_);
  and (_16102_, _16056_, _15715_);
  not (_16103_, _16102_);
  or (_16104_, _16103_, _14474_);
  and (_16105_, _16060_, _07581_);
  not (_16106_, _16105_);
  or (_16107_, _16102_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_16108_, _16107_, _16106_);
  and (_16109_, _16108_, _16104_);
  and (_16110_, _16105_, _15885_);
  or (_40461_, _16110_, _16109_);
  or (_16111_, _16103_, _14684_);
  or (_16112_, _16102_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_16113_, _16112_, _16106_);
  and (_16114_, _16113_, _16111_);
  and (_16115_, _16105_, _15891_);
  or (_40462_, _16115_, _16114_);
  or (_16116_, _16103_, _14876_);
  or (_16117_, _16102_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_16118_, _16117_, _16106_);
  and (_16119_, _16118_, _16116_);
  and (_16120_, _16105_, _15897_);
  or (_40464_, _16120_, _16119_);
  or (_16121_, _16103_, _15071_);
  or (_16122_, _16102_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_16123_, _16122_, _16106_);
  and (_16124_, _16123_, _16121_);
  and (_16125_, _16105_, _15804_);
  or (_40465_, _16125_, _16124_);
  or (_16126_, _16103_, _15299_);
  or (_16127_, _16102_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_16128_, _16127_, _16106_);
  and (_16129_, _16128_, _16126_);
  and (_16130_, _16105_, _15810_);
  or (_40466_, _16130_, _16129_);
  or (_16131_, _16103_, _15496_);
  or (_16132_, _16102_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_16133_, _16132_, _16106_);
  and (_16134_, _16133_, _16131_);
  and (_16135_, _16105_, _15816_);
  or (_40467_, _16135_, _16134_);
  or (_16136_, _16103_, _15698_);
  or (_16137_, _16102_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_16138_, _16137_, _16106_);
  and (_16139_, _16138_, _16136_);
  and (_16140_, _16105_, _15868_);
  or (_40468_, _16140_, _16139_);
  or (_16141_, _16103_, _09452_);
  or (_16142_, _16102_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_16143_, _16142_, _16106_);
  and (_16144_, _16143_, _16141_);
  and (_16145_, _16105_, _09476_);
  or (_40470_, _16145_, _16144_);
  and (_16146_, _16056_, _15781_);
  nor (_16147_, _16146_, _07111_);
  not (_16148_, _08641_);
  and (_16149_, _15085_, _07857_);
  nand (_16150_, _16149_, _07862_);
  or (_16151_, _16150_, _16148_);
  nand (_16152_, _16146_, _14474_);
  nand (_16153_, _16152_, _16151_);
  or (_16154_, _16153_, _16147_);
  and (_16155_, _16060_, _08641_);
  not (_16156_, _16155_);
  or (_16157_, _16156_, _15885_);
  and (_40473_, _16157_, _16154_);
  not (_16158_, _16146_);
  or (_16159_, _16158_, _14684_);
  or (_16160_, _16146_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_16161_, _16160_, _16156_);
  and (_16162_, _16161_, _16159_);
  and (_16163_, _16155_, _15891_);
  or (_40475_, _16163_, _16162_);
  or (_16164_, _16158_, _14876_);
  or (_16165_, _16146_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_16166_, _16165_, _16156_);
  and (_16167_, _16166_, _16164_);
  and (_16168_, _16155_, _15897_);
  or (_40476_, _16168_, _16167_);
  or (_16169_, _16158_, _15071_);
  or (_16170_, _16146_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_16171_, _16170_, _16156_);
  and (_16172_, _16171_, _16169_);
  and (_16173_, _16155_, _15804_);
  or (_40477_, _16173_, _16172_);
  or (_16174_, _16158_, _15299_);
  or (_16175_, _16146_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_16176_, _16175_, _16156_);
  and (_16177_, _16176_, _16174_);
  and (_16178_, _16155_, _15810_);
  or (_40478_, _16178_, _16177_);
  or (_16179_, _16158_, _15496_);
  or (_16180_, _16146_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_16181_, _16180_, _16156_);
  and (_16182_, _16181_, _16179_);
  and (_16183_, _16155_, _15816_);
  or (_40479_, _16183_, _16182_);
  or (_16184_, _16158_, _15698_);
  or (_16185_, _16146_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_16186_, _16185_, _16156_);
  and (_16187_, _16186_, _16184_);
  and (_16188_, _16155_, _15868_);
  or (_40481_, _16188_, _16187_);
  and (_16189_, _16146_, _09452_);
  or (_16190_, _16146_, _08001_);
  nand (_16191_, _16190_, _16151_);
  or (_16192_, _16191_, _16189_);
  or (_16193_, _16156_, _09476_);
  and (_40482_, _16193_, _16192_);
  not (_16194_, _07272_);
  or (_16195_, _16150_, _16194_);
  or (_16196_, _16195_, _14493_);
  and (_16197_, _16056_, _07525_);
  and (_16198_, _16197_, _14474_);
  or (_16199_, _16197_, _07109_);
  nand (_16200_, _16199_, _16195_);
  or (_16201_, _16200_, _16198_);
  and (_40485_, _16201_, _16196_);
  and (_16202_, _16060_, _07272_);
  not (_16203_, _16202_);
  or (_16204_, _16197_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_16205_, _16204_, _16203_);
  not (_16206_, _16197_);
  or (_16207_, _16206_, _14684_);
  and (_16208_, _16207_, _16205_);
  and (_16209_, _16202_, _15891_);
  or (_40487_, _16209_, _16208_);
  nor (_16210_, _16197_, _07734_);
  and (_16211_, _16197_, _14876_);
  or (_16212_, _16211_, _16210_);
  and (_16213_, _16212_, _16195_);
  and (_16214_, _16202_, _15897_);
  or (_40488_, _16214_, _16213_);
  or (_16215_, _16197_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_16216_, _16215_, _16203_);
  or (_16217_, _16206_, _15071_);
  and (_16218_, _16217_, _16216_);
  and (_16219_, _16202_, _15804_);
  or (_40489_, _16219_, _16218_);
  or (_16220_, _16197_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_16221_, _16220_, _16203_);
  or (_16222_, _16206_, _15299_);
  and (_16223_, _16222_, _16221_);
  and (_16224_, _16202_, _15810_);
  or (_40490_, _16224_, _16223_);
  or (_16225_, _16197_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_16226_, _16225_, _16203_);
  or (_16227_, _16206_, _15496_);
  and (_16228_, _16227_, _16226_);
  and (_16229_, _16202_, _15816_);
  or (_40491_, _16229_, _16228_);
  or (_16230_, _16206_, _15698_);
  or (_16231_, _16197_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_16232_, _16231_, _16203_);
  and (_16233_, _16232_, _16230_);
  and (_16234_, _16202_, _15868_);
  or (_40493_, _16234_, _16233_);
  or (_16235_, _16197_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_16236_, _16235_, _16203_);
  or (_16237_, _16206_, _09452_);
  and (_16238_, _16237_, _16236_);
  and (_16239_, _16202_, _09476_);
  or (_40494_, _16239_, _16238_);
  not (_16240_, _07846_);
  and (_16241_, _14477_, _16240_);
  and (_16242_, _14476_, _16241_);
  not (_16243_, _16242_);
  or (_16244_, _16243_, _14474_);
  and (_16245_, _07864_, _07273_);
  not (_16246_, _16245_);
  or (_16247_, _16242_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_16248_, _16247_, _16246_);
  and (_16249_, _16248_, _16244_);
  and (_16250_, _16245_, _15885_);
  or (_40498_, _16250_, _16249_);
  or (_16251_, _16243_, _14684_);
  or (_16252_, _16242_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_16253_, _16252_, _16246_);
  and (_16254_, _16253_, _16251_);
  and (_16255_, _16245_, _15891_);
  or (_40499_, _16255_, _16254_);
  or (_16256_, _16242_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_16257_, _16256_, _16246_);
  or (_16258_, _16243_, _14876_);
  and (_16259_, _16258_, _16257_);
  and (_16260_, _16245_, _15897_);
  or (_40500_, _16260_, _16259_);
  or (_16261_, _16242_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_16262_, _16261_, _16246_);
  or (_16263_, _16243_, _15071_);
  and (_16264_, _16263_, _16262_);
  and (_16265_, _16245_, _15804_);
  or (_40501_, _16265_, _16264_);
  or (_16266_, _16242_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_16267_, _16266_, _16246_);
  or (_16268_, _16243_, _15299_);
  and (_16269_, _16268_, _16267_);
  and (_16270_, _16245_, _15810_);
  or (_40503_, _16270_, _16269_);
  or (_16271_, _16243_, _15496_);
  or (_16272_, _16242_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_16273_, _16272_, _16246_);
  and (_16274_, _16273_, _16271_);
  and (_16275_, _16245_, _15816_);
  or (_40504_, _16275_, _16274_);
  or (_16276_, _16243_, _15698_);
  or (_16277_, _16242_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_16278_, _16277_, _16246_);
  and (_16279_, _16278_, _16276_);
  and (_16280_, _16245_, _15868_);
  or (_40505_, _16280_, _16279_);
  or (_16281_, _16242_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_16282_, _16281_, _16246_);
  or (_16283_, _16243_, _09452_);
  and (_16284_, _16283_, _16282_);
  and (_16285_, _16245_, _09476_);
  or (_40506_, _16285_, _16284_);
  and (_16286_, _15715_, _16241_);
  not (_16287_, _16286_);
  or (_16288_, _16287_, _14474_);
  and (_16289_, _07864_, _07581_);
  not (_16290_, _16289_);
  or (_16291_, _16286_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_16292_, _16291_, _16290_);
  and (_16293_, _16292_, _16288_);
  and (_16294_, _16289_, _15885_);
  or (_40510_, _16294_, _16293_);
  or (_16295_, _16287_, _14684_);
  or (_16296_, _16286_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_16297_, _16296_, _16290_);
  and (_16298_, _16297_, _16295_);
  and (_16299_, _16289_, _15891_);
  or (_40511_, _16299_, _16298_);
  or (_16300_, _16286_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_16301_, _16300_, _16290_);
  or (_16302_, _16287_, _14876_);
  and (_16303_, _16302_, _16301_);
  and (_16304_, _16289_, _15897_);
  or (_40512_, _16304_, _16303_);
  or (_16305_, _16286_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_16306_, _16305_, _16290_);
  or (_16307_, _16287_, _15071_);
  and (_16308_, _16307_, _16306_);
  and (_16309_, _16289_, _15804_);
  or (_40513_, _16309_, _16308_);
  or (_16310_, _16286_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_16311_, _16310_, _16290_);
  or (_16312_, _16287_, _15299_);
  and (_16313_, _16312_, _16311_);
  and (_16314_, _16289_, _15810_);
  or (_40515_, _16314_, _16313_);
  or (_16315_, _16286_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_16316_, _16315_, _16290_);
  or (_16317_, _16287_, _15496_);
  and (_16318_, _16317_, _16316_);
  and (_16319_, _16289_, _15816_);
  or (_40516_, _16319_, _16318_);
  or (_16320_, _16286_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_16321_, _16320_, _16290_);
  or (_16322_, _16287_, _15698_);
  and (_16323_, _16322_, _16321_);
  and (_16324_, _16289_, _15868_);
  or (_40517_, _16324_, _16323_);
  or (_16325_, _16286_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_16326_, _16325_, _16290_);
  or (_16327_, _16287_, _09452_);
  and (_16328_, _16327_, _16326_);
  and (_16329_, _16289_, _09476_);
  or (_40518_, _16329_, _16328_);
  and (_16330_, _15719_, _07857_);
  nand (_16331_, _08641_, _16330_);
  or (_16332_, _16331_, _15885_);
  and (_16333_, _15781_, _07849_);
  and (_16334_, _16333_, _14474_);
  or (_16335_, _16333_, _07123_);
  nand (_16336_, _16335_, _16331_);
  or (_16337_, _16336_, _16334_);
  and (_40522_, _16337_, _16332_);
  and (_16338_, _08641_, _07864_);
  not (_16339_, _16338_);
  or (_16340_, _16333_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_16341_, _16340_, _16339_);
  not (_16342_, _16333_);
  or (_16343_, _16342_, _14684_);
  and (_16344_, _16343_, _16341_);
  and (_16345_, _16338_, _15891_);
  or (_40523_, _16345_, _16344_);
  nor (_16346_, _16333_, _07748_);
  and (_16347_, _16333_, _14876_);
  or (_16348_, _16347_, _16346_);
  and (_16349_, _16348_, _16331_);
  and (_16350_, _16338_, _15897_);
  or (_40524_, _16350_, _16349_);
  or (_16351_, _16333_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_16352_, _16351_, _16339_);
  or (_16353_, _16342_, _15071_);
  and (_16354_, _16353_, _16352_);
  and (_16355_, _16338_, _15804_);
  or (_40526_, _16355_, _16354_);
  or (_16356_, _16333_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_16357_, _16356_, _16339_);
  or (_16358_, _16342_, _15299_);
  and (_16359_, _16358_, _16357_);
  and (_16360_, _16338_, _15810_);
  or (_40527_, _16360_, _16359_);
  or (_16361_, _16333_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_16362_, _16361_, _16339_);
  or (_16363_, _16342_, _15496_);
  and (_16364_, _16363_, _16362_);
  and (_16365_, _16338_, _15816_);
  or (_40528_, _16365_, _16364_);
  or (_16366_, _16333_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_16367_, _16366_, _16339_);
  or (_16368_, _16342_, _15698_);
  and (_16369_, _16368_, _16367_);
  and (_16370_, _16338_, _15868_);
  or (_40529_, _16370_, _16369_);
  or (_16371_, _16333_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_16372_, _16371_, _16339_);
  or (_16373_, _16342_, _09452_);
  and (_16374_, _16373_, _16372_);
  and (_16375_, _16338_, _09476_);
  or (_40530_, _16375_, _16374_);
  and (_16376_, _16330_, _07272_);
  not (_16377_, _16376_);
  or (_16378_, _15885_, _16377_);
  and (_16379_, _14474_, _07850_);
  nor (_16380_, _07850_, _07121_);
  or (_16381_, _16380_, _16376_);
  or (_16382_, _16381_, _16379_);
  and (_40533_, _16382_, _16378_);
  or (_16383_, _07850_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_16384_, _16383_, _07866_);
  or (_16385_, _14684_, _07868_);
  and (_16386_, _16385_, _16384_);
  and (_16387_, _15891_, _07865_);
  or (_40534_, _16387_, _16386_);
  nor (_16388_, _07850_, _07746_);
  and (_16389_, _14876_, _07850_);
  or (_16390_, _16389_, _16388_);
  and (_16391_, _16390_, _16377_);
  and (_16392_, _15897_, _07865_);
  or (_40535_, _16392_, _16391_);
  or (_16393_, _15071_, _07868_);
  nor (_16394_, _07850_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor (_16395_, _16394_, _16376_);
  and (_16396_, _16395_, _16393_);
  and (_16397_, _15804_, _07865_);
  or (_40537_, _16397_, _16396_);
  or (_16398_, _07850_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_16399_, _16398_, _07866_);
  or (_16400_, _15299_, _07868_);
  and (_16401_, _16400_, _16399_);
  and (_16402_, _15810_, _07865_);
  or (_40538_, _16402_, _16401_);
  nor (_16403_, _07850_, _08215_);
  and (_16404_, _15496_, _07850_);
  or (_16405_, _16404_, _16403_);
  and (_16406_, _16405_, _16377_);
  and (_16407_, _15816_, _16376_);
  or (_40539_, _16407_, _16406_);
  or (_16408_, _07850_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_16409_, _16408_, _07866_);
  or (_16410_, _15698_, _07868_);
  and (_16411_, _16410_, _16409_);
  and (_16412_, _15868_, _07865_);
  or (_40540_, _16412_, _16411_);
  nor (_16413_, _01320_, _10086_);
  nand (_16414_, _11254_, _07933_);
  nor (_16415_, _07933_, _10086_);
  nor (_16416_, _16415_, _07217_);
  nand (_16417_, _16416_, _16414_);
  nor (_16418_, _08374_, _10453_);
  or (_16419_, _16418_, _16415_);
  or (_16420_, _16419_, _06286_);
  and (_16421_, _07933_, \oc8051_golden_model_1.ACC [0]);
  or (_16422_, _16421_, _16415_);
  and (_16423_, _16422_, _07143_);
  nor (_16424_, _07143_, _10086_);
  or (_16425_, _16424_, _06285_);
  or (_16426_, _16425_, _16423_);
  and (_16427_, _16426_, _06282_);
  and (_16428_, _16427_, _16420_);
  and (_16429_, _14326_, _08594_);
  nor (_16430_, _08594_, _10086_);
  or (_16431_, _16430_, _16429_);
  and (_16432_, _16431_, _06281_);
  or (_16433_, _16432_, _16428_);
  and (_16434_, _16433_, _07169_);
  and (_16435_, _07933_, _07135_);
  or (_16436_, _16435_, _16415_);
  and (_16437_, _16436_, _06354_);
  or (_16438_, _16437_, _06345_);
  or (_16439_, _16438_, _16434_);
  or (_16440_, _16422_, _06346_);
  and (_16441_, _16440_, _06278_);
  and (_16442_, _16441_, _16439_);
  and (_16443_, _16415_, _06277_);
  or (_16444_, _16443_, _06270_);
  or (_16445_, _16444_, _16442_);
  or (_16446_, _16419_, _06271_);
  and (_16447_, _16446_, _16445_);
  or (_16448_, _16447_, _09520_);
  nor (_16449_, _10028_, _10026_);
  nor (_16450_, _16449_, _10029_);
  or (_16451_, _16450_, _10059_);
  and (_16452_, _16451_, _06267_);
  and (_16453_, _16452_, _16448_);
  and (_16454_, _14358_, _08594_);
  or (_16455_, _16454_, _16430_);
  and (_16456_, _16455_, _06266_);
  or (_16457_, _16456_, _06259_);
  or (_16458_, _16457_, _16453_);
  or (_16459_, _16436_, _06260_);
  and (_16460_, _16459_, _06258_);
  and (_16461_, _16460_, _16458_);
  and (_16462_, _09384_, _07933_);
  or (_16463_, _16462_, _16415_);
  and (_16464_, _16463_, _09486_);
  or (_16465_, _16464_, _05972_);
  or (_16466_, _16465_, _16461_);
  and (_16467_, _14413_, _07933_);
  or (_16468_, _16415_, _06251_);
  or (_16469_, _16468_, _16467_);
  and (_16470_, _16469_, _09481_);
  and (_16471_, _16470_, _16466_);
  nand (_16472_, _10419_, _06018_);
  and (_16473_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_16474_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_16475_, _16474_, _16473_);
  or (_16476_, _10419_, _16475_);
  and (_16477_, _16476_, _09480_);
  and (_16478_, _16477_, _16472_);
  or (_16479_, _16478_, _10080_);
  or (_16480_, _16479_, _16471_);
  and (_16481_, _14311_, _07933_);
  or (_16482_, _16415_, _09025_);
  or (_16483_, _16482_, _16481_);
  and (_16484_, _07933_, _08929_);
  or (_16485_, _16484_, _16415_);
  or (_16486_, _16485_, _06216_);
  and (_16487_, _16486_, _09030_);
  and (_16488_, _16487_, _16483_);
  and (_16489_, _16488_, _16480_);
  nor (_16490_, _12532_, _10453_);
  or (_16491_, _16490_, _16415_);
  and (_16492_, _16414_, _06524_);
  and (_16493_, _16492_, _16491_);
  or (_16494_, _16493_, _16489_);
  and (_16495_, _16494_, _07219_);
  nand (_16496_, _16485_, _06426_);
  nor (_16497_, _16496_, _16418_);
  or (_16498_, _16497_, _06532_);
  or (_16499_, _16498_, _16495_);
  and (_16500_, _16499_, _16417_);
  or (_16501_, _16500_, _06437_);
  and (_16502_, _14307_, _07933_);
  or (_16503_, _16415_, _07229_);
  or (_16504_, _16503_, _16502_);
  and (_16505_, _16504_, _07231_);
  and (_16506_, _16505_, _16501_);
  and (_16507_, _16491_, _06535_);
  or (_16508_, _16507_, _06559_);
  or (_16509_, _16508_, _16506_);
  or (_16510_, _16419_, _07240_);
  and (_16511_, _16510_, _16509_);
  or (_16512_, _16511_, _05932_);
  or (_16513_, _16415_, _05933_);
  and (_16514_, _16513_, _16512_);
  or (_16515_, _16514_, _06566_);
  or (_16516_, _16419_, _06570_);
  and (_16517_, _16516_, _01320_);
  and (_16518_, _16517_, _16515_);
  or (_16519_, _16518_, _16413_);
  and (_42890_, _16519_, _42355_);
  nor (_16520_, _01320_, _10081_);
  nor (_16521_, _07933_, _10081_);
  nor (_16522_, _11252_, _10453_);
  or (_16523_, _16522_, _16521_);
  or (_16524_, _16523_, _07231_);
  or (_16525_, _07933_, \oc8051_golden_model_1.B [1]);
  nand (_16526_, _07933_, _07031_);
  and (_16527_, _16526_, _06215_);
  and (_16528_, _16527_, _16525_);
  nor (_16529_, _08594_, _10081_);
  and (_16530_, _14511_, _08594_);
  or (_16531_, _16530_, _16529_);
  and (_16532_, _16531_, _06277_);
  and (_16533_, _07933_, _09422_);
  or (_16534_, _16533_, _16521_);
  or (_16535_, _16534_, _07169_);
  and (_16536_, _14520_, _07933_);
  not (_16537_, _16536_);
  and (_16538_, _16537_, _16525_);
  or (_16539_, _16538_, _06286_);
  and (_16540_, _07933_, \oc8051_golden_model_1.ACC [1]);
  or (_16541_, _16540_, _16521_);
  and (_16542_, _16541_, _07143_);
  nor (_16543_, _07143_, _10081_);
  or (_16544_, _16543_, _06285_);
  or (_16545_, _16544_, _16542_);
  and (_16546_, _16545_, _06282_);
  and (_16547_, _16546_, _16539_);
  and (_16548_, _14508_, _08594_);
  or (_16549_, _16548_, _16529_);
  and (_16550_, _16549_, _06281_);
  or (_16551_, _16550_, _06354_);
  or (_16552_, _16551_, _16547_);
  and (_16553_, _16552_, _16535_);
  or (_16554_, _16553_, _06345_);
  or (_16555_, _16541_, _06346_);
  and (_16556_, _16555_, _06278_);
  and (_16557_, _16556_, _16554_);
  or (_16558_, _16557_, _16532_);
  and (_16559_, _16558_, _06271_);
  and (_16560_, _16548_, _14507_);
  or (_16561_, _16560_, _16529_);
  and (_16562_, _16561_, _06270_);
  or (_16563_, _16562_, _09520_);
  or (_16564_, _16563_, _16559_);
  or (_16565_, _09972_, _09971_);
  nand (_16566_, _16565_, _10030_);
  or (_16567_, _16565_, _10030_);
  and (_16568_, _16567_, _16566_);
  or (_16569_, _16568_, _10059_);
  and (_16570_, _16569_, _06267_);
  and (_16571_, _16570_, _16564_);
  or (_16572_, _16529_, _14551_);
  and (_16573_, _16572_, _06266_);
  and (_16574_, _16573_, _16549_);
  or (_16575_, _16574_, _06259_);
  or (_16576_, _16575_, _16571_);
  or (_16577_, _16534_, _06260_);
  and (_16578_, _16577_, _16576_);
  or (_16579_, _16578_, _09486_);
  and (_16580_, _09339_, _07933_);
  or (_16581_, _16521_, _06258_);
  or (_16582_, _16581_, _16580_);
  and (_16583_, _16582_, _06251_);
  and (_16584_, _16583_, _16579_);
  or (_16585_, _14607_, _10453_);
  and (_16586_, _16525_, _05972_);
  and (_16587_, _16586_, _16585_);
  or (_16588_, _16587_, _09480_);
  or (_16589_, _16588_, _16584_);
  nor (_16590_, _10414_, _10413_);
  or (_16591_, _16590_, _10415_);
  nor (_16592_, _16591_, _10419_);
  and (_16593_, _10419_, _10385_);
  or (_16594_, _16593_, _16592_);
  or (_16595_, _16594_, _09481_);
  and (_16596_, _16595_, _06216_);
  and (_16597_, _16596_, _16589_);
  or (_16598_, _16597_, _16528_);
  and (_16599_, _16598_, _09025_);
  or (_16600_, _14505_, _10453_);
  and (_16601_, _16525_, _06398_);
  and (_16602_, _16601_, _16600_);
  or (_16603_, _16602_, _06524_);
  or (_16604_, _16603_, _16599_);
  and (_16605_, _11253_, _07933_);
  or (_16606_, _16605_, _16521_);
  or (_16607_, _16606_, _09030_);
  and (_16608_, _16607_, _07219_);
  and (_16609_, _16608_, _16604_);
  or (_16610_, _14503_, _10453_);
  and (_16611_, _16525_, _06426_);
  and (_16612_, _16611_, _16610_);
  or (_16613_, _16612_, _06532_);
  or (_16614_, _16613_, _16609_);
  and (_16615_, _16540_, _08325_);
  or (_16616_, _16521_, _07217_);
  or (_16617_, _16616_, _16615_);
  and (_16618_, _16617_, _07229_);
  and (_16619_, _16618_, _16614_);
  or (_16620_, _16526_, _08325_);
  and (_16621_, _16525_, _06437_);
  and (_16622_, _16621_, _16620_);
  or (_16623_, _16622_, _06535_);
  or (_16624_, _16623_, _16619_);
  and (_16625_, _16624_, _16524_);
  or (_16626_, _16625_, _06559_);
  or (_16627_, _16538_, _07240_);
  and (_16628_, _16627_, _05933_);
  and (_16629_, _16628_, _16626_);
  and (_16630_, _16531_, _05932_);
  or (_16631_, _16630_, _06566_);
  or (_16632_, _16631_, _16629_);
  or (_16633_, _16521_, _06570_);
  or (_16634_, _16633_, _16536_);
  and (_16635_, _16634_, _01320_);
  and (_16636_, _16635_, _16632_);
  or (_16637_, _16636_, _16520_);
  and (_42891_, _16637_, _42355_);
  nor (_16638_, _01320_, _10096_);
  nor (_16639_, _07933_, _10096_);
  and (_16640_, _07933_, _08662_);
  or (_16641_, _16640_, _16639_);
  or (_16642_, _16641_, _06260_);
  and (_16643_, _14716_, _08594_);
  and (_16644_, _16643_, _14731_);
  nor (_16645_, _08594_, _10096_);
  or (_16646_, _16645_, _06271_);
  or (_16647_, _16646_, _16644_);
  or (_16648_, _16641_, _07169_);
  and (_16649_, _14703_, _07933_);
  or (_16650_, _16649_, _16639_);
  or (_16651_, _16650_, _06286_);
  and (_16652_, _07933_, \oc8051_golden_model_1.ACC [2]);
  or (_16653_, _16652_, _16639_);
  and (_16654_, _16653_, _07143_);
  nor (_16655_, _07143_, _10096_);
  or (_16656_, _16655_, _06285_);
  or (_16657_, _16656_, _16654_);
  and (_16658_, _16657_, _06282_);
  and (_16659_, _16658_, _16651_);
  or (_16660_, _16645_, _16643_);
  and (_16661_, _16660_, _06281_);
  or (_16662_, _16661_, _06354_);
  or (_16663_, _16662_, _16659_);
  and (_16664_, _16663_, _16648_);
  or (_16665_, _16664_, _06345_);
  or (_16666_, _16653_, _06346_);
  and (_16667_, _16666_, _06278_);
  and (_16668_, _16667_, _16665_);
  and (_16669_, _14699_, _08594_);
  or (_16670_, _16669_, _16645_);
  and (_16671_, _16670_, _06277_);
  or (_16672_, _16671_, _06270_);
  or (_16673_, _16672_, _16668_);
  and (_16674_, _16673_, _16647_);
  or (_16675_, _16674_, _09520_);
  or (_16676_, _10032_, _09928_);
  and (_16677_, _16676_, _10033_);
  or (_16678_, _16677_, _10059_);
  and (_16679_, _16678_, _06267_);
  and (_16680_, _16679_, _16675_);
  and (_16681_, _14749_, _08594_);
  or (_16682_, _16681_, _16645_);
  and (_16683_, _16682_, _06266_);
  or (_16684_, _16683_, _06259_);
  or (_16685_, _16684_, _16680_);
  and (_16686_, _16685_, _16642_);
  or (_16687_, _16686_, _09486_);
  and (_16688_, _09293_, _07933_);
  or (_16689_, _16639_, _06258_);
  or (_16690_, _16689_, _16688_);
  and (_16691_, _16690_, _16687_);
  or (_16692_, _16691_, _05972_);
  and (_16693_, _14804_, _07933_);
  or (_16694_, _16639_, _06251_);
  or (_16695_, _16694_, _16693_);
  and (_16696_, _16695_, _09481_);
  and (_16697_, _16696_, _16692_);
  nor (_16698_, _10415_, _10386_);
  not (_16699_, _16698_);
  and (_16700_, _16699_, _10379_);
  nor (_16701_, _16699_, _10379_);
  nor (_16702_, _16701_, _16700_);
  or (_16703_, _16702_, _10419_);
  nand (_16704_, _10419_, _10376_);
  and (_16705_, _16704_, _09480_);
  and (_16706_, _16705_, _16703_);
  or (_16707_, _16706_, _10080_);
  or (_16708_, _16707_, _16697_);
  and (_16709_, _14697_, _07933_);
  or (_16710_, _16639_, _09025_);
  or (_16711_, _16710_, _16709_);
  and (_16712_, _07933_, _08980_);
  or (_16713_, _16712_, _16639_);
  or (_16714_, _16713_, _06216_);
  and (_16715_, _16714_, _09030_);
  and (_16716_, _16715_, _16711_);
  and (_16717_, _16716_, _16708_);
  and (_16718_, _11250_, _07933_);
  or (_16719_, _16718_, _16639_);
  and (_16720_, _16719_, _06524_);
  or (_16721_, _16720_, _16717_);
  and (_16722_, _16721_, _07219_);
  or (_16723_, _16639_, _08424_);
  and (_16724_, _16713_, _06426_);
  and (_16725_, _16724_, _16723_);
  or (_16726_, _16725_, _16722_);
  and (_16727_, _16726_, _07217_);
  and (_16728_, _16653_, _06532_);
  and (_16729_, _16728_, _16723_);
  or (_16730_, _16729_, _06437_);
  or (_16731_, _16730_, _16727_);
  and (_16732_, _14694_, _07933_);
  or (_16733_, _16639_, _07229_);
  or (_16734_, _16733_, _16732_);
  and (_16735_, _16734_, _07231_);
  and (_16736_, _16735_, _16731_);
  nor (_16737_, _11249_, _10453_);
  or (_16738_, _16737_, _16639_);
  and (_16739_, _16738_, _06535_);
  or (_16740_, _16739_, _06559_);
  or (_16741_, _16740_, _16736_);
  or (_16742_, _16650_, _07240_);
  and (_16743_, _16742_, _05933_);
  and (_16744_, _16743_, _16741_);
  and (_16745_, _16670_, _05932_);
  or (_16746_, _16745_, _06566_);
  or (_16747_, _16746_, _16744_);
  and (_16748_, _14873_, _07933_);
  or (_16749_, _16639_, _06570_);
  or (_16750_, _16749_, _16748_);
  and (_16751_, _16750_, _01320_);
  and (_16752_, _16751_, _16747_);
  or (_16753_, _16752_, _16638_);
  and (_42892_, _16753_, _42355_);
  nor (_16754_, _01320_, _10097_);
  nor (_16755_, _07933_, _10097_);
  and (_16756_, _14998_, _07933_);
  or (_16757_, _16756_, _16755_);
  and (_16758_, _16757_, _05972_);
  nor (_16759_, _08594_, _10097_);
  and (_16760_, _14897_, _08594_);
  or (_16761_, _16760_, _16759_);
  or (_16762_, _16759_, _14926_);
  and (_16763_, _16762_, _16761_);
  or (_16764_, _16763_, _06271_);
  and (_16765_, _14900_, _07933_);
  or (_16766_, _16765_, _16755_);
  or (_16767_, _16766_, _06286_);
  and (_16768_, _07933_, \oc8051_golden_model_1.ACC [3]);
  or (_16769_, _16768_, _16755_);
  and (_16770_, _16769_, _07143_);
  nor (_16771_, _07143_, _10097_);
  or (_16772_, _16771_, _06285_);
  or (_16773_, _16772_, _16770_);
  and (_16774_, _16773_, _06282_);
  and (_16775_, _16774_, _16767_);
  and (_16776_, _16761_, _06281_);
  or (_16777_, _16776_, _06354_);
  or (_16778_, _16777_, _16775_);
  and (_16779_, _07933_, _09421_);
  or (_16780_, _16779_, _16755_);
  or (_16781_, _16780_, _07169_);
  and (_16782_, _16781_, _16778_);
  or (_16783_, _16782_, _06345_);
  or (_16784_, _16769_, _06346_);
  and (_16785_, _16784_, _06278_);
  and (_16786_, _16785_, _16783_);
  and (_16787_, _14895_, _08594_);
  or (_16788_, _16787_, _16759_);
  and (_16789_, _16788_, _06277_);
  or (_16790_, _16789_, _06270_);
  or (_16791_, _16790_, _16786_);
  and (_16792_, _16791_, _16764_);
  or (_16793_, _16792_, _09520_);
  nor (_16794_, _10035_, _09870_);
  nor (_16795_, _16794_, _10036_);
  or (_16796_, _16795_, _10059_);
  and (_16797_, _16796_, _06267_);
  and (_16798_, _16797_, _16793_);
  and (_16799_, _14943_, _08594_);
  or (_16800_, _16799_, _16759_);
  and (_16801_, _16800_, _06266_);
  or (_16802_, _16801_, _06259_);
  or (_16803_, _16802_, _16798_);
  or (_16804_, _16780_, _06260_);
  and (_16805_, _16804_, _16803_);
  or (_16806_, _16805_, _09486_);
  and (_16807_, _09247_, _07933_);
  or (_16808_, _16755_, _06258_);
  or (_16809_, _16808_, _16807_);
  and (_16810_, _16809_, _06251_);
  and (_16811_, _16810_, _16806_);
  or (_16812_, _16811_, _16758_);
  and (_16813_, _16812_, _09481_);
  nor (_16814_, _16700_, _10378_);
  nor (_16815_, _16814_, _10371_);
  and (_16816_, _16814_, _10371_);
  or (_16817_, _16816_, _16815_);
  or (_16818_, _16817_, _10419_);
  not (_16819_, _10419_);
  or (_16820_, _16819_, _10368_);
  and (_16821_, _16820_, _09480_);
  and (_16822_, _16821_, _16818_);
  or (_16823_, _16822_, _10080_);
  or (_16824_, _16823_, _16813_);
  and (_16825_, _14893_, _07933_);
  or (_16826_, _16755_, _09025_);
  or (_16827_, _16826_, _16825_);
  and (_16828_, _07933_, _08809_);
  or (_16829_, _16828_, _16755_);
  or (_16830_, _16829_, _06216_);
  and (_16831_, _16830_, _09030_);
  and (_16832_, _16831_, _16827_);
  and (_16833_, _16832_, _16824_);
  and (_16834_, _12529_, _07933_);
  or (_16835_, _16834_, _16755_);
  and (_16836_, _16835_, _06524_);
  or (_16837_, _16836_, _16833_);
  and (_16838_, _16837_, _07219_);
  or (_16839_, _16755_, _08280_);
  and (_16840_, _16829_, _06426_);
  and (_16841_, _16840_, _16839_);
  or (_16842_, _16841_, _16838_);
  and (_16843_, _16842_, _07217_);
  and (_16844_, _16769_, _06532_);
  and (_16845_, _16844_, _16839_);
  or (_16846_, _16845_, _06437_);
  or (_16847_, _16846_, _16843_);
  and (_16848_, _14890_, _07933_);
  or (_16849_, _16755_, _07229_);
  or (_16850_, _16849_, _16848_);
  and (_16851_, _16850_, _07231_);
  and (_16852_, _16851_, _16847_);
  nor (_16853_, _11247_, _10453_);
  or (_16854_, _16853_, _16755_);
  and (_16855_, _16854_, _06535_);
  or (_16856_, _16855_, _06559_);
  or (_16857_, _16856_, _16852_);
  or (_16858_, _16766_, _07240_);
  and (_16859_, _16858_, _05933_);
  and (_16860_, _16859_, _16857_);
  and (_16861_, _16788_, _05932_);
  or (_16862_, _16861_, _06566_);
  or (_16863_, _16862_, _16860_);
  and (_16864_, _15068_, _07933_);
  or (_16865_, _16755_, _06570_);
  or (_16866_, _16865_, _16864_);
  and (_16867_, _16866_, _01320_);
  and (_16868_, _16867_, _16863_);
  or (_16869_, _16868_, _16754_);
  and (_42893_, _16869_, _42355_);
  nor (_16870_, _01320_, _10098_);
  nor (_16871_, _07933_, _10098_);
  and (_16872_, _15226_, _07933_);
  or (_16873_, _16872_, _16871_);
  and (_16874_, _16873_, _05972_);
  and (_16875_, _09420_, _07933_);
  or (_16876_, _16875_, _16871_);
  or (_16877_, _16876_, _06260_);
  nor (_16878_, _08594_, _10098_);
  and (_16879_, _15145_, _08594_);
  or (_16880_, _16879_, _16878_);
  and (_16881_, _16880_, _06277_);
  and (_16882_, _15133_, _07933_);
  or (_16883_, _16882_, _16871_);
  or (_16884_, _16883_, _06286_);
  and (_16885_, _07933_, \oc8051_golden_model_1.ACC [4]);
  or (_16886_, _16885_, _16871_);
  and (_16887_, _16886_, _07143_);
  nor (_16888_, _07143_, _10098_);
  or (_16889_, _16888_, _06285_);
  or (_16890_, _16889_, _16887_);
  and (_16891_, _16890_, _06282_);
  and (_16892_, _16891_, _16884_);
  and (_16893_, _15116_, _08594_);
  or (_16894_, _16893_, _16878_);
  and (_16895_, _16894_, _06281_);
  or (_16896_, _16895_, _06354_);
  or (_16897_, _16896_, _16892_);
  or (_16898_, _16876_, _07169_);
  and (_16899_, _16898_, _16897_);
  or (_16900_, _16899_, _06345_);
  or (_16901_, _16886_, _06346_);
  and (_16902_, _16901_, _06278_);
  and (_16903_, _16902_, _16900_);
  or (_16904_, _16903_, _16881_);
  and (_16905_, _16904_, _06271_);
  or (_16906_, _16878_, _15152_);
  and (_16907_, _16906_, _06270_);
  and (_16908_, _16907_, _16894_);
  or (_16909_, _16908_, _09520_);
  or (_16910_, _16909_, _16905_);
  or (_16911_, _10039_, _10037_);
  and (_16912_, _16911_, _10040_);
  or (_16913_, _16912_, _10059_);
  and (_16914_, _16913_, _06267_);
  and (_16915_, _16914_, _16910_);
  and (_16916_, _15170_, _08594_);
  or (_16917_, _16916_, _16878_);
  and (_16918_, _16917_, _06266_);
  or (_16919_, _16918_, _06259_);
  or (_16920_, _16919_, _16915_);
  and (_16921_, _16920_, _16877_);
  or (_16922_, _16921_, _09486_);
  and (_16923_, _09437_, _07933_);
  or (_16924_, _16871_, _06258_);
  or (_16925_, _16924_, _16923_);
  and (_16926_, _16925_, _06251_);
  and (_16927_, _16926_, _16922_);
  or (_16928_, _16927_, _16874_);
  and (_16929_, _16928_, _09481_);
  or (_16930_, _16819_, _10360_);
  nor (_16931_, _16814_, _10369_);
  or (_16932_, _16931_, _10370_);
  nand (_16933_, _16932_, _10408_);
  or (_16934_, _16932_, _10408_);
  and (_16935_, _16934_, _16933_);
  or (_16936_, _16935_, _10419_);
  and (_16937_, _16936_, _09480_);
  and (_16938_, _16937_, _16930_);
  or (_16939_, _16938_, _10080_);
  or (_16940_, _16939_, _16929_);
  and (_16941_, _15114_, _07933_);
  or (_16942_, _16871_, _09025_);
  or (_16943_, _16942_, _16941_);
  and (_16944_, _08919_, _07933_);
  or (_16945_, _16944_, _16871_);
  or (_16946_, _16945_, _06216_);
  and (_16947_, _16946_, _09030_);
  and (_16948_, _16947_, _16943_);
  and (_16949_, _16948_, _16940_);
  and (_16950_, _11245_, _07933_);
  or (_16951_, _16950_, _16871_);
  and (_16952_, _16951_, _06524_);
  or (_16953_, _16952_, _16949_);
  and (_16954_, _16953_, _07219_);
  or (_16955_, _16871_, _08528_);
  and (_16956_, _16945_, _06426_);
  and (_16957_, _16956_, _16955_);
  or (_16958_, _16957_, _16954_);
  and (_16959_, _16958_, _07217_);
  and (_16960_, _16886_, _06532_);
  and (_16961_, _16960_, _16955_);
  or (_16962_, _16961_, _06437_);
  or (_16963_, _16962_, _16959_);
  and (_16964_, _15111_, _07933_);
  or (_16965_, _16871_, _07229_);
  or (_16966_, _16965_, _16964_);
  and (_16967_, _16966_, _07231_);
  and (_16968_, _16967_, _16963_);
  nor (_16969_, _11244_, _10453_);
  or (_16970_, _16969_, _16871_);
  and (_16971_, _16970_, _06535_);
  or (_16972_, _16971_, _06559_);
  or (_16973_, _16972_, _16968_);
  or (_16974_, _16883_, _07240_);
  and (_16975_, _16974_, _05933_);
  and (_16976_, _16975_, _16973_);
  and (_16977_, _16880_, _05932_);
  or (_16978_, _16977_, _06566_);
  or (_16979_, _16978_, _16976_);
  and (_16980_, _15296_, _07933_);
  or (_16981_, _16871_, _06570_);
  or (_16982_, _16981_, _16980_);
  and (_16983_, _16982_, _01320_);
  and (_16984_, _16983_, _16979_);
  or (_16985_, _16984_, _16870_);
  and (_42894_, _16985_, _42355_);
  nor (_16986_, _01320_, _10099_);
  nor (_16987_, _07933_, _10099_);
  and (_16988_, _15421_, _07933_);
  or (_16989_, _16988_, _16987_);
  and (_16990_, _16989_, _05972_);
  and (_16991_, _09419_, _07933_);
  or (_16992_, _16991_, _16987_);
  or (_16993_, _16992_, _06260_);
  nor (_16994_, _08594_, _10099_);
  and (_16995_, _15342_, _08594_);
  or (_16996_, _16995_, _16994_);
  and (_16997_, _16996_, _06277_);
  and (_16998_, _15330_, _07933_);
  or (_16999_, _16998_, _16987_);
  or (_17000_, _16999_, _06286_);
  and (_17001_, _07933_, \oc8051_golden_model_1.ACC [5]);
  or (_17002_, _17001_, _16987_);
  and (_17003_, _17002_, _07143_);
  nor (_17004_, _07143_, _10099_);
  or (_17005_, _17004_, _06285_);
  or (_17006_, _17005_, _17003_);
  and (_17007_, _17006_, _06282_);
  and (_17008_, _17007_, _17000_);
  and (_17009_, _15315_, _08594_);
  or (_17010_, _17009_, _16994_);
  and (_17011_, _17010_, _06281_);
  or (_17012_, _17011_, _06354_);
  or (_17013_, _17012_, _17008_);
  or (_17014_, _16992_, _07169_);
  and (_17015_, _17014_, _17013_);
  or (_17016_, _17015_, _06345_);
  or (_17017_, _17002_, _06346_);
  and (_17018_, _17017_, _06278_);
  and (_17019_, _17018_, _17016_);
  or (_17020_, _17019_, _16997_);
  and (_17021_, _17020_, _06271_);
  or (_17022_, _16994_, _15349_);
  and (_17023_, _17022_, _06270_);
  and (_17024_, _17023_, _17010_);
  or (_17025_, _17024_, _09520_);
  or (_17026_, _17025_, _17021_);
  nor (_17027_, _10042_, _09731_);
  nor (_17028_, _17027_, _10043_);
  or (_17029_, _17028_, _10059_);
  and (_17030_, _17029_, _06267_);
  and (_17031_, _17030_, _17026_);
  or (_17032_, _16994_, _15365_);
  and (_17033_, _17032_, _06266_);
  and (_17034_, _17033_, _17010_);
  or (_17035_, _17034_, _06259_);
  or (_17036_, _17035_, _17031_);
  and (_17037_, _17036_, _16993_);
  or (_17038_, _17037_, _09486_);
  and (_17039_, _09436_, _07933_);
  or (_17040_, _16987_, _06258_);
  or (_17041_, _17040_, _17039_);
  and (_17042_, _17041_, _06251_);
  and (_17043_, _17042_, _17038_);
  or (_17044_, _17043_, _16990_);
  and (_17045_, _17044_, _09481_);
  not (_17046_, _10397_);
  and (_17047_, _16933_, _17046_);
  nor (_17048_, _17047_, _10409_);
  and (_17049_, _17047_, _10409_);
  or (_17050_, _17049_, _17048_);
  nor (_17051_, _10419_, _09481_);
  and (_17052_, _17051_, _17050_);
  and (_17053_, _10352_, _09480_);
  and (_17054_, _17053_, _10419_);
  or (_17055_, _17054_, _10080_);
  or (_17056_, _17055_, _17052_);
  or (_17057_, _17056_, _17045_);
  and (_17058_, _15313_, _07933_);
  or (_17059_, _16987_, _09025_);
  or (_17060_, _17059_, _17058_);
  and (_17061_, _08913_, _07933_);
  or (_17062_, _17061_, _16987_);
  or (_17063_, _17062_, _06216_);
  and (_17064_, _17063_, _09030_);
  and (_17065_, _17064_, _17060_);
  and (_17066_, _17065_, _17057_);
  and (_17067_, _12536_, _07933_);
  or (_17068_, _17067_, _16987_);
  and (_17069_, _17068_, _06524_);
  or (_17070_, _17069_, _17066_);
  and (_17071_, _17070_, _07219_);
  or (_17072_, _16987_, _08231_);
  and (_17073_, _17062_, _06426_);
  and (_17074_, _17073_, _17072_);
  or (_17075_, _17074_, _17071_);
  and (_17076_, _17075_, _07217_);
  and (_17077_, _17002_, _06532_);
  and (_17078_, _17077_, _17072_);
  or (_17079_, _17078_, _06437_);
  or (_17080_, _17079_, _17076_);
  and (_17081_, _15310_, _07933_);
  or (_17082_, _16987_, _07229_);
  or (_17083_, _17082_, _17081_);
  and (_17084_, _17083_, _07231_);
  and (_17085_, _17084_, _17080_);
  nor (_17086_, _11241_, _10453_);
  or (_17087_, _17086_, _16987_);
  and (_17088_, _17087_, _06535_);
  or (_17089_, _17088_, _06559_);
  or (_17090_, _17089_, _17085_);
  or (_17091_, _16999_, _07240_);
  and (_17092_, _17091_, _05933_);
  and (_17093_, _17092_, _17090_);
  and (_17094_, _16996_, _05932_);
  or (_17095_, _17094_, _06566_);
  or (_17096_, _17095_, _17093_);
  and (_17097_, _15493_, _07933_);
  or (_17098_, _16987_, _06570_);
  or (_17099_, _17098_, _17097_);
  and (_17100_, _17099_, _01320_);
  and (_17101_, _17100_, _17096_);
  or (_17102_, _17101_, _16986_);
  and (_42896_, _17102_, _42355_);
  nor (_17103_, _01320_, _10337_);
  nor (_17104_, _07933_, _10337_);
  and (_17105_, _15623_, _07933_);
  or (_17106_, _17105_, _17104_);
  and (_17107_, _17106_, _05972_);
  and (_17108_, _09418_, _07933_);
  or (_17109_, _17108_, _17104_);
  or (_17110_, _17109_, _06260_);
  nor (_17111_, _08594_, _10337_);
  and (_17112_, _15544_, _08594_);
  or (_17113_, _17112_, _17111_);
  and (_17114_, _17113_, _06277_);
  and (_17115_, _15521_, _07933_);
  or (_17116_, _17115_, _17104_);
  or (_17117_, _17116_, _06286_);
  and (_17118_, _07933_, \oc8051_golden_model_1.ACC [6]);
  or (_17119_, _17118_, _17104_);
  and (_17120_, _17119_, _07143_);
  nor (_17121_, _07143_, _10337_);
  or (_17122_, _17121_, _06285_);
  or (_17123_, _17122_, _17120_);
  and (_17124_, _17123_, _06282_);
  and (_17125_, _17124_, _17117_);
  and (_17126_, _15535_, _08594_);
  or (_17127_, _17126_, _17111_);
  and (_17128_, _17127_, _06281_);
  or (_17129_, _17128_, _06354_);
  or (_17130_, _17129_, _17125_);
  or (_17131_, _17109_, _07169_);
  and (_17132_, _17131_, _17130_);
  or (_17133_, _17132_, _06345_);
  or (_17134_, _17119_, _06346_);
  and (_17135_, _17134_, _06278_);
  and (_17136_, _17135_, _17133_);
  or (_17137_, _17136_, _17114_);
  and (_17138_, _17137_, _06271_);
  or (_17139_, _17111_, _15551_);
  and (_17140_, _17139_, _06270_);
  and (_17141_, _17140_, _17127_);
  or (_17142_, _17141_, _09520_);
  or (_17143_, _17142_, _17138_);
  not (_17144_, _10058_);
  or (_17145_, _10057_, _10044_);
  and (_17146_, _17145_, _17144_);
  or (_17147_, _17146_, _10059_);
  and (_17148_, _17147_, _06267_);
  and (_17149_, _17148_, _17143_);
  and (_17150_, _15568_, _08594_);
  or (_17151_, _17150_, _17111_);
  and (_17152_, _17151_, _06266_);
  or (_17153_, _17152_, _06259_);
  or (_17154_, _17153_, _17149_);
  and (_17155_, _17154_, _17110_);
  or (_17156_, _17155_, _09486_);
  and (_17157_, _09435_, _07933_);
  or (_17158_, _17104_, _06258_);
  or (_17159_, _17158_, _17157_);
  and (_17160_, _17159_, _06251_);
  and (_17161_, _17160_, _17156_);
  or (_17162_, _17161_, _17107_);
  and (_17163_, _17162_, _09481_);
  nor (_17164_, _17047_, _10353_);
  or (_17165_, _17164_, _10354_);
  or (_17166_, _17165_, _10406_);
  nand (_17167_, _17165_, _10406_);
  and (_17168_, _17167_, _17166_);
  or (_17169_, _17168_, _10419_);
  or (_17170_, _16819_, _10343_);
  and (_17171_, _17170_, _09480_);
  and (_17172_, _17171_, _17169_);
  or (_17173_, _17172_, _10080_);
  or (_17174_, _17173_, _17163_);
  and (_17175_, _15517_, _07933_);
  or (_17176_, _17104_, _09025_);
  or (_17177_, _17176_, _17175_);
  and (_17178_, _08845_, _07933_);
  or (_17179_, _17178_, _17104_);
  or (_17180_, _17179_, _06216_);
  and (_17181_, _17180_, _09030_);
  and (_17182_, _17181_, _17177_);
  and (_17183_, _17182_, _17174_);
  and (_17184_, _11239_, _07933_);
  or (_17185_, _17184_, _17104_);
  and (_17186_, _17185_, _06524_);
  or (_17187_, _17186_, _17183_);
  and (_17188_, _17187_, _07219_);
  or (_17189_, _17104_, _08128_);
  and (_17190_, _17179_, _06426_);
  and (_17191_, _17190_, _17189_);
  or (_17192_, _17191_, _17188_);
  and (_17193_, _17192_, _07217_);
  and (_17194_, _17119_, _06532_);
  and (_17195_, _17194_, _17189_);
  or (_17196_, _17195_, _06437_);
  or (_17197_, _17196_, _17193_);
  and (_17198_, _15514_, _07933_);
  or (_17199_, _17104_, _07229_);
  or (_17200_, _17199_, _17198_);
  and (_17201_, _17200_, _07231_);
  and (_17202_, _17201_, _17197_);
  nor (_17203_, _11238_, _10453_);
  or (_17204_, _17203_, _17104_);
  and (_17205_, _17204_, _06535_);
  or (_17206_, _17205_, _06559_);
  or (_17207_, _17206_, _17202_);
  or (_17208_, _17116_, _07240_);
  and (_17209_, _17208_, _05933_);
  and (_17210_, _17209_, _17207_);
  and (_17211_, _17113_, _05932_);
  or (_17212_, _17211_, _06566_);
  or (_17213_, _17212_, _17210_);
  and (_17214_, _15695_, _07933_);
  or (_17215_, _17104_, _06570_);
  or (_17216_, _17215_, _17214_);
  and (_17217_, _17216_, _01320_);
  and (_17218_, _17217_, _17213_);
  or (_17219_, _17218_, _17103_);
  and (_42897_, _17219_, _42355_);
  nor (_17220_, _01320_, _06018_);
  and (_17221_, _11320_, \oc8051_golden_model_1.ACC [1]);
  nand (_17222_, _10472_, _08737_);
  nand (_17223_, _12533_, _06292_);
  and (_17224_, _17223_, _10475_);
  and (_17225_, _06702_, _05993_);
  nand (_17226_, _11111_, _10774_);
  nand (_17227_, _11006_, _12551_);
  and (_17228_, _06414_, _06007_);
  not (_17229_, _17228_);
  not (_17230_, _10955_);
  and (_17231_, _17230_, _11164_);
  or (_17232_, _06248_, _05985_);
  nor (_17233_, _07930_, _06018_);
  and (_17234_, _14413_, _07930_);
  or (_17235_, _17234_, _17233_);
  and (_17236_, _17235_, _05972_);
  and (_17237_, _07930_, _07135_);
  or (_17238_, _17237_, _17233_);
  or (_17239_, _17238_, _06260_);
  nor (_17240_, _10603_, _06018_);
  or (_17241_, _17240_, _10604_);
  or (_17242_, _17241_, _10555_);
  or (_17243_, _10623_, _07135_);
  nor (_17244_, _10633_, _07159_);
  or (_17245_, _17244_, _09384_);
  and (_17246_, _10645_, _07135_);
  nor (_17247_, _06755_, _06018_);
  and (_17248_, _06755_, _06018_);
  nor (_17249_, _17248_, _17247_);
  nor (_17250_, _17249_, _10645_);
  or (_17251_, _17250_, _10633_);
  or (_17252_, _17251_, _17246_);
  and (_17253_, _17252_, _05960_);
  or (_17254_, _17253_, _07159_);
  and (_17255_, _17254_, _06286_);
  and (_17256_, _17255_, _17245_);
  not (_17257_, _07930_);
  nor (_17258_, _08374_, _17257_);
  or (_17259_, _17258_, _17233_);
  and (_17260_, _17259_, _06285_);
  or (_17261_, _17260_, _06281_);
  or (_17262_, _17261_, _17256_);
  and (_17263_, _14326_, _08596_);
  nor (_17264_, _08596_, _06018_);
  or (_17265_, _17264_, _06282_);
  or (_17266_, _17265_, _17263_);
  and (_17267_, _17266_, _07169_);
  and (_17268_, _17267_, _17262_);
  and (_17269_, _17238_, _06354_);
  or (_17270_, _17269_, _10622_);
  or (_17271_, _17270_, _17268_);
  and (_17272_, _17271_, _17243_);
  or (_17273_, _17272_, _07174_);
  or (_17274_, _09384_, _10692_);
  and (_17275_, _17274_, _06346_);
  and (_17276_, _17275_, _17273_);
  and (_17277_, _08374_, _06345_);
  or (_17278_, _17277_, _10696_);
  or (_17279_, _17278_, _17276_);
  nand (_17280_, _10696_, _10123_);
  and (_17281_, _17280_, _17279_);
  or (_17282_, _17281_, _06277_);
  or (_17283_, _17233_, _06278_);
  and (_17284_, _17283_, _06271_);
  and (_17285_, _17284_, _17282_);
  and (_17286_, _17259_, _06270_);
  or (_17287_, _17286_, _09520_);
  or (_17288_, _17287_, _17285_);
  or (_17289_, _16473_, _10059_);
  and (_17290_, _17289_, _10719_);
  and (_17291_, _17290_, _10723_);
  and (_17292_, _17291_, _17288_);
  not (_17293_, _10724_);
  nor (_17294_, _10776_, _06018_);
  or (_17295_, _17294_, _10777_);
  and (_17296_, _17295_, _17293_);
  or (_17297_, _17296_, _10727_);
  or (_17298_, _17297_, _17292_);
  and (_17299_, _17298_, _17242_);
  or (_17300_, _17299_, _06380_);
  nor (_17301_, _10535_, _06018_);
  or (_17302_, _17301_, _10536_);
  or (_17303_, _17302_, _06386_);
  and (_17304_, _17303_, _10487_);
  and (_17305_, _17304_, _17300_);
  nor (_17306_, _10842_, _06018_);
  or (_17307_, _17306_, _10843_);
  and (_17308_, _17307_, _10486_);
  or (_17309_, _17308_, _05976_);
  or (_17310_, _17309_, _17305_);
  or (_17311_, _06248_, _05940_);
  and (_17312_, _17311_, _06267_);
  and (_17313_, _17312_, _17310_);
  and (_17314_, _14358_, _08596_);
  or (_17315_, _17314_, _17264_);
  and (_17316_, _17315_, _06266_);
  or (_17317_, _17316_, _06259_);
  or (_17318_, _17317_, _17313_);
  and (_17319_, _17318_, _17239_);
  or (_17320_, _17319_, _09486_);
  and (_17321_, _09384_, _07930_);
  or (_17322_, _17233_, _06258_);
  or (_17323_, _17322_, _17321_);
  and (_17324_, _17323_, _06251_);
  and (_17325_, _17324_, _17320_);
  or (_17326_, _17325_, _17236_);
  and (_17327_, _17326_, _09481_);
  or (_17328_, _17051_, _05984_);
  or (_17329_, _17328_, _17327_);
  and (_17330_, _17329_, _17232_);
  or (_17331_, _17330_, _06215_);
  and (_17332_, _07930_, _08929_);
  or (_17333_, _17332_, _17233_);
  or (_17334_, _17333_, _06216_);
  and (_17335_, _17334_, _10892_);
  and (_17336_, _17335_, _17331_);
  and (_17337_, _10891_, _06248_);
  or (_17338_, _17337_, _10899_);
  or (_17339_, _17338_, _17336_);
  and (_17340_, _07157_, _06018_);
  nor (_17341_, _17340_, _11164_);
  or (_17342_, _10905_, _17341_);
  and (_17343_, _17342_, _10909_);
  and (_17345_, _17343_, _17339_);
  and (_17346_, _10908_, _17341_);
  or (_17347_, _17346_, _10913_);
  or (_17348_, _17347_, _17345_);
  or (_17349_, _10919_, _17341_);
  and (_17350_, _17349_, _10918_);
  and (_17351_, _17350_, _17348_);
  nor (_17352_, _09384_, \oc8051_golden_model_1.ACC [0]);
  nor (_17353_, _17352_, _11217_);
  and (_17354_, _17353_, _10917_);
  or (_17356_, _17354_, _06526_);
  or (_17357_, _17356_, _17351_);
  nand (_17358_, _12533_, _06526_);
  and (_17359_, _17358_, _17357_);
  and (_17360_, _17359_, _10935_);
  and (_17361_, _10481_, _12552_);
  or (_17362_, _17361_, _06398_);
  or (_17363_, _17362_, _17360_);
  and (_17364_, _14311_, _07930_);
  or (_17365_, _17364_, _17233_);
  or (_17367_, _17365_, _09025_);
  and (_17368_, _17367_, _09030_);
  and (_17369_, _17368_, _17363_);
  and (_17370_, _17233_, _06524_);
  or (_17371_, _17370_, _10944_);
  or (_17372_, _17371_, _17369_);
  or (_17373_, _11164_, _10948_);
  and (_17374_, _17373_, _10955_);
  and (_17375_, _17374_, _17372_);
  or (_17376_, _17375_, _17231_);
  and (_17378_, _17376_, _10951_);
  and (_17379_, _11164_, _10950_);
  or (_17380_, _17379_, _17378_);
  and (_17381_, _17380_, _10964_);
  and (_17382_, _10959_, _11217_);
  or (_17383_, _17382_, _06530_);
  or (_17384_, _17383_, _17381_);
  or (_17385_, _11254_, _06531_);
  and (_17386_, _17385_, _10974_);
  and (_17387_, _17386_, _17384_);
  and (_17389_, _10968_, _11293_);
  or (_17390_, _17389_, _17387_);
  and (_17391_, _17390_, _07219_);
  nand (_17392_, _17333_, _06426_);
  nor (_17393_, _17392_, _17258_);
  and (_17394_, _05887_, _06007_);
  or (_17395_, _17394_, _17393_);
  or (_17396_, _17395_, _17391_);
  nor (_17397_, _17394_, _07060_);
  nor (_17398_, _17340_, _07060_);
  or (_17400_, _17398_, _17397_);
  and (_17401_, _17400_, _17396_);
  nor (_17402_, _17340_, _07061_);
  or (_17403_, _17402_, _17401_);
  and (_17404_, _17403_, _17229_);
  nor (_17405_, _17340_, _17229_);
  or (_17406_, _17405_, _11000_);
  or (_17407_, _17406_, _17404_);
  nand (_17408_, _11000_, _17352_);
  and (_17409_, _17408_, _06538_);
  and (_17410_, _17409_, _17407_);
  nand (_17411_, _11009_, _12532_);
  and (_17412_, _17411_, _11008_);
  or (_17413_, _17412_, _17410_);
  and (_17414_, _17413_, _17227_);
  or (_17415_, _17414_, _06437_);
  and (_17416_, _14307_, _07930_);
  or (_17417_, _17233_, _07229_);
  or (_17418_, _17417_, _17416_);
  and (_17419_, _17418_, _11023_);
  and (_17420_, _17419_, _17415_);
  and (_17421_, _11024_, _17295_);
  or (_17422_, _17421_, _13990_);
  or (_17423_, _17422_, _17420_);
  or (_17424_, _11027_, _17241_);
  and (_17425_, _17424_, _17423_);
  or (_17426_, _17425_, _06522_);
  or (_17427_, _17302_, _06523_);
  and (_17428_, _17427_, _11083_);
  and (_17429_, _17428_, _17426_);
  and (_17430_, _11082_, _17307_);
  or (_17431_, _17430_, _11111_);
  or (_17432_, _17431_, _17429_);
  and (_17433_, _17432_, _17226_);
  or (_17434_, _17433_, _17225_);
  and (_17435_, _05887_, _05993_);
  nand (_17436_, _17341_, _05926_);
  nand (_17437_, _17436_, _17435_);
  and (_17438_, _06801_, _05993_);
  and (_17439_, _10953_, _05993_);
  nor (_17440_, _17439_, _17438_);
  and (_17441_, _17440_, _17437_);
  and (_17442_, _17441_, _17434_);
  or (_17443_, _17439_, _06715_);
  or (_17444_, _17443_, _17438_);
  and (_17445_, _17444_, _17341_);
  or (_17446_, _17445_, _11189_);
  or (_17447_, _17446_, _17442_);
  not (_17448_, _11188_);
  not (_17449_, _11189_);
  or (_17450_, _17449_, _17353_);
  and (_17451_, _17450_, _17448_);
  and (_17452_, _17451_, _17447_);
  and (_17453_, _17353_, _11188_);
  or (_17454_, _17453_, _06292_);
  or (_17455_, _17454_, _17452_);
  and (_17456_, _17455_, _17224_);
  and (_17457_, _12552_, _10474_);
  or (_17458_, _17457_, _10472_);
  or (_17459_, _17458_, _17456_);
  and (_17460_, _17459_, _17222_);
  or (_17461_, _17460_, _06559_);
  or (_17462_, _17259_, _07240_);
  and (_17463_, _17462_, _11316_);
  and (_17464_, _17463_, _17461_);
  and (_17465_, _11315_, _06018_);
  or (_17466_, _17465_, _17464_);
  and (_17467_, _17466_, _14289_);
  or (_17468_, _17467_, _17221_);
  and (_17469_, _17468_, _05933_);
  and (_17470_, _17233_, _05932_);
  or (_17471_, _17470_, _06566_);
  or (_17472_, _17471_, _17469_);
  or (_17473_, _17259_, _06570_);
  and (_17474_, _17473_, _11339_);
  and (_17475_, _17474_, _17472_);
  nor (_17476_, _11345_, _06018_);
  nor (_17477_, _17476_, _13027_);
  or (_17478_, _17477_, _17475_);
  nand (_17479_, _11345_, _06044_);
  and (_17480_, _17479_, _01320_);
  and (_17481_, _17480_, _17478_);
  or (_17482_, _17481_, _17220_);
  and (_42898_, _17482_, _42355_);
  nor (_17483_, _01320_, _06044_);
  nor (_17484_, _11217_, _11216_);
  nor (_17485_, _17484_, _11218_);
  or (_17486_, _17485_, _17449_);
  or (_17487_, _11092_, _11091_);
  nor (_17488_, _11093_, _06523_);
  and (_17489_, _17488_, _17487_);
  not (_17490_, _11026_);
  nor (_17491_, _11063_, _11062_);
  nor (_17492_, _17491_, _11064_);
  or (_17493_, _17492_, _17490_);
  nor (_17494_, _11162_, _07060_);
  or (_17495_, _17494_, _17397_);
  and (_17496_, _11161_, _10950_);
  or (_17497_, _11253_, _06527_);
  nor (_17498_, _07930_, _06044_);
  and (_17499_, _07930_, _09422_);
  or (_17500_, _17499_, _17498_);
  or (_17501_, _17500_, _06260_);
  nor (_17502_, _08596_, _06044_);
  and (_17503_, _14508_, _08596_);
  or (_17504_, _17503_, _17502_);
  or (_17505_, _17502_, _14507_);
  and (_17506_, _17505_, _06270_);
  and (_17507_, _17506_, _17504_);
  or (_17508_, _10623_, _09422_);
  or (_17509_, _17244_, _09339_);
  and (_17510_, _10645_, _09422_);
  or (_17511_, _06755_, \oc8051_golden_model_1.ACC [1]);
  nand (_17512_, _06755_, \oc8051_golden_model_1.ACC [1]);
  nand (_17513_, _17512_, _17511_);
  nor (_17514_, _17513_, _10645_);
  or (_17515_, _17514_, _10633_);
  or (_17516_, _17515_, _17510_);
  and (_17517_, _17516_, _05960_);
  or (_17518_, _17517_, _07159_);
  and (_17519_, _17518_, _17509_);
  or (_17520_, _17519_, _06285_);
  or (_17521_, _07930_, \oc8051_golden_model_1.ACC [1]);
  and (_17522_, _14520_, _07930_);
  not (_17523_, _17522_);
  and (_17524_, _17523_, _17521_);
  or (_17525_, _17524_, _06286_);
  and (_17526_, _17525_, _17520_);
  or (_17527_, _17526_, _10656_);
  nor (_17528_, _10660_, \oc8051_golden_model_1.PSW [6]);
  nor (_17529_, _17528_, \oc8051_golden_model_1.ACC [1]);
  and (_17530_, _17528_, \oc8051_golden_model_1.ACC [1]);
  nor (_17531_, _17530_, _17529_);
  nand (_17532_, _17531_, _10656_);
  and (_17533_, _17532_, _06361_);
  and (_17534_, _17533_, _17527_);
  and (_17535_, _17504_, _06281_);
  and (_17536_, _17500_, _06354_);
  or (_17537_, _17536_, _10622_);
  or (_17538_, _17537_, _17535_);
  or (_17539_, _17538_, _17534_);
  and (_17540_, _17539_, _17508_);
  or (_17541_, _17540_, _07174_);
  or (_17542_, _09339_, _10692_);
  and (_17543_, _17542_, _06346_);
  and (_17544_, _17543_, _17541_);
  nor (_17545_, _08324_, _06346_);
  or (_17546_, _17545_, _10696_);
  or (_17547_, _17546_, _17544_);
  nand (_17548_, _10696_, _10152_);
  and (_17549_, _17548_, _17547_);
  or (_17550_, _17549_, _06277_);
  and (_17551_, _14511_, _08596_);
  or (_17552_, _17551_, _17502_);
  or (_17553_, _17552_, _06278_);
  and (_17554_, _17553_, _06271_);
  and (_17555_, _17554_, _17550_);
  or (_17556_, _17555_, _17507_);
  and (_17557_, _17556_, _10059_);
  nor (_17558_, _10007_, _10006_);
  nor (_17559_, _17558_, _10008_);
  nand (_17560_, _17559_, _09520_);
  nand (_17561_, _17560_, _10724_);
  or (_17562_, _17561_, _17557_);
  nor (_17563_, _10769_, _06018_);
  or (_17564_, _17563_, _10775_);
  and (_17565_, _17564_, _11163_);
  nor (_17566_, _17564_, _11163_);
  or (_17567_, _17566_, _17565_);
  or (_17568_, _17567_, _10724_);
  and (_17569_, _17568_, _10555_);
  and (_17570_, _17569_, _17562_);
  not (_17571_, _11216_);
  nor (_17572_, _10556_, _06018_);
  or (_17573_, _17572_, _10602_);
  nand (_17574_, _17573_, _17571_);
  or (_17575_, _17573_, _17571_);
  and (_17576_, _17575_, _10727_);
  and (_17577_, _17576_, _17574_);
  or (_17578_, _17577_, _06380_);
  or (_17579_, _17578_, _17570_);
  nor (_17580_, _10488_, _06018_);
  or (_17581_, _17580_, _10534_);
  nor (_17582_, _17581_, _11253_);
  and (_17583_, _17581_, _11253_);
  or (_17584_, _17583_, _06386_);
  or (_17585_, _17584_, _17582_);
  and (_17586_, _17585_, _10487_);
  and (_17587_, _17586_, _17579_);
  nor (_17588_, _08786_, _06018_);
  nor (_17589_, _17588_, _10841_);
  or (_17590_, _17589_, _11292_);
  nand (_17591_, _17589_, _11292_);
  and (_17592_, _17591_, _10486_);
  and (_17593_, _17592_, _17590_);
  or (_17594_, _17593_, _05976_);
  or (_17595_, _17594_, _17587_);
  nand (_17596_, _06995_, _05976_);
  and (_17597_, _17596_, _06267_);
  and (_17598_, _17597_, _17595_);
  or (_17599_, _17502_, _14551_);
  and (_17600_, _17599_, _06266_);
  and (_17601_, _17600_, _17504_);
  or (_17602_, _17601_, _06259_);
  or (_17603_, _17602_, _17598_);
  and (_17604_, _17603_, _17501_);
  or (_17605_, _17604_, _09486_);
  and (_17606_, _09339_, _07930_);
  or (_17607_, _17498_, _06258_);
  or (_17608_, _17607_, _17606_);
  and (_17609_, _17608_, _06251_);
  and (_17610_, _17609_, _17605_);
  or (_17611_, _14607_, _17257_);
  and (_17612_, _17521_, _05972_);
  and (_17613_, _17612_, _17611_);
  or (_17614_, _17613_, _09480_);
  or (_17615_, _17614_, _17610_);
  nand (_17616_, _10330_, _09480_);
  and (_17617_, _17616_, _17615_);
  or (_17618_, _17617_, _05984_);
  nand (_17619_, _06995_, _05984_);
  and (_17620_, _17619_, _06216_);
  and (_17621_, _17620_, _17618_);
  nand (_17622_, _07930_, _07031_);
  and (_17623_, _17622_, _06215_);
  and (_17624_, _17623_, _17521_);
  or (_17625_, _17624_, _10891_);
  or (_17626_, _17625_, _17621_);
  nand (_17627_, _10891_, _06995_);
  and (_17628_, _17627_, _10905_);
  and (_17629_, _17628_, _17626_);
  and (_17630_, _10899_, _11163_);
  or (_17631_, _17630_, _17629_);
  and (_17632_, _17631_, _12693_);
  not (_17633_, _12693_);
  and (_17634_, _17633_, _11163_);
  or (_17635_, _17634_, _06866_);
  or (_17636_, _17635_, _17632_);
  or (_17637_, _11163_, _06867_);
  and (_17638_, _17637_, _10918_);
  and (_17639_, _17638_, _17636_);
  and (_17640_, _11216_, _10917_);
  or (_17641_, _17640_, _06526_);
  or (_17642_, _17641_, _17639_);
  and (_17643_, _17642_, _17497_);
  or (_17644_, _17643_, _10481_);
  or (_17645_, _10935_, _11292_);
  and (_17646_, _17645_, _09025_);
  and (_17647_, _17646_, _17644_);
  or (_17648_, _14505_, _17257_);
  and (_17649_, _17521_, _06398_);
  and (_17650_, _17649_, _17648_);
  or (_17651_, _17650_, _17647_);
  and (_17652_, _17651_, _09030_);
  nand (_17653_, _17498_, _06524_);
  and (_17654_, _07466_, _06012_);
  not (_17655_, _17654_);
  and (_17656_, _09006_, _06012_);
  or (_17657_, _17656_, _07065_);
  nor (_17658_, _07472_, _06875_);
  nor (_17659_, _17658_, _17657_);
  and (_17660_, _17659_, _17655_);
  nand (_17661_, _17660_, _17653_);
  or (_17662_, _17661_, _17652_);
  or (_17663_, _17660_, _11161_);
  and (_17664_, _17663_, _10951_);
  and (_17665_, _17664_, _17662_);
  or (_17666_, _17665_, _17496_);
  and (_17667_, _17666_, _10964_);
  and (_17668_, _10959_, _11213_);
  or (_17669_, _17668_, _06530_);
  or (_17670_, _17669_, _17667_);
  or (_17671_, _11251_, _06531_);
  and (_17672_, _17671_, _10974_);
  and (_17673_, _17672_, _17670_);
  and (_17674_, _10968_, _11290_);
  or (_17675_, _17674_, _17673_);
  and (_17676_, _17675_, _07219_);
  or (_17677_, _14503_, _17257_);
  and (_17678_, _17521_, _06426_);
  and (_17679_, _17678_, _17677_);
  or (_17680_, _17679_, _17394_);
  or (_17681_, _17680_, _17676_);
  and (_17682_, _17681_, _17495_);
  nor (_17683_, _11162_, _07061_);
  or (_17684_, _17683_, _17682_);
  and (_17685_, _17684_, _17229_);
  nor (_17686_, _11162_, _17229_);
  or (_17687_, _17686_, _11000_);
  or (_17688_, _17687_, _17685_);
  not (_17689_, _11000_);
  or (_17690_, _17689_, _11215_);
  and (_17691_, _17690_, _06538_);
  and (_17692_, _17691_, _17688_);
  nand (_17693_, _11009_, _11252_);
  and (_17694_, _17693_, _11008_);
  or (_17695_, _17694_, _17692_);
  nand (_17696_, _11006_, _11291_);
  and (_17697_, _17696_, _07229_);
  and (_17698_, _17697_, _17695_);
  or (_17699_, _17622_, _08325_);
  and (_17700_, _17699_, _06437_);
  and (_17701_, _17700_, _17521_);
  or (_17702_, _17701_, _11017_);
  or (_17703_, _17702_, _17698_);
  nor (_17704_, _11036_, _11035_);
  nor (_17705_, _17704_, _11037_);
  or (_17706_, _17705_, _11018_);
  nand (_17707_, _17706_, _17703_);
  nand (_17708_, _17707_, _11021_);
  or (_17709_, _17705_, _11021_);
  and (_17710_, _17709_, _11020_);
  and (_17711_, _17710_, _17708_);
  and (_17712_, _17705_, _11019_);
  or (_17713_, _17712_, _11026_);
  or (_17714_, _17713_, _17711_);
  and (_17715_, _17714_, _17493_);
  or (_17716_, _17715_, _06892_);
  not (_17717_, _06892_);
  or (_17718_, _17492_, _17717_);
  and (_17719_, _17718_, _06523_);
  and (_17720_, _17719_, _17716_);
  or (_17721_, _17720_, _17489_);
  and (_17722_, _17721_, _11083_);
  or (_17723_, _11120_, _11119_);
  nor (_17724_, _11121_, _11083_);
  and (_17725_, _17724_, _17723_);
  or (_17726_, _17725_, _11111_);
  or (_17727_, _17726_, _17722_);
  nand (_17728_, _11111_, _06018_);
  and (_17729_, _17728_, _11185_);
  and (_17730_, _17729_, _17727_);
  or (_17731_, _11164_, _11163_);
  nor (_17732_, _11185_, _11165_);
  and (_17733_, _17732_, _17731_);
  or (_17734_, _17733_, _11189_);
  or (_17735_, _17734_, _17730_);
  and (_17736_, _17735_, _17486_);
  or (_17737_, _17736_, _11188_);
  or (_17738_, _17485_, _17448_);
  and (_17739_, _17738_, _06293_);
  and (_17740_, _17739_, _17737_);
  nor (_17741_, _11254_, _11253_);
  nor (_17742_, _17741_, _11255_);
  or (_17743_, _17742_, _10474_);
  and (_17744_, _17743_, _12979_);
  or (_17745_, _17744_, _17740_);
  nor (_17746_, _11293_, _11292_);
  nor (_17747_, _17746_, _11294_);
  or (_17748_, _17747_, _10475_);
  and (_17749_, _17748_, _12981_);
  and (_17750_, _17749_, _17745_);
  and (_17751_, _10472_, \oc8051_golden_model_1.ACC [0]);
  or (_17752_, _17751_, _06559_);
  or (_17753_, _17752_, _17750_);
  or (_17754_, _17524_, _07240_);
  and (_17755_, _17754_, _11316_);
  and (_17756_, _17755_, _17753_);
  nor (_17757_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor (_17758_, _11346_, _17757_);
  nor (_17759_, _17758_, _11316_);
  or (_17760_, _17759_, _11320_);
  or (_17761_, _17760_, _17756_);
  nand (_17762_, _11320_, _10198_);
  and (_17763_, _17762_, _05933_);
  and (_17764_, _17763_, _17761_);
  and (_17765_, _17552_, _05932_);
  or (_17766_, _17765_, _06566_);
  or (_17767_, _17766_, _17764_);
  or (_17768_, _17522_, _17498_);
  or (_17769_, _17768_, _06570_);
  and (_17770_, _17769_, _11339_);
  and (_17771_, _17770_, _17767_);
  and (_17772_, _17758_, _11338_);
  or (_17773_, _17772_, _11345_);
  or (_17774_, _17773_, _17771_);
  nand (_17775_, _11345_, _10198_);
  and (_17776_, _17775_, _01320_);
  and (_17777_, _17776_, _17774_);
  or (_17778_, _17777_, _17483_);
  and (_42900_, _17778_, _42355_);
  nor (_17779_, _01320_, _10198_);
  nand (_17780_, _10472_, _06044_);
  and (_17781_, _11038_, _10767_);
  nor (_17782_, _17781_, _11039_);
  and (_17783_, _17782_, _11024_);
  and (_17784_, _06414_, _06012_);
  not (_17785_, _17784_);
  nor (_17786_, _07509_, _06875_);
  and (_17787_, _17786_, _11158_);
  or (_17788_, _11211_, _10918_);
  and (_17789_, _06407_, _06000_);
  nand (_17790_, _05887_, _06000_);
  or (_17791_, _17790_, _11160_);
  nand (_17792_, _06646_, _05984_);
  nor (_17793_, _07930_, _10198_);
  and (_17794_, _07930_, _08662_);
  or (_17795_, _17794_, _17793_);
  or (_17796_, _17795_, _06260_);
  or (_17797_, _10623_, _08662_);
  or (_17798_, _17244_, _09293_);
  and (_17799_, _10645_, _08662_);
  or (_17800_, _06755_, \oc8051_golden_model_1.ACC [2]);
  nand (_17801_, _06755_, \oc8051_golden_model_1.ACC [2]);
  nand (_17802_, _17801_, _17800_);
  nor (_17803_, _17802_, _10645_);
  or (_17804_, _17803_, _10633_);
  or (_17805_, _17804_, _17799_);
  and (_17806_, _17805_, _05960_);
  or (_17807_, _17806_, _07159_);
  and (_17808_, _17807_, _17798_);
  or (_17809_, _17808_, _06285_);
  and (_17810_, _14703_, _07930_);
  or (_17811_, _17810_, _17793_);
  or (_17812_, _17811_, _06286_);
  and (_17813_, _17812_, _17809_);
  or (_17814_, _17813_, _10656_);
  nor (_17815_, _17529_, _10198_);
  and (_17816_, _10659_, \oc8051_golden_model_1.PSW [6]);
  nor (_17817_, _17816_, _17815_);
  nand (_17818_, _17817_, _10656_);
  and (_17819_, _17818_, _06361_);
  and (_17820_, _17819_, _17814_);
  nor (_17821_, _08596_, _10198_);
  and (_17822_, _14716_, _08596_);
  or (_17823_, _17822_, _17821_);
  and (_17824_, _17823_, _06281_);
  and (_17825_, _17795_, _06354_);
  or (_17826_, _17825_, _10622_);
  or (_17827_, _17826_, _17824_);
  or (_17828_, _17827_, _17820_);
  and (_17829_, _17828_, _17797_);
  or (_17830_, _17829_, _07174_);
  or (_17831_, _09293_, _10692_);
  and (_17832_, _17831_, _06346_);
  and (_17833_, _17832_, _17830_);
  nor (_17834_, _08423_, _06346_);
  or (_17835_, _17834_, _10696_);
  or (_17836_, _17835_, _17833_);
  nand (_17837_, _10696_, _10105_);
  and (_17838_, _17837_, _17836_);
  or (_17839_, _17838_, _06277_);
  and (_17840_, _14699_, _08596_);
  or (_17841_, _17840_, _17821_);
  or (_17842_, _17841_, _06278_);
  and (_17843_, _17842_, _06271_);
  and (_17844_, _17843_, _17839_);
  or (_17845_, _17821_, _14731_);
  and (_17846_, _17823_, _06270_);
  and (_17847_, _17846_, _17845_);
  or (_17848_, _17847_, _09520_);
  or (_17849_, _17848_, _17844_);
  nor (_17850_, _10010_, _10008_);
  or (_17851_, _17850_, _10011_);
  nand (_17852_, _17851_, _09520_);
  and (_17853_, _17852_, _10724_);
  and (_17854_, _17853_, _17849_);
  and (_17855_, _07334_, \oc8051_golden_model_1.ACC [1]);
  and (_17856_, _07135_, _06018_);
  nor (_17857_, _17856_, _11163_);
  nor (_17858_, _17857_, _17855_);
  nor (_17859_, _11160_, _17858_);
  and (_17860_, _11160_, _17858_);
  nor (_17861_, _17860_, _17859_);
  nor (_17862_, _17341_, _11163_);
  and (_17863_, _17862_, \oc8051_golden_model_1.PSW [7]);
  or (_17864_, _17863_, _17861_);
  nand (_17865_, _17863_, _17861_);
  and (_17866_, _17865_, _17293_);
  and (_17867_, _17866_, _17864_);
  or (_17868_, _17867_, _10727_);
  or (_17869_, _17868_, _17854_);
  or (_17870_, _09339_, _06044_);
  and (_17871_, _09384_, _06018_);
  or (_17872_, _17871_, _11216_);
  and (_17873_, _17872_, _17870_);
  nor (_17874_, _11211_, _17873_);
  and (_17875_, _11211_, _17873_);
  or (_17876_, _17875_, _17874_);
  nor (_17877_, _17353_, _11216_);
  and (_17878_, _17877_, \oc8051_golden_model_1.PSW [7]);
  nor (_17879_, _17878_, _17876_);
  and (_17880_, _17878_, _17876_);
  or (_17881_, _17880_, _10555_);
  or (_17882_, _17881_, _17879_);
  and (_17883_, _17882_, _17869_);
  or (_17884_, _17883_, _06380_);
  and (_17885_, _08324_, \oc8051_golden_model_1.ACC [1]);
  and (_17886_, _08374_, _06018_);
  nor (_17887_, _14097_, _17886_);
  nor (_17888_, _17887_, _17885_);
  nor (_17889_, _11250_, _17888_);
  and (_17890_, _11250_, _17888_);
  nor (_17891_, _17890_, _17889_);
  and (_17892_, _12534_, \oc8051_golden_model_1.PSW [7]);
  or (_17893_, _17892_, _17891_);
  nand (_17894_, _17892_, _17891_);
  and (_17895_, _17894_, _17893_);
  or (_17896_, _17895_, _06386_);
  and (_17897_, _17896_, _10487_);
  and (_17898_, _17897_, _17884_);
  and (_17899_, _06248_, _06018_);
  nor (_17900_, _17899_, _11292_);
  nor (_17901_, _17900_, _14109_);
  not (_17902_, _11289_);
  nor (_17903_, _17902_, _17901_);
  and (_17904_, _17902_, _17901_);
  nor (_17905_, _17904_, _17903_);
  and (_17906_, _12553_, \oc8051_golden_model_1.PSW [7]);
  not (_17907_, _17906_);
  or (_17908_, _17907_, _17905_);
  nand (_17909_, _17907_, _17905_);
  nand (_17910_, _17909_, _17908_);
  and (_17911_, _17910_, _10486_);
  or (_17912_, _17911_, _05976_);
  or (_17913_, _17912_, _17898_);
  nand (_17914_, _06646_, _05976_);
  and (_17915_, _17914_, _06267_);
  and (_17916_, _17915_, _17913_);
  and (_17917_, _14749_, _08596_);
  or (_17918_, _17917_, _17821_);
  and (_17919_, _17918_, _06266_);
  or (_17920_, _17919_, _06259_);
  or (_17921_, _17920_, _17916_);
  and (_17922_, _17921_, _17796_);
  or (_17923_, _17922_, _09486_);
  and (_17924_, _09293_, _07930_);
  or (_17925_, _17793_, _06258_);
  or (_17926_, _17925_, _17924_);
  and (_17927_, _17926_, _06251_);
  and (_17928_, _17927_, _17923_);
  and (_17929_, _14804_, _07930_);
  or (_17930_, _17929_, _17793_);
  and (_17931_, _17930_, _05972_);
  or (_17932_, _17931_, _09480_);
  or (_17933_, _17932_, _17928_);
  or (_17934_, _10266_, _09481_);
  and (_17935_, _17934_, _17933_);
  or (_17936_, _17935_, _05984_);
  and (_17937_, _17936_, _17792_);
  or (_17938_, _17937_, _06215_);
  and (_17939_, _07930_, _08980_);
  or (_17940_, _17939_, _17793_);
  or (_17941_, _17940_, _06216_);
  and (_17942_, _17941_, _10892_);
  and (_17943_, _17942_, _17938_);
  or (_17944_, _10892_, _06646_);
  nand (_17945_, _17944_, _17790_);
  or (_17946_, _17945_, _17943_);
  and (_17947_, _17946_, _17791_);
  or (_17948_, _17947_, _17789_);
  not (_17949_, _17789_);
  or (_17950_, _11160_, _17949_);
  and (_17951_, _05882_, _05934_);
  and (_17952_, _17951_, _06000_);
  not (_17953_, _17952_);
  and (_17954_, _17953_, _17950_);
  and (_17955_, _17954_, _17948_);
  and (_17956_, _17952_, _11160_);
  or (_17957_, _17956_, _10917_);
  or (_17958_, _17957_, _17955_);
  and (_17959_, _17958_, _17788_);
  or (_17960_, _17959_, _06526_);
  or (_17961_, _11250_, _06527_);
  and (_17962_, _17961_, _10935_);
  and (_17963_, _17962_, _17960_);
  nor (_17964_, _10935_, _11289_);
  or (_17965_, _17964_, _06398_);
  or (_17966_, _17965_, _17963_);
  and (_17967_, _14697_, _07930_);
  or (_17969_, _17967_, _17793_);
  or (_17970_, _17969_, _09025_);
  and (_17971_, _17970_, _17966_);
  or (_17972_, _17971_, _06524_);
  not (_17973_, _17786_);
  or (_17974_, _17793_, _09030_);
  and (_17975_, _17974_, _17973_);
  and (_17976_, _17975_, _17972_);
  or (_17977_, _17976_, _17787_);
  and (_17978_, _17977_, _17785_);
  and (_17979_, _11158_, _17784_);
  or (_17980_, _17979_, _17978_);
  and (_17981_, _17980_, _10964_);
  and (_17982_, _10959_, _11208_);
  or (_17983_, _17982_, _06530_);
  or (_17984_, _17983_, _17981_);
  or (_17985_, _11248_, _06531_);
  and (_17986_, _17985_, _10974_);
  and (_17987_, _17986_, _17984_);
  and (_17988_, _10968_, _11286_);
  or (_17989_, _17988_, _17987_);
  and (_17990_, _17989_, _07219_);
  nand (_17991_, _17940_, _06426_);
  nor (_17992_, _17991_, _11249_);
  or (_17993_, _17992_, _17990_);
  and (_17994_, _17993_, _10987_);
  nor (_17995_, _10987_, _11159_);
  or (_17996_, _17995_, _10991_);
  or (_17997_, _17996_, _17994_);
  nand (_17998_, _10991_, _11159_);
  and (_17999_, _17998_, _10995_);
  and (_18000_, _17999_, _17997_);
  nor (_18001_, _11159_, _10995_);
  or (_18002_, _18001_, _11000_);
  or (_18003_, _18002_, _18000_);
  or (_18004_, _17689_, _11210_);
  and (_18005_, _18004_, _06538_);
  and (_18006_, _18005_, _18003_);
  nand (_18007_, _11009_, _11249_);
  and (_18008_, _18007_, _11008_);
  or (_18009_, _18008_, _18006_);
  nand (_18010_, _06646_, _10198_);
  or (_18011_, _11009_, _18010_);
  and (_18012_, _18011_, _18009_);
  or (_18013_, _18012_, _06437_);
  and (_18014_, _14694_, _07930_);
  or (_18015_, _17793_, _07229_);
  or (_18016_, _18015_, _18014_);
  and (_18017_, _18016_, _11023_);
  and (_18018_, _18017_, _18013_);
  or (_18019_, _18018_, _17783_);
  and (_18020_, _18019_, _17490_);
  and (_18021_, _11065_, _10596_);
  nor (_18022_, _18021_, _11066_);
  and (_18023_, _18022_, _11026_);
  or (_18024_, _18023_, _06892_);
  or (_18025_, _18024_, _18020_);
  or (_18026_, _18022_, _17717_);
  and (_18027_, _18026_, _06523_);
  and (_18028_, _18027_, _18025_);
  and (_18029_, _11094_, _10528_);
  nor (_18030_, _18029_, _11095_);
  and (_18031_, _18030_, _06522_);
  or (_18032_, _18031_, _11082_);
  or (_18033_, _18032_, _18028_);
  and (_18034_, _11122_, _10835_);
  nor (_18035_, _18034_, _11123_);
  or (_18036_, _18035_, _11083_);
  and (_18037_, _18036_, _18033_);
  or (_18038_, _18037_, _11111_);
  nand (_18039_, _11111_, _06044_);
  and (_18040_, _18039_, _11185_);
  and (_18041_, _18040_, _18038_);
  or (_18042_, _11167_, _11160_);
  nor (_18043_, _11185_, _11168_);
  and (_18044_, _18043_, _18042_);
  or (_18045_, _18044_, _11189_);
  or (_18046_, _18045_, _18041_);
  and (_18047_, _11219_, _11212_);
  nor (_18048_, _18047_, _11220_);
  and (_18049_, _18048_, _17448_);
  or (_18050_, _18049_, _11190_);
  and (_18051_, _18050_, _18046_);
  and (_18052_, _18048_, _11188_);
  or (_18053_, _18052_, _06292_);
  or (_18054_, _18053_, _18051_);
  nor (_18055_, _11257_, _11250_);
  nor (_18056_, _18055_, _11258_);
  or (_18057_, _18056_, _06293_);
  and (_18058_, _18057_, _10475_);
  and (_18059_, _18058_, _18054_);
  nand (_18060_, _11295_, _11289_);
  nor (_18061_, _11296_, _10475_);
  and (_18062_, _18061_, _18060_);
  or (_18063_, _18062_, _10472_);
  or (_18064_, _18063_, _18059_);
  and (_18065_, _18064_, _17780_);
  or (_18066_, _18065_, _06559_);
  or (_18067_, _17811_, _07240_);
  and (_18068_, _18067_, _11316_);
  and (_18069_, _18068_, _18066_);
  nor (_18070_, _17757_, _10198_);
  or (_18071_, _18070_, _11321_);
  and (_18072_, _18071_, _11315_);
  or (_18073_, _18072_, _11320_);
  or (_18074_, _18073_, _18069_);
  nand (_18075_, _11320_, _10248_);
  and (_18076_, _18075_, _05933_);
  and (_18077_, _18076_, _18074_);
  and (_18078_, _17841_, _05932_);
  or (_18079_, _18078_, _06566_);
  or (_18080_, _18079_, _18077_);
  and (_18081_, _14873_, _07930_);
  or (_18082_, _18081_, _17793_);
  or (_18083_, _18082_, _06570_);
  and (_18084_, _18083_, _11339_);
  and (_18085_, _18084_, _18080_);
  nor (_18086_, _11346_, \oc8051_golden_model_1.ACC [2]);
  nor (_18087_, _18086_, _11347_);
  and (_18088_, _18087_, _11338_);
  or (_18089_, _18088_, _11345_);
  or (_18090_, _18089_, _18085_);
  nand (_18091_, _11345_, _10248_);
  and (_18092_, _18091_, _01320_);
  and (_18093_, _18092_, _18090_);
  or (_18094_, _18093_, _17779_);
  and (_42901_, _18094_, _42355_);
  nor (_18095_, _01320_, _10248_);
  and (_18096_, _11040_, _10761_);
  nor (_18097_, _18096_, _11041_);
  or (_18098_, _18097_, _11023_);
  nor (_18099_, _11157_, _07060_);
  or (_18100_, _18099_, _17397_);
  and (_18101_, _17786_, _11156_);
  or (_18102_, _12529_, _06527_);
  and (_18103_, _18102_, _10935_);
  nand (_18104_, _06212_, _05984_);
  nor (_18105_, _07930_, _10248_);
  and (_18106_, _07930_, _09421_);
  or (_18107_, _18106_, _18105_);
  or (_18108_, _18107_, _06260_);
  and (_18109_, _07760_, \oc8051_golden_model_1.ACC [2]);
  nor (_18110_, _17859_, _18109_);
  nor (_18111_, _11157_, _11156_);
  nor (_18112_, _18111_, _18110_);
  and (_18113_, _18111_, _18110_);
  nor (_18114_, _18113_, _18112_);
  and (_18115_, _18114_, \oc8051_golden_model_1.PSW [7]);
  nor (_18116_, _18114_, \oc8051_golden_model_1.PSW [7]);
  nor (_18117_, _18116_, _18115_);
  not (_18118_, _18117_);
  and (_18119_, _17861_, \oc8051_golden_model_1.PSW [7]);
  nor (_18120_, _17862_, _10774_);
  nor (_18121_, _18120_, _18119_);
  nor (_18122_, _18121_, _18118_);
  and (_18123_, _18121_, _18118_);
  or (_18124_, _18123_, _18122_);
  nand (_18125_, _18124_, _17293_);
  nor (_18126_, _08596_, _10248_);
  and (_18127_, _14897_, _08596_);
  or (_18128_, _18127_, _18126_);
  or (_18129_, _18126_, _14926_);
  and (_18130_, _18129_, _06270_);
  and (_18131_, _18130_, _18128_);
  or (_18132_, _10623_, _09421_);
  or (_18133_, _18128_, _06282_);
  and (_18134_, _18133_, _07169_);
  and (_18135_, _14900_, _07930_);
  or (_18136_, _18135_, _18105_);
  and (_18137_, _18136_, _06285_);
  not (_18138_, _10645_);
  or (_18139_, _18138_, _09421_);
  or (_18140_, _06755_, \oc8051_golden_model_1.ACC [3]);
  nand (_18141_, _06755_, \oc8051_golden_model_1.ACC [3]);
  and (_18142_, _18141_, _18140_);
  or (_18143_, _18142_, _10645_);
  and (_18144_, _18143_, _10634_);
  and (_18145_, _18144_, _18139_);
  and (_18146_, _18145_, _08639_);
  or (_18147_, _18146_, _09247_);
  or (_18148_, _18145_, _10633_);
  and (_18149_, _18148_, _05960_);
  or (_18150_, _18149_, _07159_);
  and (_18151_, _18150_, _06286_);
  and (_18152_, _18151_, _18147_);
  or (_18153_, _18152_, _18137_);
  and (_18154_, _18153_, _10657_);
  not (_18155_, \oc8051_golden_model_1.PSW [6]);
  nor (_18156_, _10659_, _18155_);
  nor (_18157_, _18156_, \oc8051_golden_model_1.ACC [3]);
  nor (_18158_, _18157_, _10660_);
  and (_18159_, _18158_, _10656_);
  or (_18160_, _18159_, _06281_);
  or (_18161_, _18160_, _18154_);
  and (_18162_, _18161_, _18134_);
  and (_18163_, _18107_, _06354_);
  or (_18164_, _18163_, _10622_);
  or (_18165_, _18164_, _18162_);
  and (_18166_, _18165_, _18132_);
  or (_18167_, _18166_, _07174_);
  or (_18168_, _09247_, _10692_);
  and (_18169_, _18168_, _06346_);
  and (_18170_, _18169_, _18167_);
  nor (_18171_, _08279_, _06346_);
  or (_18172_, _18171_, _10696_);
  or (_18173_, _18172_, _18170_);
  nand (_18174_, _10696_, _08737_);
  and (_18175_, _18174_, _18173_);
  or (_18176_, _18175_, _06277_);
  and (_18177_, _14895_, _08596_);
  or (_18178_, _18177_, _18126_);
  or (_18179_, _18178_, _06278_);
  and (_18180_, _18179_, _06271_);
  and (_18181_, _18180_, _18176_);
  or (_18182_, _18181_, _18131_);
  and (_18183_, _18182_, _10059_);
  or (_18184_, _10013_, _10011_);
  nor (_18185_, _10014_, _10059_);
  nand (_18186_, _18185_, _18184_);
  nand (_18187_, _18186_, _10724_);
  or (_18188_, _18187_, _18183_);
  and (_18189_, _18188_, _18125_);
  or (_18190_, _18189_, _10727_);
  nand (_18191_, _17877_, _17876_);
  and (_18192_, _18191_, \oc8051_golden_model_1.PSW [7]);
  nor (_18193_, _09293_, _10198_);
  nor (_18194_, _17874_, _18193_);
  nor (_18195_, _11207_, _11206_);
  not (_18196_, _18195_);
  nand (_18197_, _18196_, _18194_);
  or (_18198_, _18196_, _18194_);
  and (_18199_, _18198_, _18197_);
  or (_18200_, _18199_, _10774_);
  nand (_18201_, _18199_, _10774_);
  and (_18202_, _18201_, _18200_);
  nand (_18203_, _18202_, _18192_);
  or (_18204_, _18202_, _18192_);
  and (_18205_, _18204_, _18203_);
  or (_18206_, _18205_, _10555_);
  and (_18207_, _18206_, _06386_);
  and (_18208_, _18207_, _18190_);
  and (_18209_, _12535_, \oc8051_golden_model_1.PSW [7]);
  and (_18210_, _08423_, \oc8051_golden_model_1.ACC [2]);
  nor (_18211_, _17889_, _18210_);
  nor (_18212_, _12529_, _18211_);
  and (_18213_, _12529_, _18211_);
  nor (_18214_, _18213_, _18212_);
  not (_18215_, _12534_);
  or (_18216_, _18215_, _17891_);
  or (_18217_, _18216_, _10774_);
  and (_18218_, _18217_, _18214_);
  or (_18219_, _18218_, _10486_);
  or (_18220_, _18219_, _18209_);
  and (_18221_, _18220_, _12600_);
  or (_18222_, _18221_, _18208_);
  nor (_18223_, _17903_, _11287_);
  not (_18224_, _12549_);
  and (_18225_, _18224_, _18223_);
  nor (_18226_, _18224_, _18223_);
  nor (_18227_, _18226_, _18225_);
  and (_18228_, _17908_, _18227_);
  nor (_18229_, _17908_, _18227_);
  or (_18230_, _18229_, _10487_);
  or (_18231_, _18230_, _18228_);
  and (_18232_, _18231_, _18222_);
  or (_18233_, _18232_, _05976_);
  nand (_18234_, _06212_, _05976_);
  and (_18235_, _18234_, _06267_);
  and (_18236_, _18235_, _18233_);
  and (_18237_, _14943_, _08596_);
  or (_18238_, _18237_, _18126_);
  and (_18239_, _18238_, _06266_);
  or (_18240_, _18239_, _06259_);
  or (_18241_, _18240_, _18236_);
  and (_18242_, _18241_, _18108_);
  or (_18243_, _18242_, _09486_);
  and (_18244_, _09247_, _07930_);
  or (_18245_, _18105_, _06258_);
  or (_18246_, _18245_, _18244_);
  and (_18247_, _18246_, _06251_);
  and (_18248_, _18247_, _18243_);
  and (_18249_, _14998_, _07930_);
  or (_18250_, _18249_, _18105_);
  and (_18251_, _18250_, _05972_);
  or (_18252_, _18251_, _09480_);
  or (_18253_, _18252_, _18248_);
  or (_18254_, _10215_, _09481_);
  and (_18255_, _18254_, _18253_);
  or (_18256_, _18255_, _05984_);
  and (_18257_, _18256_, _18104_);
  or (_18258_, _18257_, _06215_);
  and (_18259_, _07930_, _08809_);
  or (_18260_, _18259_, _18105_);
  or (_18261_, _18260_, _06216_);
  and (_18262_, _18261_, _10892_);
  and (_18263_, _18262_, _18258_);
  or (_18264_, _10892_, _06212_);
  nand (_18265_, _18264_, _12694_);
  or (_18266_, _18265_, _18263_);
  or (_18267_, _12694_, _18111_);
  and (_18268_, _18267_, _06867_);
  and (_18269_, _18268_, _18266_);
  and (_18270_, _18111_, _06866_);
  or (_18271_, _18270_, _10916_);
  or (_18272_, _18271_, _18269_);
  nand (_18273_, _18196_, _10916_);
  nand (_18274_, _18273_, _18272_);
  nor (_18275_, _18274_, _06868_);
  and (_18276_, _18195_, _06868_);
  or (_18277_, _18276_, _06526_);
  or (_18278_, _18277_, _18275_);
  and (_18279_, _18278_, _18103_);
  nor (_18280_, _10935_, _12549_);
  or (_18281_, _18280_, _06398_);
  or (_18282_, _18281_, _18279_);
  and (_18283_, _14893_, _07930_);
  or (_18284_, _18283_, _18105_);
  or (_18285_, _18284_, _09025_);
  and (_18286_, _18285_, _18282_);
  or (_18287_, _18286_, _06524_);
  or (_18288_, _18105_, _09030_);
  and (_18289_, _18288_, _17973_);
  and (_18290_, _18289_, _18287_);
  or (_18291_, _18290_, _18101_);
  and (_18292_, _18291_, _17785_);
  and (_18293_, _11156_, _17784_);
  or (_18294_, _18293_, _18292_);
  and (_18295_, _18294_, _10964_);
  and (_18296_, _10959_, _11206_);
  or (_18297_, _18296_, _06530_);
  or (_18298_, _18297_, _18295_);
  or (_18299_, _11246_, _06531_);
  and (_18300_, _18299_, _10974_);
  and (_18301_, _18300_, _18298_);
  and (_18302_, _10968_, _11284_);
  or (_18303_, _18302_, _18301_);
  and (_18304_, _18303_, _07219_);
  nand (_18305_, _18260_, _06426_);
  nor (_18306_, _18305_, _11247_);
  or (_18307_, _18306_, _17394_);
  or (_18308_, _18307_, _18304_);
  and (_18309_, _18308_, _18100_);
  nor (_18310_, _11157_, _07061_);
  or (_18311_, _18310_, _18309_);
  and (_18312_, _18311_, _17229_);
  nor (_18313_, _11157_, _17229_);
  or (_18314_, _18313_, _11000_);
  or (_18315_, _18314_, _18312_);
  nand (_18316_, _11000_, _11207_);
  and (_18317_, _18316_, _06538_);
  and (_18318_, _18317_, _18315_);
  nand (_18319_, _11009_, _11247_);
  and (_18320_, _18319_, _11008_);
  or (_18321_, _18320_, _18318_);
  or (_18322_, _11009_, _11285_);
  and (_18323_, _18322_, _07229_);
  and (_18324_, _18323_, _18321_);
  and (_18325_, _14890_, _07930_);
  or (_18326_, _18325_, _18105_);
  and (_18327_, _18326_, _06437_);
  or (_18328_, _18327_, _11024_);
  or (_18329_, _18328_, _18324_);
  and (_18330_, _18329_, _18098_);
  or (_18331_, _18330_, _13990_);
  and (_18332_, _11067_, _10591_);
  nor (_18333_, _18332_, _11068_);
  or (_18334_, _18333_, _11027_);
  and (_18335_, _18334_, _06523_);
  and (_18336_, _18335_, _18331_);
  nand (_18337_, _11096_, _10523_);
  nor (_18338_, _11097_, _06523_);
  and (_18339_, _18338_, _18337_);
  or (_18340_, _18339_, _11082_);
  or (_18341_, _18340_, _18336_);
  and (_18342_, _11124_, _10830_);
  nor (_18343_, _18342_, _11125_);
  or (_18344_, _18343_, _11083_);
  and (_18345_, _18344_, _12775_);
  and (_18346_, _18345_, _18341_);
  or (_18347_, _17439_, _17435_);
  and (_18348_, _11111_, \oc8051_golden_model_1.ACC [2]);
  or (_18349_, _18348_, _18347_);
  or (_18350_, _18349_, _18346_);
  not (_18351_, _17438_);
  nor (_18352_, _11169_, _18111_);
  and (_18353_, _11169_, _18111_);
  or (_18354_, _18353_, _18352_);
  and (_18355_, _18354_, _18351_);
  or (_18356_, _18355_, _11185_);
  and (_18357_, _18356_, _18350_);
  and (_18358_, _18354_, _17438_);
  or (_18359_, _18358_, _11191_);
  or (_18360_, _18359_, _18357_);
  and (_18361_, _11221_, _18195_);
  nor (_18362_, _11221_, _18195_);
  or (_18363_, _18362_, _18361_);
  or (_18364_, _18363_, _11190_);
  and (_18365_, _18364_, _06293_);
  and (_18366_, _18365_, _18360_);
  and (_18367_, _11259_, _12529_);
  nor (_18368_, _11259_, _12529_);
  or (_18369_, _18368_, _18367_);
  and (_18370_, _18369_, _06292_);
  or (_18371_, _18370_, _10474_);
  or (_18372_, _18371_, _18366_);
  and (_18373_, _11297_, _18224_);
  nor (_18374_, _11297_, _18224_);
  or (_18375_, _18374_, _10475_);
  or (_18376_, _18375_, _18373_);
  and (_18377_, _18376_, _12981_);
  and (_18378_, _18377_, _18372_);
  and (_18379_, _10472_, \oc8051_golden_model_1.ACC [2]);
  or (_18380_, _18379_, _06559_);
  or (_18381_, _18380_, _18378_);
  or (_18382_, _18136_, _07240_);
  and (_18383_, _18382_, _11316_);
  and (_18384_, _18383_, _18381_);
  nor (_18385_, _11321_, _10248_);
  or (_18386_, _18385_, _11322_);
  and (_18387_, _18386_, _11315_);
  or (_18388_, _18387_, _11320_);
  or (_18389_, _18388_, _18384_);
  nand (_18390_, _11320_, _10123_);
  and (_18391_, _18390_, _05933_);
  and (_18392_, _18391_, _18389_);
  and (_18393_, _18178_, _05932_);
  or (_18394_, _18393_, _06566_);
  or (_18395_, _18394_, _18392_);
  and (_18396_, _15068_, _07930_);
  or (_18397_, _18396_, _18105_);
  or (_18398_, _18397_, _06570_);
  and (_18399_, _18398_, _11339_);
  and (_18400_, _18399_, _18395_);
  nor (_18401_, _11347_, \oc8051_golden_model_1.ACC [3]);
  nor (_18402_, _18401_, _11348_);
  and (_18403_, _18402_, _11338_);
  or (_18404_, _18403_, _11345_);
  or (_18405_, _18404_, _18400_);
  nand (_18406_, _11345_, _10123_);
  and (_18407_, _18406_, _01320_);
  and (_18408_, _18407_, _18405_);
  or (_18409_, _18408_, _18095_);
  and (_42902_, _18409_, _42355_);
  nor (_18410_, _01320_, _10123_);
  or (_18411_, _11223_, _11205_);
  and (_18412_, _18411_, _11224_);
  or (_18413_, _18412_, _17449_);
  or (_18414_, _11245_, _06527_);
  and (_18415_, _18414_, _10935_);
  not (_18416_, _12692_);
  and (_18417_, _11155_, _06869_);
  nand (_18418_, _06961_, _05984_);
  nor (_18419_, _07930_, _10123_);
  and (_18420_, _09420_, _07930_);
  or (_18421_, _18420_, _18419_);
  or (_18422_, _18421_, _06260_);
  nor (_18423_, _12535_, _10774_);
  or (_18424_, _18211_, _14093_);
  and (_18425_, _18424_, _14092_);
  nor (_18426_, _11245_, _18425_);
  and (_18427_, _11245_, _18425_);
  nor (_18428_, _18427_, _18426_);
  and (_18429_, _18428_, \oc8051_golden_model_1.PSW [7]);
  nor (_18430_, _18428_, \oc8051_golden_model_1.PSW [7]);
  nor (_18431_, _18430_, _18429_);
  and (_18432_, _18431_, _18423_);
  nor (_18433_, _18431_, _18423_);
  nor (_18434_, _18433_, _18432_);
  or (_18435_, _18434_, _06386_);
  and (_18436_, _18435_, _10487_);
  or (_18437_, _18122_, _18115_);
  and (_18438_, _09421_, _10248_);
  or (_18439_, _09421_, _10248_);
  and (_18440_, _18439_, _18110_);
  or (_18441_, _18440_, _18438_);
  nor (_18442_, _11155_, _18441_);
  and (_18443_, _11155_, _18441_);
  nor (_18444_, _18443_, _18442_);
  and (_18445_, _18444_, \oc8051_golden_model_1.PSW [7]);
  nor (_18446_, _18444_, \oc8051_golden_model_1.PSW [7]);
  nor (_18447_, _18446_, _18445_);
  or (_18448_, _18447_, _18437_);
  and (_18449_, _18447_, _18437_);
  nor (_18450_, _18449_, _10724_);
  and (_18451_, _18450_, _18448_);
  or (_18452_, _10623_, _09420_);
  nor (_18453_, _08596_, _10123_);
  and (_18454_, _15116_, _08596_);
  or (_18455_, _18454_, _18453_);
  or (_18456_, _18455_, _06282_);
  and (_18457_, _18456_, _07169_);
  and (_18458_, _15133_, _07930_);
  or (_18459_, _18458_, _18419_);
  and (_18460_, _18459_, _06285_);
  or (_18461_, _10634_, _09437_);
  and (_18462_, _10645_, _09420_);
  or (_18463_, _06755_, \oc8051_golden_model_1.ACC [4]);
  nand (_18464_, _06755_, \oc8051_golden_model_1.ACC [4]);
  nand (_18465_, _18464_, _18463_);
  nor (_18466_, _18465_, _10645_);
  or (_18467_, _18466_, _10633_);
  or (_18468_, _18467_, _18462_);
  and (_18469_, _18468_, _10636_);
  and (_18470_, _18469_, _18461_);
  or (_18471_, _18470_, _18460_);
  and (_18472_, _18471_, _10657_);
  nor (_18473_, _10660_, \oc8051_golden_model_1.ACC [4]);
  nor (_18474_, _18473_, _10661_);
  and (_18475_, _18474_, _10656_);
  or (_18476_, _18475_, _06281_);
  or (_18477_, _18476_, _18472_);
  and (_18478_, _18477_, _18457_);
  and (_18479_, _18421_, _06354_);
  or (_18480_, _18479_, _10622_);
  or (_18481_, _18480_, _18478_);
  and (_18482_, _18481_, _18452_);
  or (_18483_, _18482_, _07174_);
  or (_18484_, _09437_, _10692_);
  and (_18485_, _18484_, _06346_);
  and (_18486_, _18485_, _18483_);
  nor (_18487_, _08527_, _06346_);
  or (_18488_, _18487_, _10696_);
  or (_18489_, _18488_, _18486_);
  nand (_18490_, _10696_, _06018_);
  and (_18491_, _18490_, _18489_);
  or (_18492_, _18491_, _06277_);
  and (_18493_, _15145_, _08596_);
  or (_18494_, _18493_, _18453_);
  or (_18495_, _18494_, _06278_);
  and (_18496_, _18495_, _06271_);
  and (_18497_, _18496_, _18492_);
  or (_18498_, _18453_, _15152_);
  and (_18499_, _18498_, _06270_);
  and (_18500_, _18499_, _18455_);
  or (_18501_, _18500_, _09520_);
  or (_18502_, _18501_, _18497_);
  nor (_18503_, _10016_, _10014_);
  nor (_18504_, _18503_, _10017_);
  or (_18505_, _18504_, _10059_);
  and (_18506_, _18505_, _10724_);
  and (_18507_, _18506_, _18502_);
  or (_18508_, _18507_, _18451_);
  and (_18509_, _18508_, _10555_);
  nand (_18510_, _18203_, _18200_);
  and (_18511_, _09247_, _10248_);
  or (_18512_, _09247_, _10248_);
  and (_18513_, _18512_, _18194_);
  or (_18514_, _18513_, _18511_);
  nor (_18515_, _11205_, _18514_);
  not (_18516_, _18515_);
  nand (_18517_, _11205_, _18514_);
  and (_18518_, _18517_, _18516_);
  nand (_18519_, _18518_, \oc8051_golden_model_1.PSW [7]);
  or (_18520_, _18518_, \oc8051_golden_model_1.PSW [7]);
  and (_18521_, _18520_, _18519_);
  or (_18522_, _18521_, _18510_);
  nand (_18523_, _18521_, _18510_);
  and (_18524_, _10727_, _18523_);
  and (_18525_, _18524_, _18522_);
  or (_18526_, _18525_, _06380_);
  or (_18527_, _18526_, _18509_);
  and (_18528_, _18527_, _18436_);
  nor (_18529_, _12554_, _10774_);
  nor (_18530_, _18223_, _12547_);
  nor (_18531_, _18530_, _12548_);
  nor (_18532_, _11283_, _18531_);
  and (_18533_, _11283_, _18531_);
  nor (_18534_, _18533_, _18532_);
  and (_18535_, _18534_, \oc8051_golden_model_1.PSW [7]);
  nor (_18536_, _18534_, \oc8051_golden_model_1.PSW [7]);
  nor (_18537_, _18536_, _18535_);
  or (_18538_, _18537_, _18529_);
  and (_18539_, _18537_, _18529_);
  nor (_18540_, _18539_, _10487_);
  and (_18541_, _18540_, _18538_);
  or (_18542_, _18541_, _05976_);
  or (_18543_, _18542_, _18528_);
  nand (_18544_, _06961_, _05976_);
  and (_18545_, _18544_, _06267_);
  and (_18546_, _18545_, _18543_);
  and (_18547_, _15170_, _08596_);
  or (_18548_, _18547_, _18453_);
  and (_18549_, _18548_, _06266_);
  or (_18550_, _18549_, _06259_);
  or (_18551_, _18550_, _18546_);
  and (_18552_, _18551_, _18422_);
  or (_18553_, _18552_, _09486_);
  and (_18554_, _09437_, _07930_);
  or (_18555_, _18419_, _06258_);
  or (_18556_, _18555_, _18554_);
  and (_18557_, _18556_, _06251_);
  and (_18558_, _18557_, _18553_);
  and (_18559_, _15226_, _07930_);
  or (_18560_, _18559_, _18419_);
  and (_18561_, _18560_, _05972_);
  or (_18562_, _18561_, _09480_);
  or (_18563_, _18562_, _18558_);
  or (_18564_, _10165_, _09481_);
  and (_18565_, _18564_, _18563_);
  or (_18566_, _18565_, _05984_);
  and (_18567_, _18566_, _18418_);
  or (_18568_, _18567_, _06215_);
  and (_18569_, _08919_, _07930_);
  or (_18570_, _18569_, _18419_);
  or (_18571_, _18570_, _06216_);
  and (_18572_, _18571_, _10892_);
  and (_18573_, _18572_, _18568_);
  and (_18574_, _06338_, _06000_);
  nor (_18575_, _10892_, _06961_);
  or (_18576_, _18575_, _18574_);
  or (_18577_, _18576_, _18573_);
  and (_18578_, _11155_, _06255_);
  or (_18579_, _18578_, _17790_);
  and (_18580_, _18579_, _18577_);
  nor (_18581_, _17790_, _06255_);
  and (_18582_, _18581_, _11155_);
  or (_18583_, _18582_, _17789_);
  or (_18584_, _18583_, _18580_);
  not (_18585_, _06869_);
  or (_18586_, _11155_, _17949_);
  and (_18587_, _18586_, _18585_);
  and (_18588_, _18587_, _18584_);
  or (_18589_, _18588_, _18417_);
  and (_18590_, _18589_, _18416_);
  and (_18591_, _12692_, _11155_);
  or (_18592_, _18591_, _06866_);
  or (_18593_, _18592_, _18590_);
  or (_18594_, _11155_, _06867_);
  and (_18595_, _18594_, _10918_);
  and (_18596_, _18595_, _18593_);
  and (_18597_, _11205_, _10917_);
  or (_18598_, _18597_, _06526_);
  or (_18599_, _18598_, _18596_);
  and (_18600_, _18599_, _18415_);
  nor (_18601_, _10935_, _11282_);
  or (_18602_, _18601_, _06398_);
  or (_18603_, _18602_, _18600_);
  and (_18604_, _15114_, _07930_);
  or (_18605_, _18604_, _18419_);
  or (_18606_, _18605_, _09025_);
  and (_18607_, _18606_, _18603_);
  or (_18608_, _18607_, _06524_);
  or (_18609_, _18419_, _09030_);
  and (_18610_, _18609_, _12243_);
  and (_18611_, _18610_, _18608_);
  or (_18612_, _10959_, _11152_);
  and (_18613_, _18612_, _12720_);
  or (_18614_, _18613_, _18611_);
  or (_18615_, _10964_, _11202_);
  and (_18616_, _18615_, _18614_);
  or (_18617_, _18616_, _06530_);
  or (_18618_, _11242_, _06531_);
  and (_18619_, _18618_, _10974_);
  and (_18620_, _18619_, _18617_);
  and (_18621_, _10968_, _11279_);
  or (_18622_, _18621_, _18620_);
  and (_18623_, _18622_, _07219_);
  not (_18624_, _17397_);
  nand (_18625_, _18570_, _06426_);
  nor (_18626_, _18625_, _11244_);
  or (_18627_, _18626_, _18624_);
  or (_18628_, _18627_, _18623_);
  or (_18629_, _17397_, _11154_);
  and (_18630_, _18629_, _17229_);
  and (_18631_, _18630_, _18628_);
  and (_18632_, _11154_, _17228_);
  or (_18633_, _18632_, _11000_);
  or (_18634_, _18633_, _18631_);
  or (_18635_, _17689_, _11204_);
  and (_18636_, _18635_, _06538_);
  and (_18637_, _18636_, _18634_);
  nand (_18638_, _11009_, _11244_);
  and (_18639_, _18638_, _11008_);
  or (_18640_, _18639_, _18637_);
  nand (_18641_, _11006_, _11281_);
  and (_18642_, _18641_, _18640_);
  or (_18643_, _18642_, _06437_);
  and (_18644_, _15111_, _07930_);
  or (_18645_, _18419_, _07229_);
  or (_18646_, _18645_, _18644_);
  and (_18647_, _18646_, _11023_);
  and (_18648_, _18647_, _18643_);
  or (_18649_, _11042_, _10754_);
  and (_18650_, _18649_, _11043_);
  and (_18651_, _18650_, _11024_);
  or (_18652_, _18651_, _11026_);
  or (_18653_, _18652_, _18648_);
  or (_18654_, _11069_, _10585_);
  and (_18655_, _18654_, _11070_);
  or (_18656_, _18655_, _17490_);
  and (_18657_, _18656_, _18653_);
  or (_18658_, _18657_, _06892_);
  or (_18659_, _18655_, _17717_);
  and (_18660_, _18659_, _06523_);
  and (_18661_, _18660_, _18658_);
  or (_18662_, _11098_, _10517_);
  and (_18663_, _11099_, _06522_);
  and (_18664_, _18663_, _18662_);
  or (_18665_, _18664_, _18661_);
  and (_18666_, _18665_, _11083_);
  or (_18667_, _11126_, _10824_);
  and (_18668_, _11127_, _11082_);
  and (_18669_, _18668_, _18667_);
  or (_18670_, _18669_, _11111_);
  or (_18671_, _18670_, _18666_);
  nand (_18672_, _11111_, _10248_);
  and (_18673_, _18672_, _11185_);
  and (_18674_, _18673_, _18671_);
  or (_18675_, _11171_, _11155_);
  nor (_18676_, _11185_, _11172_);
  and (_18677_, _18676_, _18675_);
  or (_18678_, _18677_, _11189_);
  or (_18679_, _18678_, _18674_);
  and (_18680_, _18679_, _18413_);
  or (_18681_, _18680_, _11188_);
  or (_18682_, _18412_, _17448_);
  and (_18683_, _18682_, _06293_);
  and (_18684_, _18683_, _18681_);
  or (_18685_, _11261_, _11245_);
  and (_18686_, _18685_, _11262_);
  or (_18687_, _18686_, _10474_);
  and (_18688_, _18687_, _12979_);
  or (_18689_, _18688_, _18684_);
  or (_18690_, _11300_, _11283_);
  and (_18691_, _18690_, _11301_);
  or (_18692_, _18691_, _10475_);
  and (_18693_, _18692_, _12981_);
  and (_18694_, _18693_, _18689_);
  and (_18695_, _10472_, \oc8051_golden_model_1.ACC [3]);
  or (_18696_, _18695_, _06559_);
  or (_18697_, _18696_, _18694_);
  or (_18698_, _18459_, _07240_);
  and (_18699_, _18698_, _11316_);
  and (_18700_, _18699_, _18697_);
  nor (_18701_, _11322_, _10123_);
  or (_18702_, _18701_, _11323_);
  and (_18703_, _18702_, _11315_);
  or (_18704_, _18703_, _11320_);
  or (_18705_, _18704_, _18700_);
  nand (_18706_, _11320_, _10152_);
  and (_18707_, _18706_, _05933_);
  and (_18708_, _18707_, _18705_);
  and (_18709_, _18494_, _05932_);
  or (_18710_, _18709_, _06566_);
  or (_18711_, _18710_, _18708_);
  and (_18712_, _15296_, _07930_);
  or (_18713_, _18712_, _18419_);
  or (_18714_, _18713_, _06570_);
  and (_18715_, _18714_, _11339_);
  and (_18716_, _18715_, _18711_);
  nor (_18717_, _11348_, \oc8051_golden_model_1.ACC [4]);
  nor (_18718_, _18717_, _11349_);
  and (_18719_, _18718_, _11338_);
  or (_18720_, _18719_, _11345_);
  or (_18721_, _18720_, _18716_);
  nand (_18722_, _11345_, _10152_);
  and (_18723_, _18722_, _01320_);
  and (_18724_, _18723_, _18721_);
  or (_18725_, _18724_, _18410_);
  and (_42903_, _18725_, _42355_);
  nor (_18726_, _01320_, _10152_);
  nor (_18727_, _11174_, _11151_);
  nor (_18728_, _18727_, _11175_);
  or (_18729_, _18728_, _11185_);
  and (_18730_, _11044_, _10751_);
  nor (_18731_, _18730_, _11045_);
  or (_18732_, _18731_, _11023_);
  nand (_18733_, _10986_, _11150_);
  or (_18734_, _10964_, _11199_);
  nor (_18735_, _07930_, _10152_);
  and (_18736_, _18735_, _06524_);
  and (_18737_, _12536_, _06526_);
  and (_18738_, _06339_, _06000_);
  nor (_18739_, _18738_, _06863_);
  not (_18740_, _18739_);
  and (_18741_, _18740_, _11151_);
  nand (_18742_, _06604_, _05984_);
  and (_18743_, _09419_, _07930_);
  or (_18744_, _18743_, _18735_);
  or (_18745_, _18744_, _06260_);
  and (_18746_, _06961_, \oc8051_golden_model_1.ACC [4]);
  nor (_18747_, _18532_, _18746_);
  nor (_18748_, _12555_, _18747_);
  and (_18749_, _12555_, _18747_);
  nor (_18750_, _18749_, _18748_);
  and (_18751_, _18750_, \oc8051_golden_model_1.PSW [7]);
  nor (_18752_, _18750_, \oc8051_golden_model_1.PSW [7]);
  nor (_18753_, _18752_, _18751_);
  nor (_18754_, _18539_, _18535_);
  not (_18755_, _18754_);
  and (_18756_, _18755_, _18753_);
  nor (_18757_, _18755_, _18753_);
  nor (_18758_, _18757_, _18756_);
  or (_18759_, _18758_, _10487_);
  and (_18760_, _09202_, \oc8051_golden_model_1.ACC [4]);
  nor (_18761_, _18515_, _18760_);
  or (_18762_, _11201_, _18761_);
  nand (_18763_, _11201_, _18761_);
  and (_18764_, _18763_, _18762_);
  or (_18765_, _18764_, _10774_);
  nand (_18766_, _18764_, _10774_);
  and (_18767_, _18766_, _18765_);
  nand (_18768_, _18523_, _18519_);
  nand (_18769_, _18768_, _18767_);
  or (_18770_, _18768_, _18767_);
  and (_18771_, _18770_, _18769_);
  or (_18772_, _18771_, _10555_);
  and (_18773_, _08525_, \oc8051_golden_model_1.ACC [4]);
  nor (_18774_, _18442_, _18773_);
  nor (_18775_, _11151_, _18774_);
  and (_18777_, _11151_, _18774_);
  nor (_18778_, _18777_, _18775_);
  and (_18779_, _18778_, \oc8051_golden_model_1.PSW [7]);
  nor (_18780_, _18778_, \oc8051_golden_model_1.PSW [7]);
  nor (_18781_, _18780_, _18779_);
  nor (_18782_, _18449_, _18445_);
  not (_18783_, _18782_);
  and (_18784_, _18783_, _18781_);
  nor (_18785_, _18783_, _18781_);
  nor (_18786_, _18785_, _18784_);
  or (_18788_, _18786_, _10724_);
  nor (_18789_, _08596_, _10152_);
  and (_18790_, _15315_, _08596_);
  or (_18791_, _18790_, _18789_);
  or (_18792_, _18789_, _15349_);
  and (_18793_, _18792_, _06270_);
  and (_18794_, _18793_, _18791_);
  or (_18795_, _10623_, _09419_);
  or (_18796_, _18138_, _09419_);
  nor (_18797_, _06755_, _10152_);
  and (_18799_, _06755_, _10152_);
  or (_18800_, _18799_, _18797_);
  or (_18801_, _18800_, _10645_);
  and (_18802_, _18801_, _10634_);
  and (_18803_, _18802_, _18796_);
  and (_18804_, _10633_, _09436_);
  or (_18805_, _18804_, _18803_);
  and (_18806_, _18805_, _10636_);
  and (_18807_, _15330_, _07930_);
  or (_18808_, _18807_, _18735_);
  and (_18810_, _18808_, _06285_);
  or (_18811_, _18810_, _10656_);
  or (_18812_, _18811_, _18806_);
  nor (_18813_, _10678_, _10669_);
  nand (_18814_, _10678_, _10669_);
  nand (_18815_, _18814_, _10656_);
  or (_18816_, _18815_, _18813_);
  and (_18817_, _18816_, _06361_);
  and (_18818_, _18817_, _18812_);
  and (_18819_, _18791_, _06281_);
  and (_18821_, _18744_, _06354_);
  or (_18822_, _18821_, _10622_);
  or (_18823_, _18822_, _18819_);
  or (_18824_, _18823_, _18818_);
  and (_18825_, _18824_, _18795_);
  or (_18826_, _18825_, _07174_);
  or (_18827_, _09436_, _10692_);
  and (_18828_, _18827_, _06346_);
  and (_18829_, _18828_, _18826_);
  nor (_18830_, _08230_, _06346_);
  or (_18832_, _18830_, _10696_);
  or (_18833_, _18832_, _18829_);
  nand (_18834_, _10696_, _06044_);
  and (_18835_, _18834_, _18833_);
  or (_18836_, _18835_, _06277_);
  and (_18837_, _15342_, _08596_);
  or (_18838_, _18837_, _18789_);
  or (_18839_, _18838_, _06278_);
  and (_18840_, _18839_, _06271_);
  and (_18841_, _18840_, _18836_);
  or (_18843_, _18841_, _18794_);
  and (_18844_, _18843_, _10059_);
  or (_18845_, _10019_, _10017_);
  nor (_18846_, _10020_, _10059_);
  and (_18847_, _18846_, _18845_);
  or (_18848_, _18847_, _17293_);
  or (_18849_, _18848_, _18844_);
  and (_18850_, _18849_, _18788_);
  or (_18851_, _18850_, _10727_);
  and (_18852_, _18851_, _06386_);
  and (_18854_, _18852_, _18772_);
  and (_18855_, _08527_, \oc8051_golden_model_1.ACC [4]);
  nor (_18856_, _18426_, _18855_);
  nor (_18857_, _12536_, _18856_);
  and (_18858_, _12536_, _18856_);
  nor (_18859_, _18858_, _18857_);
  and (_18860_, _18859_, \oc8051_golden_model_1.PSW [7]);
  nor (_18861_, _18859_, \oc8051_golden_model_1.PSW [7]);
  nor (_18862_, _18861_, _18860_);
  nor (_18863_, _18432_, _18429_);
  not (_18865_, _18863_);
  and (_18866_, _18865_, _18862_);
  nor (_18867_, _18865_, _18862_);
  nor (_18868_, _18867_, _18866_);
  or (_18869_, _18868_, _10486_);
  and (_18870_, _18869_, _12600_);
  or (_18871_, _18870_, _18854_);
  and (_18872_, _18871_, _18759_);
  or (_18873_, _18872_, _05976_);
  nand (_18874_, _06604_, _05976_);
  and (_18876_, _18874_, _06267_);
  and (_18877_, _18876_, _18873_);
  or (_18878_, _18789_, _15365_);
  and (_18879_, _18878_, _06266_);
  and (_18880_, _18879_, _18791_);
  or (_18881_, _18880_, _06259_);
  or (_18882_, _18881_, _18877_);
  and (_18883_, _18882_, _18745_);
  or (_18884_, _18883_, _09486_);
  and (_18885_, _09436_, _07930_);
  or (_18887_, _18735_, _06258_);
  or (_18888_, _18887_, _18885_);
  and (_18889_, _18888_, _06251_);
  and (_18890_, _18889_, _18884_);
  and (_18891_, _15421_, _07930_);
  or (_18892_, _18891_, _18735_);
  and (_18893_, _18892_, _05972_);
  or (_18894_, _18893_, _09480_);
  or (_18895_, _18894_, _18890_);
  or (_18896_, _10137_, _09481_);
  and (_18898_, _18896_, _18895_);
  or (_18899_, _18898_, _05984_);
  and (_18900_, _18899_, _18742_);
  or (_18901_, _18900_, _06215_);
  and (_18902_, _08913_, _07930_);
  or (_18903_, _18902_, _18735_);
  or (_18904_, _18903_, _06216_);
  and (_18905_, _18904_, _10892_);
  and (_18906_, _18905_, _18901_);
  nor (_18907_, _10892_, _06604_);
  or (_18909_, _18907_, _18574_);
  or (_18910_, _18909_, _18906_);
  not (_18911_, _18574_);
  or (_18912_, _11151_, _18911_);
  and (_18913_, _18912_, _18739_);
  and (_18914_, _18913_, _18910_);
  nor (_18915_, _18914_, _18741_);
  nor (_18916_, _18915_, _06864_);
  and (_18917_, _11151_, _06864_);
  or (_18918_, _18917_, _17789_);
  or (_18920_, _18918_, _18916_);
  or (_18921_, _11151_, _17949_);
  and (_18922_, _18921_, _17953_);
  and (_18923_, _18922_, _18920_);
  and (_18924_, _17952_, _11151_);
  or (_18925_, _18924_, _10917_);
  or (_18926_, _18925_, _18923_);
  nand (_18927_, _11201_, _10917_);
  and (_18928_, _18927_, _06527_);
  and (_18929_, _18928_, _18926_);
  or (_18931_, _18929_, _18737_);
  and (_18932_, _18931_, _10935_);
  and (_18933_, _10481_, _12555_);
  or (_18934_, _18933_, _06398_);
  or (_18935_, _18934_, _18932_);
  and (_18936_, _15313_, _07930_);
  or (_18937_, _18936_, _18735_);
  or (_18938_, _18937_, _09025_);
  and (_18939_, _18938_, _09030_);
  and (_18940_, _18939_, _18935_);
  or (_18942_, _18940_, _18736_);
  and (_18943_, _18942_, _10948_);
  and (_18944_, _06714_, _06012_);
  nor (_18945_, _07066_, _18944_);
  nand (_18946_, _11149_, _10944_);
  nand (_18947_, _18946_, _18945_);
  or (_18948_, _18947_, _18943_);
  and (_18949_, _17951_, _06012_);
  nor (_18950_, _18945_, _11149_);
  nor (_18951_, _18950_, _18949_);
  and (_18952_, _18951_, _18948_);
  and (_18953_, _18949_, _11149_);
  or (_18954_, _18953_, _10959_);
  or (_18955_, _18954_, _18952_);
  and (_18956_, _18955_, _18734_);
  or (_18957_, _18956_, _06530_);
  or (_18958_, _11240_, _06531_);
  and (_18959_, _18958_, _10974_);
  and (_18960_, _18959_, _18957_);
  and (_18961_, _10968_, _11277_);
  or (_18963_, _18961_, _18960_);
  and (_18964_, _18963_, _07219_);
  nand (_18965_, _18903_, _06426_);
  nor (_18966_, _18965_, _11241_);
  or (_18967_, _18966_, _10986_);
  or (_18968_, _18967_, _18964_);
  and (_18969_, _18968_, _18733_);
  or (_18970_, _18969_, _10991_);
  nand (_18971_, _10991_, _11150_);
  and (_18972_, _18971_, _10995_);
  and (_18974_, _18972_, _18970_);
  nor (_18975_, _11150_, _10995_);
  or (_18976_, _18975_, _11000_);
  or (_18977_, _18976_, _18974_);
  nand (_18978_, _11000_, _10152_);
  or (_18979_, _18978_, _09436_);
  and (_18980_, _18979_, _06538_);
  and (_18981_, _18980_, _18977_);
  nand (_18982_, _11009_, _11241_);
  and (_18983_, _18982_, _11008_);
  or (_18985_, _18983_, _18981_);
  nand (_18986_, _11006_, _11278_);
  and (_18987_, _18986_, _07229_);
  and (_18988_, _18987_, _18985_);
  and (_18989_, _15310_, _07930_);
  or (_18990_, _18989_, _18735_);
  and (_18991_, _18990_, _06437_);
  or (_18992_, _18991_, _11024_);
  or (_18993_, _18992_, _18988_);
  and (_18994_, _18993_, _18732_);
  or (_18996_, _18994_, _13990_);
  and (_18997_, _11071_, _10582_);
  nor (_18998_, _18997_, _11072_);
  or (_18999_, _18998_, _11027_);
  and (_19000_, _18999_, _06523_);
  and (_19001_, _19000_, _18996_);
  and (_19002_, _11100_, _10514_);
  nor (_19003_, _19002_, _11101_);
  or (_19004_, _19003_, _11082_);
  and (_19005_, _19004_, _12770_);
  or (_19007_, _19005_, _19001_);
  and (_19008_, _11128_, _10818_);
  nor (_19009_, _19008_, _11129_);
  or (_19010_, _19009_, _11083_);
  and (_19011_, _19010_, _12775_);
  and (_19012_, _19011_, _19007_);
  and (_19013_, _11111_, \oc8051_golden_model_1.ACC [4]);
  or (_19014_, _11140_, _11144_);
  or (_19015_, _19014_, _19013_);
  or (_19016_, _19015_, _10476_);
  or (_19018_, _19016_, _19012_);
  and (_19019_, _19018_, _18729_);
  or (_19020_, _19019_, _11191_);
  and (_19021_, _11225_, _11201_);
  nor (_19022_, _19021_, _11226_);
  or (_19023_, _19022_, _11190_);
  and (_19024_, _19023_, _06293_);
  and (_19025_, _19024_, _19020_);
  and (_19026_, _11263_, _12536_);
  nor (_19027_, _11263_, _12536_);
  or (_19029_, _19027_, _10474_);
  or (_19030_, _19029_, _19026_);
  and (_19031_, _19030_, _12979_);
  or (_19032_, _19031_, _19025_);
  and (_19033_, _11302_, _12555_);
  nor (_19034_, _11302_, _12555_);
  or (_19035_, _19034_, _10475_);
  or (_19036_, _19035_, _19033_);
  and (_19037_, _19036_, _12981_);
  and (_19038_, _19037_, _19032_);
  and (_19040_, _10472_, \oc8051_golden_model_1.ACC [4]);
  or (_19041_, _19040_, _06559_);
  or (_19042_, _19041_, _19038_);
  or (_19043_, _18808_, _07240_);
  and (_19044_, _19043_, _11316_);
  and (_19045_, _19044_, _19042_);
  nor (_19046_, _11323_, _10152_);
  or (_19047_, _19046_, _11324_);
  and (_19048_, _19047_, _11315_);
  or (_19049_, _19048_, _11320_);
  or (_19051_, _19049_, _19045_);
  nand (_19052_, _11320_, _10105_);
  and (_19053_, _19052_, _05933_);
  and (_19054_, _19053_, _19051_);
  and (_19055_, _18838_, _05932_);
  or (_19056_, _19055_, _06566_);
  or (_19057_, _19056_, _19054_);
  and (_19058_, _15493_, _07930_);
  or (_19059_, _19058_, _18735_);
  or (_19060_, _19059_, _06570_);
  and (_19062_, _19060_, _11339_);
  and (_19063_, _19062_, _19057_);
  nor (_19064_, _11349_, \oc8051_golden_model_1.ACC [5]);
  nor (_19065_, _19064_, _11350_);
  and (_19066_, _19065_, _11338_);
  or (_19067_, _19066_, _11345_);
  or (_19068_, _19067_, _19063_);
  nand (_19069_, _11345_, _10105_);
  and (_19070_, _19069_, _01320_);
  and (_19071_, _19070_, _19068_);
  or (_19073_, _19071_, _18726_);
  and (_42904_, _19073_, _42355_);
  nor (_19074_, _01320_, _10105_);
  or (_19075_, _11102_, _10547_);
  and (_19076_, _11103_, _06522_);
  and (_19077_, _19076_, _19075_);
  nand (_19078_, _11006_, _11275_);
  or (_19079_, _11236_, _06531_);
  and (_19080_, _19079_, _10974_);
  nor (_19081_, _07930_, _10105_);
  and (_19083_, _19081_, _06524_);
  and (_19084_, _11148_, _17789_);
  and (_19085_, _15623_, _07930_);
  or (_19086_, _19085_, _19081_);
  and (_19087_, _19086_, _05972_);
  and (_19088_, _09418_, _07930_);
  or (_19089_, _19088_, _19081_);
  or (_19090_, _19089_, _06260_);
  or (_19091_, _18747_, _14119_);
  and (_19092_, _19091_, _14118_);
  nor (_19094_, _19092_, _11276_);
  and (_19095_, _19092_, _11276_);
  nor (_19096_, _19095_, _19094_);
  nor (_19097_, _18756_, _18751_);
  and (_19098_, _19097_, \oc8051_golden_model_1.PSW [7]);
  or (_19099_, _19098_, _19096_);
  nand (_19100_, _19098_, _19096_);
  and (_19101_, _19100_, _10486_);
  and (_19102_, _19101_, _19099_);
  or (_19103_, _19102_, _05976_);
  or (_19105_, _10623_, _09418_);
  or (_19106_, _10634_, _09435_);
  or (_19107_, _18138_, _09418_);
  nor (_19108_, _06755_, _10105_);
  and (_19109_, _06755_, _10105_);
  or (_19110_, _19109_, _19108_);
  or (_19111_, _19110_, _10645_);
  and (_19112_, _19111_, _19107_);
  or (_19113_, _19112_, _10633_);
  and (_19114_, _19113_, _10636_);
  and (_19116_, _19114_, _19106_);
  and (_19117_, _15521_, _07930_);
  or (_19118_, _19117_, _19081_);
  and (_19119_, _19118_, _06285_);
  or (_19120_, _19119_, _10656_);
  or (_19121_, _19120_, _19116_);
  or (_19122_, _18813_, _10671_);
  nand (_19123_, _18813_, _10671_);
  and (_19124_, _19123_, _19122_);
  or (_19125_, _19124_, _10657_);
  and (_19127_, _19125_, _06361_);
  and (_19128_, _19127_, _19121_);
  nor (_19129_, _08596_, _10105_);
  and (_19130_, _15535_, _08596_);
  or (_19131_, _19130_, _19129_);
  and (_19132_, _19131_, _06281_);
  and (_19133_, _19089_, _06354_);
  or (_19134_, _19133_, _10622_);
  or (_19135_, _19134_, _19132_);
  or (_19136_, _19135_, _19128_);
  and (_19138_, _19136_, _19105_);
  or (_19139_, _19138_, _07174_);
  or (_19140_, _09435_, _10692_);
  and (_19141_, _19140_, _06346_);
  and (_19142_, _19141_, _19139_);
  nor (_19143_, _08127_, _06346_);
  or (_19144_, _19143_, _10696_);
  or (_19145_, _19144_, _19142_);
  nand (_19146_, _10696_, _10198_);
  and (_19147_, _19146_, _19145_);
  or (_19149_, _19147_, _06277_);
  and (_19150_, _15544_, _08596_);
  or (_19151_, _19150_, _19129_);
  or (_19152_, _19151_, _06278_);
  and (_19153_, _19152_, _06271_);
  and (_19154_, _19153_, _19149_);
  or (_19155_, _19129_, _15551_);
  and (_19156_, _19155_, _06270_);
  and (_19157_, _19156_, _19131_);
  or (_19158_, _19157_, _09520_);
  or (_19160_, _19158_, _19154_);
  nor (_19161_, _10022_, _10020_);
  nor (_19162_, _19161_, _10023_);
  or (_19163_, _19162_, _10059_);
  and (_19164_, _19163_, _10724_);
  and (_19165_, _19164_, _19160_);
  or (_19166_, _09419_, _10152_);
  and (_19167_, _09419_, _10152_);
  or (_19168_, _18774_, _19167_);
  and (_19169_, _19168_, _19166_);
  nor (_19171_, _19169_, _11148_);
  and (_19172_, _19169_, _11148_);
  nor (_19173_, _19172_, _19171_);
  nor (_19174_, _18784_, _18779_);
  and (_19175_, _19174_, \oc8051_golden_model_1.PSW [7]);
  or (_19176_, _19175_, _19173_);
  nand (_19177_, _19175_, _19173_);
  and (_19178_, _19177_, _19176_);
  and (_19179_, _19178_, _17293_);
  or (_19180_, _19179_, _19165_);
  and (_19182_, _19180_, _10555_);
  or (_19183_, _09436_, _10152_);
  and (_19184_, _09436_, _10152_);
  or (_19185_, _18761_, _19184_);
  and (_19186_, _19185_, _19183_);
  nor (_19187_, _19186_, _11198_);
  and (_19188_, _19186_, _11198_);
  nor (_19189_, _19188_, _19187_);
  and (_19190_, _18769_, _18765_);
  and (_19191_, _19190_, \oc8051_golden_model_1.PSW [7]);
  nand (_19193_, _19191_, _19189_);
  or (_19194_, _19191_, _19189_);
  and (_19195_, _10727_, _19194_);
  and (_19196_, _19195_, _19193_);
  or (_19197_, _19196_, _19182_);
  and (_19198_, _19197_, _12599_);
  or (_19199_, _18856_, _14082_);
  and (_19200_, _19199_, _14081_);
  nor (_19201_, _19200_, _11239_);
  and (_19202_, _19200_, _11239_);
  nor (_19204_, _19202_, _19201_);
  nor (_19205_, _18866_, _18860_);
  and (_19206_, _19205_, \oc8051_golden_model_1.PSW [7]);
  nand (_19207_, _19206_, _19204_);
  or (_19208_, _19206_, _19204_);
  and (_19209_, _19208_, _06380_);
  and (_19210_, _19209_, _19207_);
  or (_19211_, _19210_, _19198_);
  or (_19212_, _19211_, _19103_);
  nand (_19213_, _06325_, _05976_);
  and (_19215_, _19213_, _06267_);
  and (_19216_, _19215_, _19212_);
  and (_19217_, _15568_, _08596_);
  or (_19218_, _19217_, _19129_);
  and (_19219_, _19218_, _06266_);
  or (_19220_, _19219_, _06259_);
  or (_19221_, _19220_, _19216_);
  and (_19222_, _19221_, _19090_);
  or (_19223_, _19222_, _09486_);
  and (_19224_, _09435_, _07930_);
  or (_19226_, _19081_, _06258_);
  or (_19227_, _19226_, _19224_);
  and (_19228_, _19227_, _06251_);
  and (_19229_, _19228_, _19223_);
  or (_19230_, _19229_, _19087_);
  and (_19231_, _19230_, _12252_);
  nor (_19232_, _06325_, _05985_);
  not (_19233_, _10110_);
  nor (_19234_, _19233_, _10106_);
  and (_19235_, _19234_, _05935_);
  and (_19237_, _19235_, _09480_);
  or (_19238_, _19237_, _19232_);
  or (_19239_, _19238_, _19231_);
  and (_19240_, _19239_, _06216_);
  and (_19241_, _08845_, _07930_);
  or (_19242_, _19241_, _19081_);
  and (_19243_, _19242_, _06215_);
  or (_19244_, _19243_, _10891_);
  or (_19245_, _19244_, _19240_);
  and (_19246_, _06702_, _06000_);
  and (_19248_, _10891_, _06325_);
  nor (_19249_, _19248_, _19246_);
  and (_19250_, _19249_, _19245_);
  nand (_19251_, _11148_, _19246_);
  nor (_19252_, _18738_, _06864_);
  nand (_19253_, _19252_, _19251_);
  or (_19254_, _19253_, _19250_);
  or (_19255_, _19252_, _11148_);
  and (_19256_, _19255_, _17949_);
  and (_19257_, _19256_, _19254_);
  or (_19259_, _19257_, _19084_);
  and (_19260_, _19259_, _18585_);
  and (_19261_, _11148_, _06869_);
  or (_19262_, _19261_, _19260_);
  and (_19263_, _19262_, _18416_);
  and (_19264_, _12692_, _11148_);
  or (_19265_, _19264_, _06866_);
  or (_19266_, _19265_, _19263_);
  or (_19267_, _11148_, _06867_);
  and (_19268_, _19267_, _10918_);
  and (_19270_, _19268_, _19266_);
  and (_19271_, _11198_, _10917_);
  or (_19272_, _19271_, _06526_);
  or (_19273_, _19272_, _19270_);
  or (_19274_, _11239_, _06527_);
  and (_19275_, _19274_, _10935_);
  and (_19276_, _19275_, _19273_);
  and (_19277_, _10481_, _11276_);
  or (_19278_, _19277_, _06398_);
  or (_19279_, _19278_, _19276_);
  and (_19281_, _15517_, _07930_);
  or (_19282_, _19281_, _19081_);
  or (_19283_, _19282_, _09025_);
  and (_19284_, _19283_, _09030_);
  and (_19285_, _19284_, _19279_);
  or (_19286_, _19285_, _19083_);
  and (_19287_, _19286_, _12243_);
  nor (_19288_, _12243_, _11146_);
  or (_19289_, _19288_, _19287_);
  and (_19290_, _19289_, _10964_);
  and (_19292_, _10959_, _11195_);
  or (_19293_, _19292_, _06530_);
  or (_19294_, _19293_, _19290_);
  and (_19295_, _19294_, _19080_);
  and (_19296_, _10968_, _11274_);
  or (_19297_, _19296_, _19295_);
  and (_19298_, _19297_, _07219_);
  nand (_19299_, _19242_, _06426_);
  nor (_19300_, _19299_, _11238_);
  or (_19301_, _19300_, _18624_);
  or (_19303_, _19301_, _19298_);
  or (_19304_, _17397_, _11147_);
  and (_19305_, _19304_, _17229_);
  and (_19306_, _19305_, _19303_);
  and (_19307_, _11147_, _17228_);
  or (_19308_, _19307_, _11000_);
  or (_19309_, _19308_, _19306_);
  or (_19310_, _17689_, _11197_);
  and (_19311_, _19310_, _06538_);
  and (_19312_, _19311_, _19309_);
  nand (_19314_, _11009_, _11238_);
  and (_19315_, _19314_, _11008_);
  or (_19316_, _19315_, _19312_);
  and (_19317_, _19316_, _19078_);
  or (_19318_, _19317_, _06437_);
  and (_19319_, _15514_, _07930_);
  or (_19320_, _19081_, _07229_);
  or (_19321_, _19320_, _19319_);
  and (_19322_, _19321_, _11023_);
  and (_19323_, _19322_, _19318_);
  nor (_19325_, _11046_, _10788_);
  nor (_19326_, _19325_, _11047_);
  and (_19327_, _19326_, _11024_);
  or (_19328_, _19327_, _11026_);
  or (_19329_, _19328_, _19323_);
  or (_19330_, _11073_, _10615_);
  and (_19331_, _19330_, _11074_);
  or (_19332_, _19331_, _17490_);
  and (_19333_, _19332_, _19329_);
  or (_19334_, _19333_, _06892_);
  or (_19336_, _19331_, _17717_);
  and (_19337_, _19336_, _06523_);
  and (_19338_, _19337_, _19334_);
  or (_19339_, _19338_, _19077_);
  and (_19340_, _19339_, _11083_);
  or (_19341_, _11130_, _10857_);
  and (_19342_, _11131_, _11082_);
  and (_19343_, _19342_, _19341_);
  or (_19344_, _19343_, _11111_);
  or (_19345_, _19344_, _19340_);
  nand (_19347_, _11111_, _10152_);
  and (_19348_, _19347_, _11185_);
  and (_19349_, _19348_, _19345_);
  or (_19350_, _11176_, _11148_);
  nor (_19351_, _11185_, _11177_);
  and (_19352_, _19351_, _19350_);
  or (_19353_, _19352_, _11189_);
  or (_19354_, _19353_, _19349_);
  nor (_19355_, _11227_, _11198_);
  nor (_19356_, _19355_, _11228_);
  or (_19358_, _19356_, _17449_);
  and (_19359_, _19358_, _17448_);
  and (_19360_, _19359_, _19354_);
  and (_19361_, _19356_, _11188_);
  or (_19362_, _19361_, _19360_);
  and (_19363_, _19362_, _06293_);
  or (_19364_, _11265_, _11239_);
  and (_19365_, _19364_, _11266_);
  and (_19366_, _19365_, _06292_);
  or (_19367_, _19366_, _10474_);
  or (_19369_, _19367_, _19363_);
  nor (_19370_, _11304_, _11276_);
  nor (_19371_, _19370_, _11305_);
  or (_19372_, _19371_, _10475_);
  and (_19373_, _19372_, _12981_);
  and (_19374_, _19373_, _19369_);
  and (_19375_, _10472_, \oc8051_golden_model_1.ACC [5]);
  or (_19376_, _19375_, _06559_);
  or (_19377_, _19376_, _19374_);
  or (_19378_, _19118_, _07240_);
  and (_19380_, _19378_, _11316_);
  and (_19381_, _19380_, _19377_);
  nor (_19382_, _11324_, _10105_);
  or (_19383_, _19382_, _11325_);
  and (_19384_, _19383_, _11315_);
  or (_19385_, _19384_, _11320_);
  or (_19386_, _19385_, _19381_);
  nand (_19387_, _11320_, _08737_);
  and (_19388_, _19387_, _05933_);
  and (_19389_, _19388_, _19386_);
  and (_19391_, _19151_, _05932_);
  or (_19392_, _19391_, _06566_);
  or (_19393_, _19392_, _19389_);
  and (_19394_, _15695_, _07930_);
  or (_19395_, _19394_, _19081_);
  or (_19396_, _19395_, _06570_);
  and (_19397_, _19396_, _11339_);
  and (_19398_, _19397_, _19393_);
  nor (_19399_, _11350_, \oc8051_golden_model_1.ACC [6]);
  nor (_19400_, _19399_, _11351_);
  and (_19402_, _19400_, _11338_);
  or (_19403_, _19402_, _11345_);
  or (_19404_, _19403_, _19398_);
  nand (_19405_, _11345_, _08737_);
  and (_19406_, _19405_, _01320_);
  and (_19407_, _19406_, _19404_);
  or (_19408_, _19407_, _19074_);
  and (_42905_, _19408_, _42355_);
  not (_19409_, \oc8051_golden_model_1.PCON [0]);
  nor (_19410_, _01320_, _19409_);
  nand (_19412_, _11254_, _07942_);
  nor (_19413_, _07942_, _19409_);
  nor (_19414_, _19413_, _07217_);
  nand (_19415_, _19414_, _19412_);
  and (_19416_, _07942_, \oc8051_golden_model_1.ACC [0]);
  or (_19417_, _19416_, _19413_);
  and (_19418_, _19417_, _06345_);
  or (_19419_, _19418_, _06259_);
  nor (_19420_, _08374_, _11362_);
  or (_19421_, _19420_, _19413_);
  and (_19423_, _19421_, _06285_);
  nor (_19424_, _07143_, _19409_);
  and (_19425_, _19417_, _07143_);
  or (_19426_, _19425_, _19424_);
  and (_19427_, _19426_, _06286_);
  or (_19428_, _19427_, _06354_);
  or (_19429_, _19428_, _19423_);
  and (_19430_, _19429_, _06346_);
  or (_19431_, _19430_, _19419_);
  and (_19432_, _07942_, _07135_);
  nor (_19434_, _06259_, _06354_);
  or (_19435_, _19434_, _19413_);
  or (_19436_, _19435_, _19432_);
  and (_19437_, _19436_, _19431_);
  or (_19438_, _19437_, _09486_);
  and (_19439_, _09384_, _07942_);
  or (_19440_, _19413_, _06258_);
  or (_19441_, _19440_, _19439_);
  and (_19442_, _19441_, _19438_);
  or (_19443_, _19442_, _05972_);
  and (_19445_, _14413_, _07942_);
  or (_19446_, _19413_, _06251_);
  or (_19447_, _19446_, _19445_);
  and (_19448_, _19447_, _06216_);
  and (_19449_, _19448_, _19443_);
  and (_19450_, _07942_, _08929_);
  or (_19451_, _19450_, _19413_);
  and (_19452_, _19451_, _06215_);
  or (_19453_, _19452_, _06398_);
  or (_19454_, _19453_, _19449_);
  and (_19456_, _14311_, _07942_);
  or (_19457_, _19456_, _19413_);
  or (_19458_, _19457_, _09025_);
  and (_19459_, _19458_, _09030_);
  and (_19460_, _19459_, _19454_);
  nor (_19461_, _12532_, _11362_);
  or (_19462_, _19461_, _19413_);
  and (_19463_, _19412_, _06524_);
  and (_19464_, _19463_, _19462_);
  or (_19465_, _19464_, _19460_);
  and (_19467_, _19465_, _07219_);
  nand (_19468_, _19451_, _06426_);
  nor (_19469_, _19468_, _19420_);
  or (_19470_, _19469_, _06532_);
  or (_19471_, _19470_, _19467_);
  and (_19472_, _19471_, _19415_);
  or (_19473_, _19472_, _06437_);
  and (_19474_, _14307_, _07942_);
  or (_19475_, _19474_, _19413_);
  or (_19476_, _19475_, _07229_);
  and (_19478_, _19476_, _07231_);
  and (_19479_, _19478_, _19473_);
  not (_19480_, _06651_);
  and (_19481_, _19462_, _06535_);
  or (_19482_, _19481_, _19480_);
  or (_19483_, _19482_, _19479_);
  or (_19484_, _19421_, _06651_);
  and (_19485_, _19484_, _01320_);
  and (_19486_, _19485_, _19483_);
  or (_19487_, _19486_, _19410_);
  and (_42907_, _19487_, _42355_);
  not (_19489_, \oc8051_golden_model_1.PCON [1]);
  nor (_19490_, _07942_, _19489_);
  and (_19491_, _07942_, _09422_);
  or (_19492_, _19491_, _19490_);
  or (_19493_, _19492_, _06260_);
  or (_19494_, _07942_, \oc8051_golden_model_1.PCON [1]);
  and (_19495_, _14520_, _07942_);
  not (_19496_, _19495_);
  and (_19497_, _19496_, _19494_);
  or (_19499_, _19497_, _06286_);
  and (_19500_, _07942_, \oc8051_golden_model_1.ACC [1]);
  or (_19501_, _19500_, _19490_);
  and (_19502_, _19501_, _07143_);
  nor (_19503_, _07143_, _19489_);
  or (_19504_, _19503_, _06285_);
  or (_19505_, _19504_, _19502_);
  and (_19506_, _19505_, _07169_);
  and (_19507_, _19506_, _19499_);
  and (_19508_, _19492_, _06354_);
  or (_19510_, _19508_, _19507_);
  and (_19511_, _19510_, _06346_);
  and (_19512_, _19501_, _06345_);
  or (_19513_, _19512_, _06259_);
  or (_19514_, _19513_, _19511_);
  and (_19515_, _19514_, _19493_);
  or (_19516_, _19515_, _09486_);
  and (_19517_, _09339_, _07942_);
  or (_19518_, _19490_, _06258_);
  or (_19519_, _19518_, _19517_);
  and (_19521_, _19519_, _06251_);
  and (_19522_, _19521_, _19516_);
  or (_19523_, _14607_, _11362_);
  and (_19524_, _19494_, _05972_);
  and (_19525_, _19524_, _19523_);
  or (_19526_, _19525_, _19522_);
  and (_19527_, _19526_, _06399_);
  or (_19528_, _14505_, _11362_);
  and (_19529_, _19494_, _06398_);
  and (_19530_, _19529_, _19528_);
  nand (_19532_, _07942_, _07031_);
  and (_19533_, _19532_, _06215_);
  and (_19534_, _19533_, _19494_);
  or (_19535_, _19534_, _06524_);
  or (_19536_, _19535_, _19530_);
  or (_19537_, _19536_, _19527_);
  nor (_19538_, _11252_, _11362_);
  or (_19539_, _19538_, _19490_);
  nand (_19540_, _11251_, _07942_);
  and (_19541_, _19540_, _19539_);
  or (_19543_, _19541_, _09030_);
  and (_19544_, _19543_, _07219_);
  and (_19545_, _19544_, _19537_);
  or (_19546_, _14503_, _11362_);
  and (_19547_, _19494_, _06426_);
  and (_19548_, _19547_, _19546_);
  or (_19549_, _19548_, _06532_);
  or (_19550_, _19549_, _19545_);
  nor (_19551_, _19490_, _07217_);
  nand (_19552_, _19551_, _19540_);
  and (_19554_, _19552_, _07229_);
  and (_19555_, _19554_, _19550_);
  or (_19556_, _19532_, _08325_);
  and (_19557_, _19556_, _06437_);
  and (_19558_, _19557_, _19494_);
  or (_19559_, _19558_, _06535_);
  or (_19560_, _19559_, _19555_);
  or (_19561_, _19539_, _07231_);
  and (_19562_, _19561_, _19560_);
  or (_19563_, _19562_, _06559_);
  or (_19565_, _19497_, _07240_);
  and (_19566_, _19565_, _06570_);
  and (_19567_, _19566_, _19563_);
  or (_19568_, _19495_, _19490_);
  and (_19569_, _19568_, _06566_);
  or (_19570_, _19569_, _01324_);
  or (_19571_, _19570_, _19567_);
  or (_19572_, _01320_, \oc8051_golden_model_1.PCON [1]);
  and (_19573_, _19572_, _42355_);
  and (_42908_, _19573_, _19571_);
  not (_19575_, \oc8051_golden_model_1.PCON [2]);
  nor (_19576_, _01320_, _19575_);
  nor (_19577_, _07942_, _19575_);
  and (_19578_, _09293_, _07942_);
  or (_19579_, _19578_, _19577_);
  and (_19580_, _19579_, _09486_);
  and (_19581_, _14703_, _07942_);
  or (_19582_, _19581_, _19577_);
  or (_19583_, _19582_, _06286_);
  and (_19584_, _07942_, \oc8051_golden_model_1.ACC [2]);
  or (_19586_, _19584_, _19577_);
  and (_19587_, _19586_, _07143_);
  nor (_19588_, _07143_, _19575_);
  or (_19589_, _19588_, _06285_);
  or (_19590_, _19589_, _19587_);
  and (_19591_, _19590_, _07169_);
  and (_19592_, _19591_, _19583_);
  and (_19593_, _07942_, _08662_);
  or (_19594_, _19593_, _19577_);
  and (_19595_, _19594_, _06354_);
  or (_19597_, _19595_, _19592_);
  and (_19598_, _19597_, _06346_);
  and (_19599_, _19586_, _06345_);
  or (_19600_, _19599_, _06259_);
  or (_19601_, _19600_, _19598_);
  or (_19602_, _19594_, _06260_);
  and (_19603_, _19602_, _06258_);
  and (_19604_, _19603_, _19601_);
  or (_19605_, _19604_, _05972_);
  or (_19606_, _19605_, _19580_);
  and (_19608_, _14804_, _07942_);
  or (_19609_, _19577_, _06251_);
  or (_19610_, _19609_, _19608_);
  and (_19611_, _19610_, _06216_);
  and (_19612_, _19611_, _19606_);
  and (_19613_, _07942_, _08980_);
  or (_19614_, _19613_, _19577_);
  and (_19615_, _19614_, _06215_);
  or (_19616_, _19615_, _06398_);
  or (_19617_, _19616_, _19612_);
  and (_19619_, _14697_, _07942_);
  or (_19620_, _19619_, _19577_);
  or (_19621_, _19620_, _09025_);
  and (_19622_, _19621_, _09030_);
  and (_19623_, _19622_, _19617_);
  and (_19624_, _11250_, _07942_);
  or (_19625_, _19624_, _19577_);
  and (_19626_, _19625_, _06524_);
  or (_19627_, _19626_, _19623_);
  and (_19628_, _19627_, _07219_);
  or (_19630_, _19577_, _08424_);
  and (_19631_, _19614_, _06426_);
  and (_19632_, _19631_, _19630_);
  or (_19633_, _19632_, _19628_);
  and (_19634_, _19633_, _07217_);
  and (_19635_, _19586_, _06532_);
  and (_19636_, _19635_, _19630_);
  or (_19637_, _19636_, _06437_);
  or (_19638_, _19637_, _19634_);
  and (_19639_, _14694_, _07942_);
  or (_19641_, _19577_, _07229_);
  or (_19642_, _19641_, _19639_);
  and (_19643_, _19642_, _07231_);
  and (_19644_, _19643_, _19638_);
  nor (_19645_, _11249_, _11362_);
  or (_19646_, _19645_, _19577_);
  and (_19647_, _19646_, _06535_);
  or (_19648_, _19647_, _19644_);
  and (_19649_, _19648_, _07240_);
  and (_19650_, _19582_, _06559_);
  or (_19652_, _19650_, _06566_);
  or (_19653_, _19652_, _19649_);
  and (_19654_, _14873_, _07942_);
  or (_19655_, _19577_, _06570_);
  or (_19656_, _19655_, _19654_);
  and (_19657_, _19656_, _01320_);
  and (_19658_, _19657_, _19653_);
  or (_19659_, _19658_, _19576_);
  and (_42909_, _19659_, _42355_);
  and (_19660_, _11362_, \oc8051_golden_model_1.PCON [3]);
  and (_19662_, _14900_, _07942_);
  or (_19663_, _19662_, _19660_);
  or (_19664_, _19663_, _06286_);
  and (_19665_, _07942_, \oc8051_golden_model_1.ACC [3]);
  or (_19666_, _19665_, _19660_);
  and (_19667_, _19666_, _07143_);
  and (_19668_, _07144_, \oc8051_golden_model_1.PCON [3]);
  or (_19669_, _19668_, _06285_);
  or (_19670_, _19669_, _19667_);
  and (_19671_, _19670_, _07169_);
  and (_19673_, _19671_, _19664_);
  and (_19674_, _07942_, _09421_);
  or (_19675_, _19674_, _19660_);
  and (_19676_, _19675_, _06354_);
  or (_19677_, _19676_, _19673_);
  and (_19678_, _19677_, _06346_);
  and (_19679_, _19666_, _06345_);
  or (_19680_, _19679_, _06259_);
  or (_19681_, _19680_, _19678_);
  or (_19682_, _19675_, _06260_);
  and (_19684_, _19682_, _19681_);
  or (_19685_, _19684_, _09486_);
  and (_19686_, _09247_, _07942_);
  or (_19687_, _19660_, _06258_);
  or (_19688_, _19687_, _19686_);
  and (_19689_, _19688_, _06251_);
  and (_19690_, _19689_, _19685_);
  and (_19691_, _14998_, _07942_);
  or (_19692_, _19691_, _19660_);
  and (_19693_, _19692_, _05972_);
  or (_19695_, _19693_, _10080_);
  or (_19696_, _19695_, _19690_);
  and (_19697_, _14893_, _07942_);
  or (_19698_, _19660_, _09025_);
  or (_19699_, _19698_, _19697_);
  and (_19700_, _07942_, _08809_);
  or (_19701_, _19700_, _19660_);
  or (_19702_, _19701_, _06216_);
  and (_19703_, _19702_, _09030_);
  and (_19704_, _19703_, _19699_);
  and (_19706_, _19704_, _19696_);
  and (_19707_, _12529_, _07942_);
  or (_19708_, _19707_, _19660_);
  and (_19709_, _19708_, _06524_);
  or (_19710_, _19709_, _19706_);
  and (_19711_, _19710_, _07219_);
  or (_19712_, _19660_, _08280_);
  and (_19713_, _19701_, _06426_);
  and (_19714_, _19713_, _19712_);
  or (_19715_, _19714_, _19711_);
  and (_19717_, _19715_, _07217_);
  and (_19718_, _19666_, _06532_);
  and (_19719_, _19718_, _19712_);
  or (_19720_, _19719_, _06437_);
  or (_19721_, _19720_, _19717_);
  and (_19722_, _14890_, _07942_);
  or (_19723_, _19660_, _07229_);
  or (_19724_, _19723_, _19722_);
  and (_19725_, _19724_, _07231_);
  and (_19726_, _19725_, _19721_);
  nor (_19728_, _11247_, _11362_);
  or (_19729_, _19728_, _19660_);
  and (_19730_, _19729_, _06535_);
  or (_19731_, _19730_, _06559_);
  or (_19732_, _19731_, _19726_);
  or (_19733_, _19663_, _07240_);
  and (_19734_, _19733_, _06570_);
  and (_19735_, _19734_, _19732_);
  and (_19736_, _15068_, _07942_);
  or (_19737_, _19736_, _19660_);
  and (_19739_, _19737_, _06566_);
  or (_19740_, _19739_, _01324_);
  or (_19741_, _19740_, _19735_);
  or (_19742_, _01320_, \oc8051_golden_model_1.PCON [3]);
  and (_19743_, _19742_, _42355_);
  and (_42910_, _19743_, _19741_);
  and (_19744_, _11362_, \oc8051_golden_model_1.PCON [4]);
  and (_19745_, _15133_, _07942_);
  or (_19746_, _19745_, _19744_);
  or (_19747_, _19746_, _06286_);
  and (_19749_, _07942_, \oc8051_golden_model_1.ACC [4]);
  or (_19750_, _19749_, _19744_);
  and (_19751_, _19750_, _07143_);
  and (_19752_, _07144_, \oc8051_golden_model_1.PCON [4]);
  or (_19753_, _19752_, _06285_);
  or (_19754_, _19753_, _19751_);
  and (_19755_, _19754_, _07169_);
  and (_19756_, _19755_, _19747_);
  and (_19757_, _09420_, _07942_);
  or (_19758_, _19757_, _19744_);
  and (_19760_, _19758_, _06354_);
  or (_19761_, _19760_, _19756_);
  and (_19762_, _19761_, _06346_);
  and (_19763_, _19750_, _06345_);
  or (_19764_, _19763_, _06259_);
  or (_19765_, _19764_, _19762_);
  or (_19766_, _19758_, _06260_);
  and (_19767_, _19766_, _19765_);
  or (_19768_, _19767_, _09486_);
  and (_19769_, _09437_, _07942_);
  or (_19772_, _19744_, _06258_);
  or (_19773_, _19772_, _19769_);
  and (_19774_, _19773_, _06251_);
  and (_19775_, _19774_, _19768_);
  and (_19776_, _15226_, _07942_);
  or (_19777_, _19776_, _19744_);
  and (_19778_, _19777_, _05972_);
  or (_19779_, _19778_, _19775_);
  or (_19780_, _19779_, _10080_);
  and (_19781_, _15114_, _07942_);
  or (_19784_, _19744_, _09025_);
  or (_19785_, _19784_, _19781_);
  and (_19786_, _08919_, _07942_);
  or (_19787_, _19786_, _19744_);
  or (_19788_, _19787_, _06216_);
  and (_19789_, _19788_, _09030_);
  and (_19790_, _19789_, _19785_);
  and (_19791_, _19790_, _19780_);
  and (_19792_, _11245_, _07942_);
  or (_19793_, _19792_, _19744_);
  and (_19796_, _19793_, _06524_);
  or (_19797_, _19796_, _19791_);
  and (_19798_, _19797_, _07219_);
  or (_19799_, _19744_, _08528_);
  and (_19800_, _19787_, _06426_);
  and (_19801_, _19800_, _19799_);
  or (_19802_, _19801_, _19798_);
  and (_19803_, _19802_, _07217_);
  and (_19804_, _19750_, _06532_);
  and (_19805_, _19804_, _19799_);
  or (_19808_, _19805_, _06437_);
  or (_19809_, _19808_, _19803_);
  and (_19810_, _15111_, _07942_);
  or (_19811_, _19744_, _07229_);
  or (_19812_, _19811_, _19810_);
  and (_19813_, _19812_, _07231_);
  and (_19814_, _19813_, _19809_);
  nor (_19815_, _11244_, _11362_);
  or (_19816_, _19815_, _19744_);
  and (_19817_, _19816_, _06535_);
  or (_19820_, _19817_, _06559_);
  or (_19821_, _19820_, _19814_);
  or (_19822_, _19746_, _07240_);
  and (_19823_, _19822_, _06570_);
  and (_19824_, _19823_, _19821_);
  and (_19825_, _15296_, _07942_);
  or (_19826_, _19825_, _19744_);
  and (_19827_, _19826_, _06566_);
  or (_19828_, _19827_, _01324_);
  or (_19829_, _19828_, _19824_);
  or (_19832_, _01320_, \oc8051_golden_model_1.PCON [4]);
  and (_19833_, _19832_, _42355_);
  and (_42911_, _19833_, _19829_);
  and (_19834_, _11362_, \oc8051_golden_model_1.PCON [5]);
  and (_19835_, _15330_, _07942_);
  or (_19836_, _19835_, _19834_);
  or (_19837_, _19836_, _06286_);
  and (_19838_, _07942_, \oc8051_golden_model_1.ACC [5]);
  or (_19839_, _19838_, _19834_);
  and (_19840_, _19839_, _07143_);
  and (_19843_, _07144_, \oc8051_golden_model_1.PCON [5]);
  or (_19844_, _19843_, _06285_);
  or (_19845_, _19844_, _19840_);
  and (_19846_, _19845_, _07169_);
  and (_19847_, _19846_, _19837_);
  and (_19848_, _09419_, _07942_);
  or (_19849_, _19848_, _19834_);
  and (_19850_, _19849_, _06354_);
  or (_19851_, _19850_, _19847_);
  and (_19852_, _19851_, _06346_);
  and (_19854_, _19839_, _06345_);
  or (_19855_, _19854_, _06259_);
  or (_19856_, _19855_, _19852_);
  or (_19857_, _19849_, _06260_);
  and (_19858_, _19857_, _19856_);
  or (_19859_, _19858_, _09486_);
  and (_19860_, _09436_, _07942_);
  or (_19861_, _19834_, _06258_);
  or (_19862_, _19861_, _19860_);
  and (_19863_, _19862_, _06251_);
  and (_19865_, _19863_, _19859_);
  and (_19866_, _15421_, _07942_);
  or (_19867_, _19866_, _19834_);
  and (_19868_, _19867_, _05972_);
  or (_19869_, _19868_, _10080_);
  or (_19870_, _19869_, _19865_);
  and (_19871_, _15313_, _07942_);
  or (_19872_, _19834_, _09025_);
  or (_19873_, _19872_, _19871_);
  and (_19874_, _08913_, _07942_);
  or (_19876_, _19874_, _19834_);
  or (_19877_, _19876_, _06216_);
  and (_19878_, _19877_, _09030_);
  and (_19879_, _19878_, _19873_);
  and (_19880_, _19879_, _19870_);
  and (_19881_, _12536_, _07942_);
  or (_19882_, _19881_, _19834_);
  and (_19883_, _19882_, _06524_);
  or (_19884_, _19883_, _19880_);
  and (_19885_, _19884_, _07219_);
  or (_19887_, _19834_, _08231_);
  and (_19888_, _19876_, _06426_);
  and (_19889_, _19888_, _19887_);
  or (_19890_, _19889_, _19885_);
  and (_19891_, _19890_, _07217_);
  and (_19892_, _19839_, _06532_);
  and (_19893_, _19892_, _19887_);
  or (_19894_, _19893_, _06437_);
  or (_19895_, _19894_, _19891_);
  and (_19896_, _15310_, _07942_);
  or (_19898_, _19834_, _07229_);
  or (_19899_, _19898_, _19896_);
  and (_19900_, _19899_, _07231_);
  and (_19901_, _19900_, _19895_);
  nor (_19902_, _11241_, _11362_);
  or (_19903_, _19902_, _19834_);
  and (_19904_, _19903_, _06535_);
  or (_19905_, _19904_, _06559_);
  or (_19906_, _19905_, _19901_);
  or (_19907_, _19836_, _07240_);
  and (_19909_, _19907_, _06570_);
  and (_19910_, _19909_, _19906_);
  and (_19911_, _15493_, _07942_);
  or (_19912_, _19911_, _19834_);
  and (_19913_, _19912_, _06566_);
  or (_19914_, _19913_, _01324_);
  or (_19915_, _19914_, _19910_);
  or (_19916_, _01320_, \oc8051_golden_model_1.PCON [5]);
  and (_19917_, _19916_, _42355_);
  and (_42912_, _19917_, _19915_);
  and (_19919_, _11362_, \oc8051_golden_model_1.PCON [6]);
  and (_19920_, _15521_, _07942_);
  or (_19921_, _19920_, _19919_);
  or (_19922_, _19921_, _06286_);
  and (_19923_, _07942_, \oc8051_golden_model_1.ACC [6]);
  or (_19924_, _19923_, _19919_);
  and (_19925_, _19924_, _07143_);
  and (_19926_, _07144_, \oc8051_golden_model_1.PCON [6]);
  or (_19927_, _19926_, _06285_);
  or (_19928_, _19927_, _19925_);
  and (_19930_, _19928_, _07169_);
  and (_19931_, _19930_, _19922_);
  and (_19932_, _09418_, _07942_);
  or (_19933_, _19932_, _19919_);
  and (_19934_, _19933_, _06354_);
  or (_19935_, _19934_, _19931_);
  and (_19936_, _19935_, _06346_);
  and (_19937_, _19924_, _06345_);
  or (_19938_, _19937_, _06259_);
  or (_19939_, _19938_, _19936_);
  or (_19941_, _19933_, _06260_);
  and (_19942_, _19941_, _19939_);
  or (_19943_, _19942_, _09486_);
  and (_19944_, _09435_, _07942_);
  or (_19945_, _19919_, _06258_);
  or (_19946_, _19945_, _19944_);
  and (_19947_, _19946_, _06251_);
  and (_19948_, _19947_, _19943_);
  and (_19949_, _15623_, _07942_);
  or (_19950_, _19949_, _19919_);
  and (_19952_, _19950_, _05972_);
  or (_19953_, _19952_, _10080_);
  or (_19954_, _19953_, _19948_);
  and (_19955_, _15517_, _07942_);
  or (_19956_, _19919_, _09025_);
  or (_19957_, _19956_, _19955_);
  and (_19958_, _08845_, _07942_);
  or (_19959_, _19958_, _19919_);
  or (_19960_, _19959_, _06216_);
  and (_19961_, _19960_, _09030_);
  and (_19963_, _19961_, _19957_);
  and (_19964_, _19963_, _19954_);
  and (_19965_, _11239_, _07942_);
  or (_19966_, _19965_, _19919_);
  and (_19967_, _19966_, _06524_);
  or (_19968_, _19967_, _19964_);
  and (_19969_, _19968_, _07219_);
  or (_19970_, _19919_, _08128_);
  and (_19971_, _19959_, _06426_);
  and (_19972_, _19971_, _19970_);
  or (_19974_, _19972_, _19969_);
  and (_19975_, _19974_, _07217_);
  and (_19976_, _19924_, _06532_);
  and (_19977_, _19976_, _19970_);
  or (_19978_, _19977_, _06437_);
  or (_19979_, _19978_, _19975_);
  and (_19980_, _15514_, _07942_);
  or (_19981_, _19919_, _07229_);
  or (_19982_, _19981_, _19980_);
  and (_19983_, _19982_, _07231_);
  and (_19985_, _19983_, _19979_);
  nor (_19986_, _11238_, _11362_);
  or (_19987_, _19986_, _19919_);
  and (_19988_, _19987_, _06535_);
  or (_19989_, _19988_, _06559_);
  or (_19990_, _19989_, _19985_);
  or (_19991_, _19921_, _07240_);
  and (_19992_, _19991_, _06570_);
  and (_19993_, _19992_, _19990_);
  and (_19994_, _15695_, _07942_);
  or (_19996_, _19994_, _19919_);
  and (_19997_, _19996_, _06566_);
  or (_19998_, _19997_, _01324_);
  or (_19999_, _19998_, _19993_);
  or (_20000_, _01320_, \oc8051_golden_model_1.PCON [6]);
  and (_20001_, _20000_, _42355_);
  and (_42913_, _20001_, _19999_);
  not (_20002_, \oc8051_golden_model_1.TMOD [0]);
  nor (_20003_, _01320_, _20002_);
  nand (_20004_, _11254_, _07904_);
  nor (_20006_, _07904_, _20002_);
  nor (_20007_, _20006_, _07217_);
  nand (_20008_, _20007_, _20004_);
  and (_20009_, _07904_, _07135_);
  or (_20010_, _20009_, _20006_);
  or (_20011_, _20010_, _06260_);
  nor (_20012_, _08374_, _11439_);
  or (_20013_, _20012_, _20006_);
  or (_20014_, _20013_, _06286_);
  and (_20015_, _07904_, \oc8051_golden_model_1.ACC [0]);
  or (_20017_, _20015_, _20006_);
  and (_20018_, _20017_, _07143_);
  nor (_20019_, _07143_, _20002_);
  or (_20020_, _20019_, _06285_);
  or (_20021_, _20020_, _20018_);
  and (_20022_, _20021_, _07169_);
  and (_20023_, _20022_, _20014_);
  and (_20024_, _20010_, _06354_);
  or (_20025_, _20024_, _20023_);
  and (_20026_, _20025_, _06346_);
  and (_20028_, _20017_, _06345_);
  or (_20029_, _20028_, _06259_);
  or (_20030_, _20029_, _20026_);
  and (_20031_, _20030_, _20011_);
  or (_20032_, _20031_, _09486_);
  and (_20033_, _09384_, _07904_);
  or (_20034_, _20006_, _06258_);
  or (_20035_, _20034_, _20033_);
  and (_20036_, _20035_, _20032_);
  or (_20037_, _20036_, _05972_);
  and (_20039_, _14413_, _07904_);
  or (_20040_, _20006_, _06251_);
  or (_20041_, _20040_, _20039_);
  and (_20042_, _20041_, _06216_);
  and (_20043_, _20042_, _20037_);
  and (_20044_, _07904_, _08929_);
  or (_20045_, _20044_, _20006_);
  and (_20046_, _20045_, _06215_);
  or (_20047_, _20046_, _06398_);
  or (_20048_, _20047_, _20043_);
  and (_20050_, _14311_, _07904_);
  or (_20051_, _20050_, _20006_);
  or (_20052_, _20051_, _09025_);
  and (_20053_, _20052_, _09030_);
  and (_20054_, _20053_, _20048_);
  nor (_20055_, _12532_, _11439_);
  or (_20056_, _20055_, _20006_);
  and (_20057_, _20004_, _06524_);
  and (_20058_, _20057_, _20056_);
  or (_20059_, _20058_, _20054_);
  and (_20061_, _20059_, _07219_);
  nand (_20062_, _20045_, _06426_);
  nor (_20063_, _20062_, _20012_);
  or (_20064_, _20063_, _06532_);
  or (_20065_, _20064_, _20061_);
  and (_20066_, _20065_, _20008_);
  or (_20067_, _20066_, _06437_);
  and (_20068_, _14307_, _07904_);
  or (_20069_, _20006_, _07229_);
  or (_20070_, _20069_, _20068_);
  and (_20072_, _20070_, _07231_);
  and (_20073_, _20072_, _20067_);
  and (_20074_, _20056_, _06535_);
  or (_20075_, _20074_, _19480_);
  or (_20076_, _20075_, _20073_);
  or (_20077_, _20013_, _06651_);
  and (_20078_, _20077_, _01320_);
  and (_20079_, _20078_, _20076_);
  or (_20080_, _20079_, _20003_);
  and (_42915_, _20080_, _42355_);
  and (_20082_, _11439_, \oc8051_golden_model_1.TMOD [1]);
  nor (_20083_, _11252_, _11439_);
  or (_20084_, _20083_, _20082_);
  or (_20085_, _20084_, _07231_);
  or (_20086_, _07904_, \oc8051_golden_model_1.TMOD [1]);
  and (_20087_, _14520_, _07904_);
  not (_20088_, _20087_);
  and (_20089_, _20088_, _20086_);
  or (_20090_, _20089_, _06286_);
  and (_20091_, _07904_, \oc8051_golden_model_1.ACC [1]);
  or (_20093_, _20091_, _20082_);
  and (_20094_, _20093_, _07143_);
  and (_20095_, _07144_, \oc8051_golden_model_1.TMOD [1]);
  or (_20096_, _20095_, _06285_);
  or (_20097_, _20096_, _20094_);
  and (_20098_, _20097_, _07169_);
  and (_20099_, _20098_, _20090_);
  and (_20100_, _07904_, _09422_);
  or (_20101_, _20100_, _20082_);
  and (_20102_, _20101_, _06354_);
  or (_20104_, _20102_, _20099_);
  and (_20105_, _20104_, _06346_);
  and (_20106_, _20093_, _06345_);
  or (_20107_, _20106_, _06259_);
  or (_20108_, _20107_, _20105_);
  or (_20109_, _20101_, _06260_);
  and (_20110_, _20109_, _20108_);
  or (_20111_, _20110_, _09486_);
  and (_20112_, _09339_, _07904_);
  or (_20113_, _20082_, _06258_);
  or (_20115_, _20113_, _20112_);
  and (_20116_, _20115_, _06251_);
  and (_20117_, _20116_, _20111_);
  or (_20118_, _14607_, _11439_);
  and (_20119_, _20086_, _05972_);
  and (_20120_, _20119_, _20118_);
  or (_20121_, _20120_, _20117_);
  and (_20122_, _20121_, _06399_);
  or (_20123_, _14505_, _11439_);
  and (_20124_, _20123_, _06398_);
  nand (_20126_, _07904_, _07031_);
  and (_20127_, _20126_, _06215_);
  or (_20128_, _20127_, _20124_);
  and (_20129_, _20128_, _20086_);
  or (_20130_, _20129_, _06524_);
  or (_20131_, _20130_, _20122_);
  and (_20132_, _11253_, _07904_);
  or (_20133_, _20132_, _20082_);
  or (_20134_, _20133_, _09030_);
  and (_20135_, _20134_, _07219_);
  and (_20137_, _20135_, _20131_);
  or (_20138_, _14503_, _11439_);
  and (_20139_, _20086_, _06426_);
  and (_20140_, _20139_, _20138_);
  or (_20141_, _20140_, _06532_);
  or (_20142_, _20141_, _20137_);
  and (_20143_, _20091_, _08325_);
  or (_20144_, _20082_, _07217_);
  or (_20145_, _20144_, _20143_);
  and (_20146_, _20145_, _07229_);
  and (_20148_, _20146_, _20142_);
  or (_20149_, _20126_, _08325_);
  and (_20150_, _20086_, _06437_);
  and (_20151_, _20150_, _20149_);
  or (_20152_, _20151_, _06535_);
  or (_20153_, _20152_, _20148_);
  and (_20154_, _20153_, _20085_);
  or (_20155_, _20154_, _06559_);
  or (_20156_, _20089_, _07240_);
  and (_20157_, _20156_, _06570_);
  and (_20159_, _20157_, _20155_);
  or (_20160_, _20087_, _20082_);
  and (_20161_, _20160_, _06566_);
  or (_20162_, _20161_, _01324_);
  or (_20163_, _20162_, _20159_);
  or (_20164_, _01320_, \oc8051_golden_model_1.TMOD [1]);
  and (_20165_, _20164_, _42355_);
  and (_42916_, _20165_, _20163_);
  and (_20166_, _01324_, \oc8051_golden_model_1.TMOD [2]);
  and (_20167_, _11439_, \oc8051_golden_model_1.TMOD [2]);
  and (_20169_, _09293_, _07904_);
  or (_20170_, _20169_, _20167_);
  and (_20171_, _20170_, _09486_);
  and (_20172_, _14703_, _07904_);
  or (_20173_, _20172_, _20167_);
  or (_20174_, _20173_, _06286_);
  and (_20175_, _07904_, \oc8051_golden_model_1.ACC [2]);
  or (_20176_, _20175_, _20167_);
  and (_20177_, _20176_, _07143_);
  and (_20178_, _07144_, \oc8051_golden_model_1.TMOD [2]);
  or (_20180_, _20178_, _06285_);
  or (_20181_, _20180_, _20177_);
  and (_20182_, _20181_, _07169_);
  and (_20183_, _20182_, _20174_);
  and (_20184_, _07904_, _08662_);
  or (_20185_, _20184_, _20167_);
  and (_20186_, _20185_, _06354_);
  or (_20187_, _20186_, _20183_);
  and (_20188_, _20187_, _06346_);
  and (_20189_, _20176_, _06345_);
  or (_20191_, _20189_, _06259_);
  or (_20192_, _20191_, _20188_);
  or (_20193_, _20185_, _06260_);
  and (_20194_, _20193_, _06258_);
  and (_20195_, _20194_, _20192_);
  or (_20196_, _20195_, _05972_);
  or (_20197_, _20196_, _20171_);
  and (_20198_, _14804_, _07904_);
  or (_20199_, _20167_, _06251_);
  or (_20200_, _20199_, _20198_);
  and (_20202_, _20200_, _06216_);
  and (_20203_, _20202_, _20197_);
  and (_20204_, _07904_, _08980_);
  or (_20205_, _20204_, _20167_);
  and (_20206_, _20205_, _06215_);
  or (_20207_, _20206_, _06398_);
  or (_20208_, _20207_, _20203_);
  and (_20209_, _14697_, _07904_);
  or (_20210_, _20209_, _20167_);
  or (_20211_, _20210_, _09025_);
  and (_20213_, _20211_, _09030_);
  and (_20214_, _20213_, _20208_);
  and (_20215_, _11250_, _07904_);
  or (_20216_, _20215_, _20167_);
  and (_20217_, _20216_, _06524_);
  or (_20218_, _20217_, _20214_);
  and (_20219_, _20218_, _07219_);
  or (_20220_, _20167_, _08424_);
  and (_20221_, _20205_, _06426_);
  and (_20222_, _20221_, _20220_);
  or (_20224_, _20222_, _20219_);
  and (_20225_, _20224_, _07217_);
  and (_20226_, _20176_, _06532_);
  and (_20227_, _20226_, _20220_);
  or (_20228_, _20227_, _06437_);
  or (_20229_, _20228_, _20225_);
  and (_20230_, _14694_, _07904_);
  or (_20231_, _20167_, _07229_);
  or (_20232_, _20231_, _20230_);
  and (_20233_, _20232_, _07231_);
  and (_20235_, _20233_, _20229_);
  nor (_20236_, _11249_, _11439_);
  or (_20237_, _20236_, _20167_);
  and (_20238_, _20237_, _06535_);
  or (_20239_, _20238_, _20235_);
  and (_20240_, _20239_, _07240_);
  and (_20241_, _20173_, _06559_);
  or (_20242_, _20241_, _06566_);
  or (_20243_, _20242_, _20240_);
  and (_20244_, _14873_, _07904_);
  or (_20246_, _20167_, _06570_);
  or (_20247_, _20246_, _20244_);
  and (_20248_, _20247_, _01320_);
  and (_20249_, _20248_, _20243_);
  or (_20250_, _20249_, _20166_);
  and (_42917_, _20250_, _42355_);
  and (_20251_, _11439_, \oc8051_golden_model_1.TMOD [3]);
  and (_20252_, _14900_, _07904_);
  or (_20253_, _20252_, _20251_);
  or (_20254_, _20253_, _06286_);
  and (_20256_, _07904_, \oc8051_golden_model_1.ACC [3]);
  or (_20257_, _20256_, _20251_);
  and (_20258_, _20257_, _07143_);
  and (_20259_, _07144_, \oc8051_golden_model_1.TMOD [3]);
  or (_20260_, _20259_, _06285_);
  or (_20261_, _20260_, _20258_);
  and (_20262_, _20261_, _07169_);
  and (_20263_, _20262_, _20254_);
  and (_20264_, _07904_, _09421_);
  or (_20265_, _20264_, _20251_);
  and (_20267_, _20265_, _06354_);
  or (_20268_, _20267_, _20263_);
  and (_20269_, _20268_, _06346_);
  and (_20270_, _20257_, _06345_);
  or (_20271_, _20270_, _06259_);
  or (_20272_, _20271_, _20269_);
  or (_20273_, _20265_, _06260_);
  and (_20274_, _20273_, _20272_);
  or (_20275_, _20274_, _09486_);
  and (_20276_, _09247_, _07904_);
  or (_20278_, _20251_, _06258_);
  or (_20279_, _20278_, _20276_);
  and (_20280_, _20279_, _06251_);
  and (_20281_, _20280_, _20275_);
  and (_20282_, _14998_, _07904_);
  or (_20283_, _20282_, _20251_);
  and (_20284_, _20283_, _05972_);
  or (_20285_, _20284_, _10080_);
  or (_20286_, _20285_, _20281_);
  and (_20287_, _14893_, _07904_);
  or (_20289_, _20251_, _09025_);
  or (_20290_, _20289_, _20287_);
  and (_20291_, _07904_, _08809_);
  or (_20292_, _20291_, _20251_);
  or (_20293_, _20292_, _06216_);
  and (_20294_, _20293_, _09030_);
  and (_20295_, _20294_, _20290_);
  and (_20296_, _20295_, _20286_);
  and (_20297_, _12529_, _07904_);
  or (_20298_, _20297_, _20251_);
  and (_20300_, _20298_, _06524_);
  or (_20301_, _20300_, _20296_);
  and (_20302_, _20301_, _07219_);
  or (_20303_, _20251_, _08280_);
  and (_20304_, _20292_, _06426_);
  and (_20305_, _20304_, _20303_);
  or (_20306_, _20305_, _20302_);
  and (_20307_, _20306_, _07217_);
  and (_20308_, _20257_, _06532_);
  and (_20309_, _20308_, _20303_);
  or (_20311_, _20309_, _06437_);
  or (_20312_, _20311_, _20307_);
  and (_20313_, _14890_, _07904_);
  or (_20314_, _20251_, _07229_);
  or (_20315_, _20314_, _20313_);
  and (_20316_, _20315_, _07231_);
  and (_20317_, _20316_, _20312_);
  nor (_20318_, _11247_, _11439_);
  or (_20319_, _20318_, _20251_);
  and (_20320_, _20319_, _06535_);
  or (_20322_, _20320_, _06559_);
  or (_20323_, _20322_, _20317_);
  or (_20324_, _20253_, _07240_);
  and (_20325_, _20324_, _06570_);
  and (_20326_, _20325_, _20323_);
  and (_20327_, _15068_, _07904_);
  or (_20328_, _20327_, _20251_);
  and (_20329_, _20328_, _06566_);
  or (_20330_, _20329_, _01324_);
  or (_20331_, _20330_, _20326_);
  or (_20333_, _01320_, \oc8051_golden_model_1.TMOD [3]);
  and (_20334_, _20333_, _42355_);
  and (_42919_, _20334_, _20331_);
  and (_20335_, _11439_, \oc8051_golden_model_1.TMOD [4]);
  and (_20336_, _09420_, _07904_);
  or (_20337_, _20336_, _20335_);
  or (_20338_, _20337_, _06260_);
  and (_20339_, _15133_, _07904_);
  or (_20340_, _20339_, _20335_);
  or (_20341_, _20340_, _06286_);
  and (_20343_, _07904_, \oc8051_golden_model_1.ACC [4]);
  or (_20344_, _20343_, _20335_);
  and (_20345_, _20344_, _07143_);
  and (_20346_, _07144_, \oc8051_golden_model_1.TMOD [4]);
  or (_20347_, _20346_, _06285_);
  or (_20348_, _20347_, _20345_);
  and (_20349_, _20348_, _07169_);
  and (_20350_, _20349_, _20341_);
  and (_20351_, _20337_, _06354_);
  or (_20352_, _20351_, _20350_);
  and (_20354_, _20352_, _06346_);
  and (_20355_, _20344_, _06345_);
  or (_20356_, _20355_, _06259_);
  or (_20357_, _20356_, _20354_);
  and (_20358_, _20357_, _20338_);
  or (_20359_, _20358_, _09486_);
  and (_20360_, _09437_, _07904_);
  or (_20361_, _20335_, _06258_);
  or (_20362_, _20361_, _20360_);
  and (_20363_, _20362_, _06251_);
  and (_20365_, _20363_, _20359_);
  and (_20366_, _15226_, _07904_);
  or (_20367_, _20366_, _20335_);
  and (_20368_, _20367_, _05972_);
  or (_20369_, _20368_, _20365_);
  or (_20370_, _20369_, _10080_);
  and (_20371_, _15114_, _07904_);
  or (_20372_, _20335_, _09025_);
  or (_20373_, _20372_, _20371_);
  and (_20374_, _08919_, _07904_);
  or (_20376_, _20374_, _20335_);
  or (_20377_, _20376_, _06216_);
  and (_20378_, _20377_, _09030_);
  and (_20379_, _20378_, _20373_);
  and (_20380_, _20379_, _20370_);
  and (_20381_, _11245_, _07904_);
  or (_20382_, _20381_, _20335_);
  and (_20383_, _20382_, _06524_);
  or (_20384_, _20383_, _20380_);
  and (_20385_, _20384_, _07219_);
  or (_20387_, _20335_, _08528_);
  and (_20388_, _20376_, _06426_);
  and (_20389_, _20388_, _20387_);
  or (_20390_, _20389_, _20385_);
  and (_20391_, _20390_, _07217_);
  and (_20392_, _20344_, _06532_);
  and (_20393_, _20392_, _20387_);
  or (_20394_, _20393_, _06437_);
  or (_20395_, _20394_, _20391_);
  and (_20396_, _15111_, _07904_);
  or (_20398_, _20335_, _07229_);
  or (_20399_, _20398_, _20396_);
  and (_20400_, _20399_, _07231_);
  and (_20401_, _20400_, _20395_);
  nor (_20402_, _11244_, _11439_);
  or (_20403_, _20402_, _20335_);
  and (_20404_, _20403_, _06535_);
  or (_20405_, _20404_, _06559_);
  or (_20406_, _20405_, _20401_);
  or (_20407_, _20340_, _07240_);
  and (_20409_, _20407_, _06570_);
  and (_20410_, _20409_, _20406_);
  and (_20411_, _15296_, _07904_);
  or (_20412_, _20411_, _20335_);
  and (_20413_, _20412_, _06566_);
  or (_20414_, _20413_, _01324_);
  or (_20415_, _20414_, _20410_);
  or (_20416_, _01320_, \oc8051_golden_model_1.TMOD [4]);
  and (_20417_, _20416_, _42355_);
  and (_42920_, _20417_, _20415_);
  and (_20419_, _11439_, \oc8051_golden_model_1.TMOD [5]);
  and (_20420_, _15330_, _07904_);
  or (_20421_, _20420_, _20419_);
  or (_20422_, _20421_, _06286_);
  and (_20423_, _07904_, \oc8051_golden_model_1.ACC [5]);
  or (_20424_, _20423_, _20419_);
  and (_20425_, _20424_, _07143_);
  and (_20426_, _07144_, \oc8051_golden_model_1.TMOD [5]);
  or (_20427_, _20426_, _06285_);
  or (_20428_, _20427_, _20425_);
  and (_20430_, _20428_, _07169_);
  and (_20431_, _20430_, _20422_);
  and (_20432_, _09419_, _07904_);
  or (_20433_, _20432_, _20419_);
  and (_20434_, _20433_, _06354_);
  or (_20435_, _20434_, _20431_);
  and (_20436_, _20435_, _06346_);
  and (_20437_, _20424_, _06345_);
  or (_20438_, _20437_, _06259_);
  or (_20439_, _20438_, _20436_);
  or (_20441_, _20433_, _06260_);
  and (_20442_, _20441_, _20439_);
  or (_20443_, _20442_, _09486_);
  and (_20444_, _09436_, _07904_);
  or (_20445_, _20419_, _06258_);
  or (_20446_, _20445_, _20444_);
  and (_20447_, _20446_, _06251_);
  and (_20448_, _20447_, _20443_);
  and (_20449_, _15421_, _07904_);
  or (_20450_, _20449_, _20419_);
  and (_20452_, _20450_, _05972_);
  or (_20453_, _20452_, _10080_);
  or (_20454_, _20453_, _20448_);
  and (_20455_, _15313_, _07904_);
  or (_20456_, _20419_, _09025_);
  or (_20457_, _20456_, _20455_);
  and (_20458_, _08913_, _07904_);
  or (_20459_, _20458_, _20419_);
  or (_20460_, _20459_, _06216_);
  and (_20461_, _20460_, _09030_);
  and (_20463_, _20461_, _20457_);
  and (_20464_, _20463_, _20454_);
  and (_20465_, _12536_, _07904_);
  or (_20466_, _20465_, _20419_);
  and (_20467_, _20466_, _06524_);
  or (_20468_, _20467_, _20464_);
  and (_20469_, _20468_, _07219_);
  or (_20470_, _20419_, _08231_);
  and (_20471_, _20459_, _06426_);
  and (_20472_, _20471_, _20470_);
  or (_20474_, _20472_, _20469_);
  and (_20475_, _20474_, _07217_);
  and (_20476_, _20424_, _06532_);
  and (_20477_, _20476_, _20470_);
  or (_20478_, _20477_, _06437_);
  or (_20479_, _20478_, _20475_);
  and (_20480_, _15310_, _07904_);
  or (_20481_, _20419_, _07229_);
  or (_20482_, _20481_, _20480_);
  and (_20483_, _20482_, _07231_);
  and (_20485_, _20483_, _20479_);
  nor (_20486_, _11241_, _11439_);
  or (_20487_, _20486_, _20419_);
  and (_20488_, _20487_, _06535_);
  or (_20489_, _20488_, _06559_);
  or (_20490_, _20489_, _20485_);
  or (_20491_, _20421_, _07240_);
  and (_20492_, _20491_, _06570_);
  and (_20493_, _20492_, _20490_);
  and (_20494_, _15493_, _07904_);
  or (_20496_, _20494_, _20419_);
  and (_20497_, _20496_, _06566_);
  or (_20498_, _20497_, _01324_);
  or (_20499_, _20498_, _20493_);
  or (_20500_, _01320_, \oc8051_golden_model_1.TMOD [5]);
  and (_20501_, _20500_, _42355_);
  and (_42921_, _20501_, _20499_);
  and (_20502_, _11439_, \oc8051_golden_model_1.TMOD [6]);
  and (_20503_, _15521_, _07904_);
  or (_20504_, _20503_, _20502_);
  or (_20506_, _20504_, _06286_);
  and (_20507_, _07904_, \oc8051_golden_model_1.ACC [6]);
  or (_20508_, _20507_, _20502_);
  and (_20509_, _20508_, _07143_);
  and (_20510_, _07144_, \oc8051_golden_model_1.TMOD [6]);
  or (_20511_, _20510_, _06285_);
  or (_20512_, _20511_, _20509_);
  and (_20513_, _20512_, _07169_);
  and (_20514_, _20513_, _20506_);
  and (_20515_, _09418_, _07904_);
  or (_20517_, _20515_, _20502_);
  and (_20518_, _20517_, _06354_);
  or (_20519_, _20518_, _20514_);
  and (_20520_, _20519_, _06346_);
  and (_20521_, _20508_, _06345_);
  or (_20522_, _20521_, _06259_);
  or (_20523_, _20522_, _20520_);
  or (_20524_, _20517_, _06260_);
  and (_20525_, _20524_, _20523_);
  or (_20526_, _20525_, _09486_);
  and (_20528_, _09435_, _07904_);
  or (_20529_, _20502_, _06258_);
  or (_20530_, _20529_, _20528_);
  and (_20531_, _20530_, _06251_);
  and (_20532_, _20531_, _20526_);
  and (_20533_, _15623_, _07904_);
  or (_20534_, _20533_, _20502_);
  and (_20535_, _20534_, _05972_);
  or (_20536_, _20535_, _10080_);
  or (_20537_, _20536_, _20532_);
  and (_20539_, _15517_, _07904_);
  or (_20540_, _20502_, _09025_);
  or (_20541_, _20540_, _20539_);
  and (_20542_, _08845_, _07904_);
  or (_20543_, _20542_, _20502_);
  or (_20544_, _20543_, _06216_);
  and (_20545_, _20544_, _09030_);
  and (_20546_, _20545_, _20541_);
  and (_20547_, _20546_, _20537_);
  and (_20548_, _11239_, _07904_);
  or (_20550_, _20548_, _20502_);
  and (_20551_, _20550_, _06524_);
  or (_20552_, _20551_, _20547_);
  and (_20553_, _20552_, _07219_);
  or (_20554_, _20502_, _08128_);
  and (_20555_, _20543_, _06426_);
  and (_20556_, _20555_, _20554_);
  or (_20557_, _20556_, _20553_);
  and (_20558_, _20557_, _07217_);
  and (_20559_, _20508_, _06532_);
  and (_20561_, _20559_, _20554_);
  or (_20562_, _20561_, _06437_);
  or (_20563_, _20562_, _20558_);
  and (_20564_, _15514_, _07904_);
  or (_20565_, _20502_, _07229_);
  or (_20566_, _20565_, _20564_);
  and (_20567_, _20566_, _07231_);
  and (_20568_, _20567_, _20563_);
  nor (_20569_, _11238_, _11439_);
  or (_20570_, _20569_, _20502_);
  and (_20572_, _20570_, _06535_);
  or (_20573_, _20572_, _06559_);
  or (_20574_, _20573_, _20568_);
  or (_20575_, _20504_, _07240_);
  and (_20576_, _20575_, _06570_);
  and (_20577_, _20576_, _20574_);
  and (_20578_, _15695_, _07904_);
  or (_20579_, _20578_, _20502_);
  and (_20580_, _20579_, _06566_);
  or (_20581_, _20580_, _01324_);
  or (_20583_, _20581_, _20577_);
  or (_20584_, _01320_, \oc8051_golden_model_1.TMOD [6]);
  and (_20585_, _20584_, _42355_);
  and (_42922_, _20585_, _20583_);
  not (_20586_, \oc8051_golden_model_1.DPL [0]);
  nor (_20587_, _01320_, _20586_);
  and (_20588_, _07950_, \oc8051_golden_model_1.ACC [0]);
  and (_20589_, _20588_, _08374_);
  nor (_20590_, _07950_, _20586_);
  or (_20591_, _20590_, _07217_);
  or (_20593_, _20591_, _20589_);
  and (_20594_, _09384_, _07950_);
  or (_20595_, _20594_, _20590_);
  and (_20596_, _20595_, _09486_);
  and (_20597_, _07950_, _07135_);
  or (_20598_, _20597_, _20590_);
  or (_20599_, _20598_, _07169_);
  nor (_20600_, _08374_, _11595_);
  or (_20601_, _20600_, _20590_);
  and (_20602_, _20601_, _06285_);
  nor (_20604_, _07143_, _20586_);
  or (_20605_, _20590_, _20588_);
  and (_20606_, _20605_, _07143_);
  or (_20607_, _20606_, _20604_);
  and (_20608_, _20607_, _06286_);
  or (_20609_, _20608_, _06354_);
  or (_20610_, _20609_, _20602_);
  and (_20611_, _20610_, _20599_);
  or (_20612_, _20611_, _06345_);
  or (_20613_, _20605_, _06346_);
  and (_20615_, _20613_, _11536_);
  and (_20616_, _20615_, _20612_);
  and (_20617_, _11535_, _20586_);
  or (_20618_, _20617_, _20616_);
  and (_20619_, _20618_, _06396_);
  nor (_20620_, _06850_, _06396_);
  or (_20621_, _20620_, _06259_);
  or (_20622_, _20621_, _20619_);
  or (_20623_, _20598_, _06260_);
  and (_20624_, _20623_, _06258_);
  and (_20626_, _20624_, _20622_);
  or (_20627_, _20626_, _05972_);
  or (_20628_, _20627_, _20596_);
  and (_20629_, _14413_, _07950_);
  or (_20630_, _20590_, _06251_);
  or (_20631_, _20630_, _20629_);
  and (_20632_, _20631_, _06216_);
  and (_20633_, _20632_, _20628_);
  and (_20634_, _07950_, _08929_);
  or (_20635_, _20634_, _20590_);
  and (_20637_, _20635_, _06215_);
  or (_20638_, _20637_, _06398_);
  or (_20639_, _20638_, _20633_);
  and (_20640_, _14311_, _07950_);
  or (_20641_, _20640_, _20590_);
  or (_20642_, _20641_, _09025_);
  and (_20643_, _20642_, _09030_);
  and (_20644_, _20643_, _20639_);
  nor (_20645_, _12532_, _11595_);
  or (_20646_, _20645_, _20590_);
  nor (_20648_, _20589_, _09030_);
  and (_20649_, _20648_, _20646_);
  or (_20650_, _20649_, _20644_);
  and (_20651_, _20650_, _07219_);
  nand (_20652_, _20635_, _06426_);
  nor (_20653_, _20652_, _20600_);
  or (_20654_, _20653_, _06532_);
  or (_20655_, _20654_, _20651_);
  and (_20656_, _20655_, _20593_);
  or (_20657_, _20656_, _06437_);
  and (_20659_, _14307_, _07950_);
  or (_20660_, _20659_, _20590_);
  or (_20661_, _20660_, _07229_);
  and (_20662_, _20661_, _07231_);
  and (_20663_, _20662_, _20657_);
  and (_20664_, _20646_, _06535_);
  or (_20665_, _20664_, _19480_);
  or (_20666_, _20665_, _20663_);
  or (_20667_, _20601_, _06651_);
  and (_20668_, _20667_, _01320_);
  and (_20669_, _20668_, _20666_);
  or (_20670_, _20669_, _20587_);
  and (_42924_, _20670_, _42355_);
  not (_20671_, \oc8051_golden_model_1.DPL [1]);
  nor (_20672_, _07950_, _20671_);
  nor (_20673_, _11252_, _11595_);
  or (_20674_, _20673_, _20672_);
  or (_20675_, _20674_, _07231_);
  or (_20676_, _09339_, _11595_);
  or (_20677_, _07950_, \oc8051_golden_model_1.DPL [1]);
  and (_20679_, _20677_, _09486_);
  and (_20680_, _20679_, _20676_);
  and (_20681_, _14520_, _07950_);
  not (_20682_, _20681_);
  and (_20683_, _20682_, _20677_);
  or (_20684_, _20683_, _06286_);
  and (_20685_, _07950_, \oc8051_golden_model_1.ACC [1]);
  or (_20686_, _20685_, _20672_);
  and (_20687_, _20686_, _07143_);
  nor (_20688_, _07143_, _20671_);
  or (_20691_, _20688_, _06285_);
  or (_20692_, _20691_, _20687_);
  and (_20693_, _20692_, _07169_);
  and (_20694_, _20693_, _20684_);
  and (_20695_, _07950_, _09422_);
  or (_20696_, _20695_, _20672_);
  and (_20697_, _20696_, _06354_);
  or (_20698_, _20697_, _06345_);
  or (_20699_, _20698_, _20694_);
  or (_20700_, _20686_, _06346_);
  and (_20702_, _20700_, _11536_);
  and (_20703_, _20702_, _20699_);
  nor (_20704_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_20705_, _20704_, _11540_);
  and (_20706_, _20705_, _11535_);
  or (_20707_, _20706_, _20703_);
  and (_20708_, _20707_, _06396_);
  nor (_20709_, _07031_, _06396_);
  or (_20710_, _20709_, _06259_);
  or (_20711_, _20710_, _20708_);
  or (_20712_, _20696_, _06260_);
  and (_20713_, _20712_, _06258_);
  and (_20714_, _20713_, _20711_);
  or (_20715_, _20714_, _20680_);
  and (_20716_, _20715_, _06251_);
  or (_20717_, _14607_, _11595_);
  and (_20718_, _20677_, _05972_);
  and (_20719_, _20718_, _20717_);
  or (_20720_, _20719_, _20716_);
  and (_20721_, _20720_, _06399_);
  or (_20723_, _14505_, _11595_);
  and (_20724_, _20723_, _06398_);
  nand (_20725_, _07950_, _07031_);
  and (_20726_, _20725_, _06215_);
  or (_20727_, _20726_, _20724_);
  and (_20728_, _20727_, _20677_);
  or (_20729_, _20728_, _06524_);
  or (_20730_, _20729_, _20721_);
  nand (_20731_, _11251_, _07950_);
  and (_20732_, _20731_, _20674_);
  or (_20735_, _20732_, _09030_);
  and (_20736_, _20735_, _07219_);
  and (_20737_, _20736_, _20730_);
  or (_20738_, _14503_, _11595_);
  and (_20739_, _20677_, _06426_);
  and (_20740_, _20739_, _20738_);
  or (_20741_, _20740_, _06532_);
  or (_20742_, _20741_, _20737_);
  nor (_20743_, _20672_, _07217_);
  nand (_20744_, _20743_, _20731_);
  and (_20745_, _20744_, _07229_);
  and (_20746_, _20745_, _20742_);
  or (_20747_, _20725_, _08325_);
  and (_20748_, _20677_, _06437_);
  and (_20749_, _20748_, _20747_);
  or (_20750_, _20749_, _06535_);
  or (_20751_, _20750_, _20746_);
  and (_20752_, _20751_, _20675_);
  or (_20753_, _20752_, _06559_);
  or (_20754_, _20683_, _07240_);
  and (_20756_, _20754_, _06570_);
  and (_20757_, _20756_, _20753_);
  or (_20758_, _20681_, _20672_);
  and (_20759_, _20758_, _06566_);
  or (_20760_, _20759_, _01324_);
  or (_20761_, _20760_, _20757_);
  or (_20762_, _01320_, \oc8051_golden_model_1.DPL [1]);
  and (_20763_, _20762_, _42355_);
  and (_42925_, _20763_, _20761_);
  not (_20764_, \oc8051_golden_model_1.DPL [2]);
  nor (_20767_, _01320_, _20764_);
  nor (_20768_, _07950_, _20764_);
  and (_20769_, _07950_, _08662_);
  or (_20770_, _20769_, _20768_);
  or (_20771_, _20770_, _06260_);
  and (_20772_, _14703_, _07950_);
  or (_20773_, _20772_, _20768_);
  or (_20774_, _20773_, _06286_);
  and (_20775_, _07950_, \oc8051_golden_model_1.ACC [2]);
  or (_20776_, _20775_, _20768_);
  and (_20778_, _20776_, _07143_);
  nor (_20779_, _07143_, _20764_);
  or (_20780_, _20779_, _06285_);
  or (_20781_, _20780_, _20778_);
  and (_20782_, _20781_, _07169_);
  and (_20783_, _20782_, _20774_);
  and (_20784_, _20770_, _06354_);
  or (_20785_, _20784_, _06345_);
  or (_20786_, _20785_, _20783_);
  or (_20787_, _20776_, _06346_);
  and (_20789_, _20787_, _11536_);
  and (_20790_, _20789_, _20786_);
  nor (_20791_, _11540_, \oc8051_golden_model_1.DPL [2]);
  nor (_20792_, _20791_, _11541_);
  and (_20793_, _20792_, _11535_);
  or (_20794_, _20793_, _20790_);
  and (_20795_, _20794_, _06396_);
  nor (_20796_, _06689_, _06396_);
  or (_20797_, _20796_, _06259_);
  or (_20798_, _20797_, _20795_);
  and (_20800_, _20798_, _20771_);
  or (_20801_, _20800_, _09486_);
  and (_20802_, _09293_, _07950_);
  or (_20803_, _20768_, _06258_);
  or (_20804_, _20803_, _20802_);
  and (_20805_, _20804_, _06251_);
  and (_20806_, _20805_, _20801_);
  and (_20807_, _14804_, _07950_);
  or (_20808_, _20807_, _20768_);
  and (_20809_, _20808_, _05972_);
  or (_20810_, _20809_, _20806_);
  or (_20811_, _20810_, _10080_);
  and (_20812_, _14697_, _07950_);
  or (_20813_, _20768_, _09025_);
  or (_20814_, _20813_, _20812_);
  and (_20815_, _07950_, _08980_);
  or (_20816_, _20815_, _20768_);
  or (_20817_, _20816_, _06216_);
  and (_20818_, _20817_, _09030_);
  and (_20819_, _20818_, _20814_);
  and (_20822_, _20819_, _20811_);
  and (_20823_, _11250_, _07950_);
  or (_20824_, _20823_, _20768_);
  and (_20825_, _20824_, _06524_);
  or (_20826_, _20825_, _20822_);
  and (_20827_, _20826_, _07219_);
  or (_20828_, _20768_, _08424_);
  and (_20829_, _20816_, _06426_);
  and (_20830_, _20829_, _20828_);
  or (_20831_, _20830_, _20827_);
  and (_20833_, _20831_, _07217_);
  and (_20834_, _20776_, _06532_);
  and (_20835_, _20834_, _20828_);
  or (_20836_, _20835_, _06437_);
  or (_20837_, _20836_, _20833_);
  and (_20838_, _14694_, _07950_);
  or (_20839_, _20768_, _07229_);
  or (_20840_, _20839_, _20838_);
  and (_20841_, _20840_, _07231_);
  and (_20842_, _20841_, _20837_);
  nor (_20844_, _11249_, _11595_);
  or (_20845_, _20844_, _20768_);
  and (_20846_, _20845_, _06535_);
  or (_20847_, _20846_, _20842_);
  and (_20848_, _20847_, _07240_);
  and (_20849_, _20773_, _06559_);
  or (_20850_, _20849_, _06566_);
  or (_20851_, _20850_, _20848_);
  and (_20852_, _14873_, _07950_);
  or (_20853_, _20768_, _06570_);
  or (_20855_, _20853_, _20852_);
  and (_20856_, _20855_, _01320_);
  and (_20857_, _20856_, _20851_);
  or (_20858_, _20857_, _20767_);
  and (_42926_, _20858_, _42355_);
  and (_20859_, _11595_, \oc8051_golden_model_1.DPL [3]);
  and (_20860_, _14900_, _07950_);
  or (_20861_, _20860_, _20859_);
  or (_20862_, _20861_, _06286_);
  and (_20863_, _07950_, \oc8051_golden_model_1.ACC [3]);
  or (_20865_, _20863_, _20859_);
  and (_20866_, _20865_, _07143_);
  and (_20867_, _07144_, \oc8051_golden_model_1.DPL [3]);
  or (_20868_, _20867_, _06285_);
  or (_20869_, _20868_, _20866_);
  and (_20870_, _20869_, _07169_);
  and (_20871_, _20870_, _20862_);
  and (_20872_, _07950_, _09421_);
  or (_20873_, _20872_, _20859_);
  and (_20874_, _20873_, _06354_);
  or (_20876_, _20874_, _06345_);
  or (_20877_, _20876_, _20871_);
  or (_20878_, _20865_, _06346_);
  and (_20879_, _20878_, _11536_);
  and (_20880_, _20879_, _20877_);
  nor (_20881_, _11541_, \oc8051_golden_model_1.DPL [3]);
  nor (_20882_, _20881_, _11542_);
  and (_20883_, _20882_, _11535_);
  or (_20884_, _20883_, _20880_);
  and (_20885_, _20884_, _06396_);
  nor (_20887_, _06517_, _06396_);
  or (_20888_, _20887_, _06259_);
  or (_20889_, _20888_, _20885_);
  or (_20890_, _20873_, _06260_);
  and (_20891_, _20890_, _20889_);
  or (_20892_, _20891_, _09486_);
  and (_20893_, _09247_, _07950_);
  or (_20894_, _20859_, _06258_);
  or (_20895_, _20894_, _20893_);
  and (_20896_, _20895_, _06251_);
  and (_20898_, _20896_, _20892_);
  and (_20899_, _14998_, _07950_);
  or (_20900_, _20899_, _20859_);
  and (_20901_, _20900_, _05972_);
  or (_20902_, _20901_, _10080_);
  or (_20903_, _20902_, _20898_);
  and (_20904_, _14893_, _07950_);
  or (_20905_, _20859_, _09025_);
  or (_20906_, _20905_, _20904_);
  and (_20907_, _07950_, _08809_);
  or (_20909_, _20907_, _20859_);
  or (_20910_, _20909_, _06216_);
  and (_20911_, _20910_, _09030_);
  and (_20912_, _20911_, _20906_);
  and (_20913_, _20912_, _20903_);
  and (_20914_, _12529_, _07950_);
  or (_20915_, _20914_, _20859_);
  and (_20916_, _20915_, _06524_);
  or (_20917_, _20916_, _20913_);
  and (_20918_, _20917_, _07219_);
  or (_20920_, _20859_, _08280_);
  and (_20921_, _20909_, _06426_);
  and (_20922_, _20921_, _20920_);
  or (_20923_, _20922_, _20918_);
  and (_20924_, _20923_, _07217_);
  and (_20925_, _20865_, _06532_);
  and (_20926_, _20925_, _20920_);
  or (_20927_, _20926_, _06437_);
  or (_20928_, _20927_, _20924_);
  and (_20929_, _14890_, _07950_);
  or (_20931_, _20859_, _07229_);
  or (_20932_, _20931_, _20929_);
  and (_20933_, _20932_, _07231_);
  and (_20934_, _20933_, _20928_);
  nor (_20935_, _11247_, _11595_);
  or (_20936_, _20935_, _20859_);
  and (_20937_, _20936_, _06535_);
  or (_20938_, _20937_, _06559_);
  or (_20939_, _20938_, _20934_);
  or (_20940_, _20861_, _07240_);
  and (_20941_, _20940_, _06570_);
  and (_20942_, _20941_, _20939_);
  and (_20943_, _15068_, _07950_);
  or (_20944_, _20943_, _20859_);
  and (_20945_, _20944_, _06566_);
  or (_20946_, _20945_, _01324_);
  or (_20947_, _20946_, _20942_);
  or (_20948_, _01320_, \oc8051_golden_model_1.DPL [3]);
  and (_20949_, _20948_, _42355_);
  and (_42927_, _20949_, _20947_);
  and (_20952_, _11595_, \oc8051_golden_model_1.DPL [4]);
  and (_20953_, _09420_, _07950_);
  or (_20954_, _20953_, _20952_);
  or (_20955_, _20954_, _06260_);
  and (_20956_, _15133_, _07950_);
  or (_20957_, _20956_, _20952_);
  or (_20958_, _20957_, _06286_);
  and (_20959_, _07950_, \oc8051_golden_model_1.ACC [4]);
  or (_20960_, _20959_, _20952_);
  and (_20961_, _20960_, _07143_);
  and (_20963_, _07144_, \oc8051_golden_model_1.DPL [4]);
  or (_20964_, _20963_, _06285_);
  or (_20965_, _20964_, _20961_);
  and (_20966_, _20965_, _07169_);
  and (_20967_, _20966_, _20958_);
  and (_20968_, _20954_, _06354_);
  or (_20969_, _20968_, _06345_);
  or (_20970_, _20969_, _20967_);
  or (_20971_, _20960_, _06346_);
  and (_20972_, _20971_, _11536_);
  and (_20974_, _20972_, _20970_);
  nor (_20975_, _11542_, \oc8051_golden_model_1.DPL [4]);
  nor (_20976_, _20975_, _11543_);
  and (_20977_, _20976_, _11535_);
  or (_20978_, _20977_, _20974_);
  and (_20979_, _20978_, _06396_);
  nor (_20980_, _08879_, _06396_);
  or (_20981_, _20980_, _06259_);
  or (_20982_, _20981_, _20979_);
  and (_20983_, _20982_, _20955_);
  or (_20985_, _20983_, _09486_);
  and (_20986_, _09437_, _07950_);
  or (_20987_, _20952_, _06258_);
  or (_20988_, _20987_, _20986_);
  and (_20989_, _20988_, _06251_);
  and (_20990_, _20989_, _20985_);
  and (_20991_, _15226_, _07950_);
  or (_20992_, _20991_, _20952_);
  and (_20993_, _20992_, _05972_);
  or (_20994_, _20993_, _20990_);
  or (_20996_, _20994_, _10080_);
  and (_20997_, _15114_, _07950_);
  or (_20998_, _20952_, _09025_);
  or (_20999_, _20998_, _20997_);
  and (_21000_, _08919_, _07950_);
  or (_21001_, _21000_, _20952_);
  or (_21002_, _21001_, _06216_);
  and (_21003_, _21002_, _09030_);
  and (_21004_, _21003_, _20999_);
  and (_21005_, _21004_, _20996_);
  and (_21007_, _11245_, _07950_);
  or (_21008_, _21007_, _20952_);
  and (_21009_, _21008_, _06524_);
  or (_21010_, _21009_, _21005_);
  and (_21011_, _21010_, _07219_);
  or (_21012_, _20952_, _08528_);
  and (_21013_, _21001_, _06426_);
  and (_21014_, _21013_, _21012_);
  or (_21015_, _21014_, _21011_);
  and (_21016_, _21015_, _07217_);
  and (_21018_, _20960_, _06532_);
  and (_21019_, _21018_, _21012_);
  or (_21020_, _21019_, _06437_);
  or (_21021_, _21020_, _21016_);
  and (_21022_, _15111_, _07950_);
  or (_21023_, _20952_, _07229_);
  or (_21024_, _21023_, _21022_);
  and (_21025_, _21024_, _07231_);
  and (_21026_, _21025_, _21021_);
  nor (_21027_, _11244_, _11595_);
  or (_21029_, _21027_, _20952_);
  and (_21030_, _21029_, _06535_);
  or (_21031_, _21030_, _06559_);
  or (_21032_, _21031_, _21026_);
  or (_21033_, _20957_, _07240_);
  and (_21034_, _21033_, _06570_);
  and (_21035_, _21034_, _21032_);
  and (_21036_, _15296_, _07950_);
  or (_21037_, _21036_, _20952_);
  and (_21038_, _21037_, _06566_);
  or (_21040_, _21038_, _01324_);
  or (_21041_, _21040_, _21035_);
  or (_21042_, _01320_, \oc8051_golden_model_1.DPL [4]);
  and (_21043_, _21042_, _42355_);
  and (_42928_, _21043_, _21041_);
  and (_21044_, _11595_, \oc8051_golden_model_1.DPL [5]);
  and (_21045_, _09419_, _07950_);
  or (_21046_, _21045_, _21044_);
  or (_21047_, _21046_, _06260_);
  and (_21048_, _15330_, _07950_);
  or (_21050_, _21048_, _21044_);
  or (_21051_, _21050_, _06286_);
  and (_21052_, _07950_, \oc8051_golden_model_1.ACC [5]);
  or (_21053_, _21052_, _21044_);
  and (_21054_, _21053_, _07143_);
  and (_21055_, _07144_, \oc8051_golden_model_1.DPL [5]);
  or (_21056_, _21055_, _06285_);
  or (_21057_, _21056_, _21054_);
  and (_21058_, _21057_, _07169_);
  and (_21059_, _21058_, _21051_);
  and (_21061_, _21046_, _06354_);
  or (_21062_, _21061_, _06345_);
  or (_21063_, _21062_, _21059_);
  or (_21064_, _21053_, _06346_);
  and (_21065_, _21064_, _11536_);
  and (_21066_, _21065_, _21063_);
  nor (_21067_, _11543_, \oc8051_golden_model_1.DPL [5]);
  nor (_21068_, _21067_, _11544_);
  and (_21069_, _21068_, _11535_);
  or (_21070_, _21069_, _21066_);
  and (_21072_, _21070_, _06396_);
  and (_21073_, _08913_, _06395_);
  or (_21074_, _21073_, _06259_);
  or (_21075_, _21074_, _21072_);
  and (_21076_, _21075_, _21047_);
  or (_21077_, _21076_, _09486_);
  and (_21078_, _09436_, _07950_);
  or (_21079_, _21044_, _06258_);
  or (_21080_, _21079_, _21078_);
  and (_21081_, _21080_, _06251_);
  and (_21083_, _21081_, _21077_);
  and (_21084_, _15421_, _07950_);
  or (_21085_, _21084_, _21044_);
  and (_21086_, _21085_, _05972_);
  or (_21087_, _21086_, _21083_);
  or (_21088_, _21087_, _10080_);
  and (_21089_, _15313_, _07950_);
  or (_21090_, _21044_, _09025_);
  or (_21091_, _21090_, _21089_);
  and (_21092_, _08913_, _07950_);
  or (_21094_, _21092_, _21044_);
  or (_21095_, _21094_, _06216_);
  and (_21096_, _21095_, _09030_);
  and (_21097_, _21096_, _21091_);
  and (_21098_, _21097_, _21088_);
  and (_21099_, _12536_, _07950_);
  or (_21100_, _21099_, _21044_);
  and (_21101_, _21100_, _06524_);
  or (_21102_, _21101_, _21098_);
  and (_21103_, _21102_, _07219_);
  or (_21105_, _21044_, _08231_);
  and (_21106_, _21094_, _06426_);
  and (_21107_, _21106_, _21105_);
  or (_21108_, _21107_, _21103_);
  and (_21109_, _21108_, _07217_);
  and (_21110_, _21053_, _06532_);
  and (_21111_, _21110_, _21105_);
  or (_21112_, _21111_, _06437_);
  or (_21113_, _21112_, _21109_);
  and (_21114_, _15310_, _07950_);
  or (_21115_, _21044_, _07229_);
  or (_21116_, _21115_, _21114_);
  and (_21117_, _21116_, _07231_);
  and (_21118_, _21117_, _21113_);
  nor (_21119_, _11241_, _11595_);
  or (_21120_, _21119_, _21044_);
  and (_21121_, _21120_, _06535_);
  or (_21122_, _21121_, _06559_);
  or (_21123_, _21122_, _21118_);
  or (_21124_, _21050_, _07240_);
  and (_21127_, _21124_, _06570_);
  and (_21128_, _21127_, _21123_);
  and (_21129_, _15493_, _07950_);
  or (_21130_, _21129_, _21044_);
  and (_21131_, _21130_, _06566_);
  or (_21132_, _21131_, _01324_);
  or (_21133_, _21132_, _21128_);
  or (_21134_, _01320_, \oc8051_golden_model_1.DPL [5]);
  and (_21135_, _21134_, _42355_);
  and (_42929_, _21135_, _21133_);
  and (_21137_, _11595_, \oc8051_golden_model_1.DPL [6]);
  and (_21138_, _09418_, _07950_);
  or (_21139_, _21138_, _21137_);
  or (_21140_, _21139_, _06260_);
  and (_21141_, _15521_, _07950_);
  or (_21142_, _21141_, _21137_);
  or (_21143_, _21142_, _06286_);
  and (_21144_, _07950_, \oc8051_golden_model_1.ACC [6]);
  or (_21145_, _21144_, _21137_);
  and (_21146_, _21145_, _07143_);
  and (_21148_, _07144_, \oc8051_golden_model_1.DPL [6]);
  or (_21149_, _21148_, _06285_);
  or (_21150_, _21149_, _21146_);
  and (_21151_, _21150_, _07169_);
  and (_21152_, _21151_, _21143_);
  and (_21153_, _21139_, _06354_);
  or (_21154_, _21153_, _06345_);
  or (_21155_, _21154_, _21152_);
  or (_21156_, _21145_, _06346_);
  and (_21157_, _21156_, _11536_);
  and (_21159_, _21157_, _21155_);
  nor (_21160_, _11544_, \oc8051_golden_model_1.DPL [6]);
  nor (_21161_, _21160_, _11545_);
  and (_21162_, _21161_, _11535_);
  or (_21163_, _21162_, _21159_);
  and (_21164_, _21163_, _06396_);
  nor (_21165_, _08844_, _06396_);
  or (_21166_, _21165_, _06259_);
  or (_21167_, _21166_, _21164_);
  and (_21168_, _21167_, _21140_);
  or (_21170_, _21168_, _09486_);
  and (_21171_, _09435_, _07950_);
  or (_21172_, _21137_, _06258_);
  or (_21173_, _21172_, _21171_);
  and (_21174_, _21173_, _06251_);
  and (_21175_, _21174_, _21170_);
  and (_21176_, _15623_, _07950_);
  or (_21177_, _21176_, _21137_);
  and (_21178_, _21177_, _05972_);
  or (_21179_, _21178_, _21175_);
  or (_21181_, _21179_, _10080_);
  and (_21182_, _15517_, _07950_);
  or (_21183_, _21137_, _09025_);
  or (_21184_, _21183_, _21182_);
  and (_21185_, _08845_, _07950_);
  or (_21186_, _21185_, _21137_);
  or (_21187_, _21186_, _06216_);
  and (_21188_, _21187_, _09030_);
  and (_21189_, _21188_, _21184_);
  and (_21190_, _21189_, _21181_);
  and (_21192_, _11239_, _07950_);
  or (_21193_, _21192_, _21137_);
  and (_21194_, _21193_, _06524_);
  or (_21195_, _21194_, _21190_);
  and (_21196_, _21195_, _07219_);
  or (_21197_, _21137_, _08128_);
  and (_21198_, _21186_, _06426_);
  and (_21199_, _21198_, _21197_);
  or (_21200_, _21199_, _21196_);
  and (_21201_, _21200_, _07217_);
  and (_21203_, _21145_, _06532_);
  and (_21204_, _21203_, _21197_);
  or (_21205_, _21204_, _06437_);
  or (_21206_, _21205_, _21201_);
  and (_21207_, _15514_, _07950_);
  or (_21208_, _21137_, _07229_);
  or (_21209_, _21208_, _21207_);
  and (_21210_, _21209_, _07231_);
  and (_21211_, _21210_, _21206_);
  nor (_21212_, _11238_, _11595_);
  or (_21214_, _21212_, _21137_);
  and (_21215_, _21214_, _06535_);
  or (_21216_, _21215_, _06559_);
  or (_21217_, _21216_, _21211_);
  or (_21218_, _21142_, _07240_);
  and (_21219_, _21218_, _06570_);
  and (_21220_, _21219_, _21217_);
  and (_21221_, _15695_, _07950_);
  or (_21222_, _21221_, _21137_);
  and (_21223_, _21222_, _06566_);
  or (_21225_, _21223_, _01324_);
  or (_21226_, _21225_, _21220_);
  or (_21227_, _01320_, \oc8051_golden_model_1.DPL [6]);
  and (_21228_, _21227_, _42355_);
  and (_42930_, _21228_, _21226_);
  and (_21229_, _01324_, \oc8051_golden_model_1.DPH [0]);
  not (_21230_, _07953_);
  and (_21231_, _21230_, \oc8051_golden_model_1.DPH [0]);
  and (_21232_, _07953_, \oc8051_golden_model_1.ACC [0]);
  and (_21233_, _21232_, _08374_);
  or (_21235_, _21233_, _21231_);
  or (_21236_, _21235_, _07217_);
  nor (_21237_, _11547_, \oc8051_golden_model_1.DPH [0]);
  nor (_21238_, _21237_, _11633_);
  and (_21239_, _21238_, _11535_);
  nor (_21240_, _08374_, _11689_);
  or (_21241_, _21240_, _21231_);
  or (_21242_, _21241_, _06286_);
  or (_21243_, _21232_, _21231_);
  and (_21244_, _21243_, _07143_);
  and (_21246_, _07144_, \oc8051_golden_model_1.DPH [0]);
  or (_21247_, _21246_, _06285_);
  or (_21248_, _21247_, _21244_);
  and (_21249_, _21248_, _07169_);
  and (_21250_, _21249_, _21242_);
  and (_21251_, _08261_, _07135_);
  or (_21252_, _21251_, _21231_);
  and (_21253_, _21252_, _06354_);
  or (_21254_, _21253_, _06345_);
  or (_21255_, _21254_, _21250_);
  or (_21257_, _21243_, _06346_);
  and (_21258_, _21257_, _11536_);
  and (_21259_, _21258_, _21255_);
  or (_21260_, _21259_, _21239_);
  and (_21261_, _21260_, _06396_);
  and (_21262_, _06395_, _06248_);
  or (_21263_, _21262_, _06259_);
  or (_21264_, _21263_, _21261_);
  or (_21265_, _21252_, _06260_);
  and (_21266_, _21265_, _21264_);
  or (_21268_, _21266_, _09486_);
  and (_21269_, _09384_, _07953_);
  or (_21270_, _21231_, _06258_);
  or (_21271_, _21270_, _21269_);
  and (_21272_, _21271_, _21268_);
  or (_21273_, _21272_, _05972_);
  and (_21274_, _14413_, _08261_);
  or (_21275_, _21231_, _06251_);
  or (_21276_, _21275_, _21274_);
  and (_21277_, _21276_, _06216_);
  and (_21279_, _21277_, _21273_);
  and (_21280_, _07953_, _08929_);
  or (_21281_, _21280_, _21231_);
  and (_21282_, _21281_, _06215_);
  or (_21283_, _21282_, _06398_);
  or (_21284_, _21283_, _21279_);
  and (_21285_, _14311_, _07953_);
  or (_21286_, _21285_, _21231_);
  or (_21287_, _21286_, _09025_);
  and (_21288_, _21287_, _09030_);
  and (_21290_, _21288_, _21284_);
  nor (_21291_, _12532_, _11689_);
  or (_21292_, _21291_, _21231_);
  nor (_21293_, _21233_, _09030_);
  and (_21294_, _21293_, _21292_);
  or (_21295_, _21294_, _21290_);
  and (_21296_, _21295_, _07219_);
  nand (_21297_, _21281_, _06426_);
  nor (_21298_, _21297_, _21240_);
  or (_21299_, _21298_, _06532_);
  or (_21301_, _21299_, _21296_);
  and (_21302_, _21301_, _21236_);
  or (_21303_, _21302_, _06437_);
  and (_21304_, _14307_, _07953_);
  or (_21305_, _21304_, _21231_);
  or (_21306_, _21305_, _07229_);
  and (_21307_, _21306_, _07231_);
  and (_21308_, _21307_, _21303_);
  and (_21309_, _21292_, _06535_);
  or (_21310_, _21309_, _19480_);
  or (_21311_, _21310_, _21308_);
  or (_21312_, _21241_, _06651_);
  and (_21313_, _21312_, _01320_);
  and (_21314_, _21313_, _21311_);
  or (_21315_, _21314_, _21229_);
  and (_42932_, _21315_, _42355_);
  and (_21316_, _21230_, \oc8051_golden_model_1.DPH [1]);
  nor (_21317_, _11252_, _11689_);
  or (_21318_, _21317_, _21316_);
  or (_21319_, _21318_, _07231_);
  or (_21322_, _09339_, _11689_);
  or (_21323_, _07953_, \oc8051_golden_model_1.DPH [1]);
  and (_21324_, _21323_, _09486_);
  and (_21325_, _21324_, _21322_);
  nor (_21326_, _11633_, \oc8051_golden_model_1.DPH [1]);
  nor (_21327_, _21326_, _11634_);
  and (_21328_, _21327_, _11535_);
  and (_21329_, _14520_, _08261_);
  not (_21330_, _21329_);
  and (_21331_, _21330_, _21323_);
  or (_21333_, _21331_, _06286_);
  and (_21334_, _07953_, \oc8051_golden_model_1.ACC [1]);
  or (_21335_, _21334_, _21316_);
  and (_21336_, _21335_, _07143_);
  and (_21337_, _07144_, \oc8051_golden_model_1.DPH [1]);
  or (_21338_, _21337_, _06285_);
  or (_21339_, _21338_, _21336_);
  and (_21340_, _21339_, _07169_);
  and (_21341_, _21340_, _21333_);
  and (_21342_, _08261_, _09422_);
  or (_21344_, _21342_, _21316_);
  and (_21345_, _21344_, _06354_);
  or (_21346_, _21345_, _06345_);
  or (_21347_, _21346_, _21341_);
  or (_21348_, _21335_, _06346_);
  and (_21349_, _21348_, _11536_);
  and (_21350_, _21349_, _21347_);
  or (_21351_, _21350_, _21328_);
  and (_21352_, _21351_, _06396_);
  nor (_21353_, _06995_, _06396_);
  or (_21355_, _21353_, _06259_);
  or (_21356_, _21355_, _21352_);
  or (_21357_, _21344_, _06260_);
  and (_21358_, _21357_, _06258_);
  and (_21359_, _21358_, _21356_);
  or (_21360_, _21359_, _21325_);
  and (_21361_, _21360_, _06251_);
  and (_21362_, _14607_, _07953_);
  or (_21363_, _21362_, _21316_);
  and (_21364_, _21363_, _05972_);
  or (_21366_, _21364_, _21361_);
  and (_21367_, _21366_, _06399_);
  or (_21368_, _14505_, _11689_);
  and (_21369_, _21368_, _06398_);
  nand (_21370_, _08261_, _07031_);
  and (_21371_, _21370_, _06215_);
  or (_21372_, _21371_, _21369_);
  and (_21373_, _21372_, _21323_);
  or (_21374_, _21373_, _06524_);
  or (_21375_, _21374_, _21367_);
  nand (_21377_, _11251_, _08261_);
  and (_21378_, _21377_, _21318_);
  or (_21379_, _21378_, _09030_);
  and (_21380_, _21379_, _07219_);
  and (_21381_, _21380_, _21375_);
  or (_21382_, _14503_, _11689_);
  and (_21383_, _21323_, _06426_);
  and (_21384_, _21383_, _21382_);
  or (_21385_, _21384_, _06532_);
  or (_21386_, _21385_, _21381_);
  nor (_21388_, _21316_, _07217_);
  nand (_21389_, _21388_, _21377_);
  and (_21390_, _21389_, _07229_);
  and (_21391_, _21390_, _21386_);
  or (_21392_, _21370_, _08325_);
  and (_21393_, _21323_, _06437_);
  and (_21394_, _21393_, _21392_);
  or (_21395_, _21394_, _06535_);
  or (_21396_, _21395_, _21391_);
  and (_21397_, _21396_, _21319_);
  or (_21399_, _21397_, _06559_);
  or (_21400_, _21331_, _07240_);
  and (_21401_, _21400_, _06570_);
  and (_21402_, _21401_, _21399_);
  or (_21403_, _21329_, _21316_);
  and (_21404_, _21403_, _06566_);
  or (_21405_, _21404_, _01324_);
  or (_21406_, _21405_, _21402_);
  or (_21407_, _01320_, \oc8051_golden_model_1.DPH [1]);
  and (_21408_, _21407_, _42355_);
  and (_42933_, _21408_, _21406_);
  and (_21410_, _01324_, \oc8051_golden_model_1.DPH [2]);
  or (_21411_, _11634_, \oc8051_golden_model_1.DPH [2]);
  nor (_21412_, _11635_, _11536_);
  and (_21413_, _21412_, _21411_);
  and (_21414_, _21230_, \oc8051_golden_model_1.DPH [2]);
  and (_21415_, _08261_, _08662_);
  or (_21416_, _21415_, _21414_);
  or (_21417_, _21416_, _07169_);
  and (_21418_, _14703_, _08261_);
  or (_21420_, _21418_, _21414_);
  and (_21421_, _21420_, _06285_);
  and (_21422_, _07144_, \oc8051_golden_model_1.DPH [2]);
  and (_21423_, _07953_, \oc8051_golden_model_1.ACC [2]);
  or (_21424_, _21423_, _21414_);
  and (_21425_, _21424_, _07143_);
  or (_21426_, _21425_, _21422_);
  and (_21427_, _21426_, _06286_);
  or (_21428_, _21427_, _06354_);
  or (_21429_, _21428_, _21421_);
  and (_21431_, _21429_, _21417_);
  or (_21432_, _21431_, _06345_);
  or (_21433_, _21424_, _06346_);
  and (_21434_, _21433_, _11536_);
  and (_21435_, _21434_, _21432_);
  or (_21436_, _21435_, _21413_);
  and (_21437_, _21436_, _06396_);
  nor (_21438_, _06646_, _06396_);
  or (_21439_, _21438_, _06259_);
  or (_21440_, _21439_, _21437_);
  or (_21442_, _21416_, _06260_);
  and (_21443_, _21442_, _21440_);
  or (_21444_, _21443_, _09486_);
  and (_21445_, _09293_, _07953_);
  or (_21446_, _21414_, _06258_);
  or (_21447_, _21446_, _21445_);
  and (_21448_, _21447_, _06251_);
  and (_21449_, _21448_, _21444_);
  and (_21450_, _14804_, _08261_);
  or (_21451_, _21450_, _21414_);
  and (_21453_, _21451_, _05972_);
  or (_21454_, _21453_, _10080_);
  or (_21455_, _21454_, _21449_);
  and (_21456_, _14697_, _08261_);
  or (_21457_, _21414_, _09025_);
  or (_21458_, _21457_, _21456_);
  and (_21459_, _07953_, _08980_);
  or (_21460_, _21459_, _21414_);
  or (_21461_, _21460_, _06216_);
  and (_21462_, _21461_, _09030_);
  and (_21464_, _21462_, _21458_);
  and (_21465_, _21464_, _21455_);
  and (_21466_, _11250_, _07953_);
  or (_21467_, _21466_, _21414_);
  and (_21468_, _21467_, _06524_);
  or (_21469_, _21468_, _21465_);
  and (_21470_, _21469_, _07219_);
  or (_21471_, _21414_, _08424_);
  and (_21472_, _21460_, _06426_);
  and (_21473_, _21472_, _21471_);
  or (_21475_, _21473_, _21470_);
  and (_21476_, _21475_, _07217_);
  and (_21477_, _21424_, _06532_);
  and (_21478_, _21477_, _21471_);
  or (_21479_, _21478_, _06437_);
  or (_21480_, _21479_, _21476_);
  and (_21481_, _14694_, _08261_);
  or (_21482_, _21414_, _07229_);
  or (_21483_, _21482_, _21481_);
  and (_21484_, _21483_, _07231_);
  and (_21486_, _21484_, _21480_);
  nor (_21487_, _11249_, _11689_);
  or (_21488_, _21487_, _21414_);
  and (_21489_, _21488_, _06535_);
  or (_21490_, _21489_, _21486_);
  and (_21491_, _21490_, _07240_);
  and (_21492_, _21420_, _06559_);
  or (_21493_, _21492_, _06566_);
  or (_21494_, _21493_, _21491_);
  and (_21495_, _14873_, _08261_);
  or (_21497_, _21414_, _06570_);
  or (_21498_, _21497_, _21495_);
  and (_21499_, _21498_, _01320_);
  and (_21500_, _21499_, _21494_);
  or (_21501_, _21500_, _21410_);
  and (_42934_, _21501_, _42355_);
  or (_21502_, _11635_, \oc8051_golden_model_1.DPH [3]);
  nor (_21503_, _11636_, _11536_);
  and (_21504_, _21503_, _21502_);
  and (_21505_, _21230_, \oc8051_golden_model_1.DPH [3]);
  and (_21507_, _14900_, _08261_);
  or (_21508_, _21507_, _21505_);
  or (_21509_, _21508_, _06286_);
  and (_21510_, _07953_, \oc8051_golden_model_1.ACC [3]);
  or (_21511_, _21510_, _21505_);
  and (_21512_, _21511_, _07143_);
  and (_21513_, _07144_, \oc8051_golden_model_1.DPH [3]);
  or (_21514_, _21513_, _06285_);
  or (_21515_, _21514_, _21512_);
  and (_21516_, _21515_, _07169_);
  and (_21518_, _21516_, _21509_);
  and (_21519_, _08261_, _09421_);
  or (_21520_, _21519_, _21505_);
  and (_21521_, _21520_, _06354_);
  or (_21522_, _21521_, _06345_);
  or (_21523_, _21522_, _21518_);
  or (_21524_, _21511_, _06346_);
  and (_21525_, _21524_, _11536_);
  and (_21526_, _21525_, _21523_);
  or (_21527_, _21526_, _21504_);
  and (_21529_, _21527_, _06396_);
  nor (_21530_, _06396_, _06212_);
  or (_21531_, _21530_, _06259_);
  or (_21532_, _21531_, _21529_);
  or (_21533_, _21520_, _06260_);
  and (_21534_, _21533_, _21532_);
  or (_21535_, _21534_, _09486_);
  and (_21536_, _09247_, _07953_);
  or (_21537_, _21505_, _06258_);
  or (_21538_, _21537_, _21536_);
  and (_21540_, _21538_, _06251_);
  and (_21541_, _21540_, _21535_);
  and (_21542_, _14998_, _08261_);
  or (_21543_, _21542_, _21505_);
  and (_21544_, _21543_, _05972_);
  or (_21545_, _21544_, _10080_);
  or (_21546_, _21545_, _21541_);
  and (_21547_, _14893_, _08261_);
  or (_21548_, _21505_, _09025_);
  or (_21549_, _21548_, _21547_);
  and (_21551_, _07953_, _08809_);
  or (_21552_, _21551_, _21505_);
  or (_21553_, _21552_, _06216_);
  and (_21554_, _21553_, _09030_);
  and (_21555_, _21554_, _21549_);
  and (_21556_, _21555_, _21546_);
  and (_21557_, _12529_, _07953_);
  or (_21558_, _21557_, _21505_);
  and (_21559_, _21558_, _06524_);
  or (_21560_, _21559_, _21556_);
  and (_21562_, _21560_, _07219_);
  or (_21563_, _21505_, _08280_);
  and (_21564_, _21552_, _06426_);
  and (_21565_, _21564_, _21563_);
  or (_21566_, _21565_, _21562_);
  and (_21567_, _21566_, _07217_);
  and (_21568_, _21511_, _06532_);
  and (_21569_, _21568_, _21563_);
  or (_21570_, _21569_, _06437_);
  or (_21571_, _21570_, _21567_);
  and (_21573_, _14890_, _08261_);
  or (_21574_, _21505_, _07229_);
  or (_21575_, _21574_, _21573_);
  and (_21576_, _21575_, _07231_);
  and (_21577_, _21576_, _21571_);
  nor (_21578_, _11247_, _11689_);
  or (_21579_, _21578_, _21505_);
  and (_21580_, _21579_, _06535_);
  or (_21581_, _21580_, _06559_);
  or (_21582_, _21581_, _21577_);
  or (_21584_, _21508_, _07240_);
  and (_21585_, _21584_, _06570_);
  and (_21586_, _21585_, _21582_);
  and (_21587_, _15068_, _08261_);
  or (_21588_, _21587_, _21505_);
  and (_21589_, _21588_, _06566_);
  or (_21590_, _21589_, _01324_);
  or (_21591_, _21590_, _21586_);
  or (_21592_, _01320_, \oc8051_golden_model_1.DPH [3]);
  and (_21593_, _21592_, _42355_);
  and (_42935_, _21593_, _21591_);
  and (_21595_, _21230_, \oc8051_golden_model_1.DPH [4]);
  and (_21596_, _09420_, _08261_);
  or (_21597_, _21596_, _21595_);
  or (_21598_, _21597_, _06260_);
  and (_21599_, _15133_, _08261_);
  or (_21600_, _21599_, _21595_);
  or (_21601_, _21600_, _06286_);
  and (_21602_, _07953_, \oc8051_golden_model_1.ACC [4]);
  or (_21603_, _21602_, _21595_);
  and (_21605_, _21603_, _07143_);
  and (_21606_, _07144_, \oc8051_golden_model_1.DPH [4]);
  or (_21607_, _21606_, _06285_);
  or (_21608_, _21607_, _21605_);
  and (_21609_, _21608_, _07169_);
  and (_21610_, _21609_, _21601_);
  and (_21611_, _21597_, _06354_);
  or (_21612_, _21611_, _06345_);
  or (_21613_, _21612_, _21610_);
  or (_21614_, _21603_, _06346_);
  and (_21616_, _21614_, _11536_);
  and (_21617_, _21616_, _21613_);
  or (_21618_, _11636_, \oc8051_golden_model_1.DPH [4]);
  nor (_21619_, _11637_, _11536_);
  and (_21620_, _21619_, _21618_);
  or (_21621_, _21620_, _21617_);
  and (_21622_, _21621_, _06396_);
  nor (_21623_, _06961_, _06396_);
  or (_21624_, _21623_, _06259_);
  or (_21625_, _21624_, _21622_);
  and (_21627_, _21625_, _21598_);
  or (_21628_, _21627_, _09486_);
  or (_21629_, _21595_, _06258_);
  and (_21630_, _09437_, _07953_);
  or (_21631_, _21630_, _21629_);
  and (_21632_, _21631_, _06251_);
  and (_21633_, _21632_, _21628_);
  and (_21634_, _15226_, _07953_);
  or (_21635_, _21634_, _21595_);
  and (_21636_, _21635_, _05972_);
  or (_21638_, _21636_, _21633_);
  or (_21639_, _21638_, _10080_);
  and (_21640_, _15114_, _08261_);
  or (_21641_, _21595_, _09025_);
  or (_21642_, _21641_, _21640_);
  and (_21643_, _08919_, _07953_);
  or (_21644_, _21643_, _21595_);
  or (_21645_, _21644_, _06216_);
  and (_21646_, _21645_, _09030_);
  and (_21647_, _21646_, _21642_);
  and (_21649_, _21647_, _21639_);
  and (_21650_, _11245_, _07953_);
  or (_21651_, _21650_, _21595_);
  and (_21652_, _21651_, _06524_);
  or (_21653_, _21652_, _21649_);
  and (_21654_, _21653_, _07219_);
  or (_21655_, _21595_, _08528_);
  and (_21656_, _21644_, _06426_);
  and (_21657_, _21656_, _21655_);
  or (_21658_, _21657_, _21654_);
  and (_21659_, _21658_, _07217_);
  and (_21660_, _21603_, _06532_);
  and (_21661_, _21660_, _21655_);
  or (_21662_, _21661_, _06437_);
  or (_21663_, _21662_, _21659_);
  and (_21664_, _15111_, _08261_);
  or (_21665_, _21595_, _07229_);
  or (_21666_, _21665_, _21664_);
  and (_21667_, _21666_, _07231_);
  and (_21668_, _21667_, _21663_);
  nor (_21671_, _11244_, _11689_);
  or (_21672_, _21671_, _21595_);
  and (_21673_, _21672_, _06535_);
  or (_21674_, _21673_, _06559_);
  or (_21675_, _21674_, _21668_);
  or (_21676_, _21600_, _07240_);
  and (_21677_, _21676_, _06570_);
  and (_21678_, _21677_, _21675_);
  and (_21679_, _15296_, _08261_);
  or (_21680_, _21679_, _21595_);
  and (_21682_, _21680_, _06566_);
  or (_21683_, _21682_, _01324_);
  or (_21684_, _21683_, _21678_);
  or (_21685_, _01320_, \oc8051_golden_model_1.DPH [4]);
  and (_21686_, _21685_, _42355_);
  and (_42936_, _21686_, _21684_);
  and (_21687_, _21230_, \oc8051_golden_model_1.DPH [5]);
  and (_21688_, _09419_, _08261_);
  or (_21689_, _21688_, _21687_);
  or (_21690_, _21689_, _06260_);
  and (_21692_, _15330_, _08261_);
  or (_21693_, _21692_, _21687_);
  or (_21694_, _21693_, _06286_);
  and (_21695_, _07953_, \oc8051_golden_model_1.ACC [5]);
  or (_21696_, _21695_, _21687_);
  and (_21697_, _21696_, _07143_);
  and (_21698_, _07144_, \oc8051_golden_model_1.DPH [5]);
  or (_21699_, _21698_, _06285_);
  or (_21700_, _21699_, _21697_);
  and (_21701_, _21700_, _07169_);
  and (_21703_, _21701_, _21694_);
  and (_21704_, _21689_, _06354_);
  or (_21705_, _21704_, _06345_);
  or (_21706_, _21705_, _21703_);
  or (_21707_, _21696_, _06346_);
  and (_21708_, _21707_, _11536_);
  and (_21709_, _21708_, _21706_);
  or (_21710_, _11637_, \oc8051_golden_model_1.DPH [5]);
  nor (_21711_, _11638_, _11536_);
  and (_21712_, _21711_, _21710_);
  or (_21714_, _21712_, _21709_);
  and (_21715_, _21714_, _06396_);
  nor (_21716_, _06604_, _06396_);
  or (_21717_, _21716_, _06259_);
  or (_21718_, _21717_, _21715_);
  and (_21719_, _21718_, _21690_);
  or (_21720_, _21719_, _09486_);
  or (_21721_, _21687_, _06258_);
  and (_21722_, _09436_, _07953_);
  or (_21723_, _21722_, _21721_);
  and (_21725_, _21723_, _06251_);
  and (_21726_, _21725_, _21720_);
  and (_21727_, _15421_, _07953_);
  or (_21728_, _21727_, _21687_);
  and (_21729_, _21728_, _05972_);
  or (_21730_, _21729_, _21726_);
  or (_21731_, _21730_, _10080_);
  and (_21732_, _15313_, _08261_);
  or (_21733_, _21687_, _09025_);
  or (_21734_, _21733_, _21732_);
  and (_21736_, _08913_, _07953_);
  or (_21737_, _21736_, _21687_);
  or (_21738_, _21737_, _06216_);
  and (_21739_, _21738_, _09030_);
  and (_21740_, _21739_, _21734_);
  and (_21741_, _21740_, _21731_);
  and (_21742_, _12536_, _07953_);
  or (_21743_, _21742_, _21687_);
  and (_21744_, _21743_, _06524_);
  or (_21745_, _21744_, _21741_);
  and (_21747_, _21745_, _07219_);
  or (_21748_, _21687_, _08231_);
  and (_21749_, _21737_, _06426_);
  and (_21750_, _21749_, _21748_);
  or (_21751_, _21750_, _21747_);
  and (_21752_, _21751_, _07217_);
  and (_21753_, _21696_, _06532_);
  and (_21754_, _21753_, _21748_);
  or (_21755_, _21754_, _06437_);
  or (_21756_, _21755_, _21752_);
  and (_21758_, _15310_, _08261_);
  or (_21759_, _21687_, _07229_);
  or (_21760_, _21759_, _21758_);
  and (_21761_, _21760_, _07231_);
  and (_21762_, _21761_, _21756_);
  nor (_21763_, _11241_, _11689_);
  or (_21764_, _21763_, _21687_);
  and (_21765_, _21764_, _06535_);
  or (_21766_, _21765_, _06559_);
  or (_21767_, _21766_, _21762_);
  or (_21768_, _21693_, _07240_);
  and (_21769_, _21768_, _06570_);
  and (_21770_, _21769_, _21767_);
  and (_21771_, _15493_, _08261_);
  or (_21772_, _21771_, _21687_);
  and (_21773_, _21772_, _06566_);
  or (_21774_, _21773_, _01324_);
  or (_21775_, _21774_, _21770_);
  or (_21776_, _01320_, \oc8051_golden_model_1.DPH [5]);
  and (_21777_, _21776_, _42355_);
  and (_42938_, _21777_, _21775_);
  and (_21780_, _21230_, \oc8051_golden_model_1.DPH [6]);
  and (_21781_, _09418_, _08261_);
  or (_21782_, _21781_, _21780_);
  or (_21783_, _21782_, _06260_);
  and (_21784_, _15521_, _08261_);
  or (_21785_, _21784_, _21780_);
  or (_21786_, _21785_, _06286_);
  and (_21787_, _07953_, \oc8051_golden_model_1.ACC [6]);
  or (_21788_, _21787_, _21780_);
  and (_21790_, _21788_, _07143_);
  and (_21791_, _07144_, \oc8051_golden_model_1.DPH [6]);
  or (_21792_, _21791_, _06285_);
  or (_21793_, _21792_, _21790_);
  and (_21794_, _21793_, _07169_);
  and (_21795_, _21794_, _21786_);
  and (_21796_, _21782_, _06354_);
  or (_21797_, _21796_, _06345_);
  or (_21798_, _21797_, _21795_);
  or (_21799_, _21788_, _06346_);
  and (_21801_, _21799_, _11536_);
  and (_21802_, _21801_, _21798_);
  or (_21803_, _11638_, \oc8051_golden_model_1.DPH [6]);
  nor (_21804_, _11639_, _11536_);
  and (_21805_, _21804_, _21803_);
  or (_21806_, _21805_, _21802_);
  and (_21807_, _21806_, _06396_);
  nor (_21808_, _06396_, _06325_);
  or (_21809_, _21808_, _06259_);
  or (_21810_, _21809_, _21807_);
  and (_21812_, _21810_, _21783_);
  or (_21813_, _21812_, _09486_);
  or (_21814_, _21780_, _06258_);
  and (_21815_, _09435_, _07953_);
  or (_21816_, _21815_, _21814_);
  and (_21817_, _21816_, _06251_);
  and (_21818_, _21817_, _21813_);
  and (_21819_, _15623_, _07953_);
  or (_21820_, _21819_, _21780_);
  and (_21821_, _21820_, _05972_);
  or (_21823_, _21821_, _21818_);
  or (_21824_, _21823_, _10080_);
  and (_21825_, _15517_, _08261_);
  or (_21826_, _21780_, _09025_);
  or (_21827_, _21826_, _21825_);
  and (_21828_, _08845_, _07953_);
  or (_21829_, _21828_, _21780_);
  or (_21830_, _21829_, _06216_);
  and (_21831_, _21830_, _09030_);
  and (_21832_, _21831_, _21827_);
  and (_21834_, _21832_, _21824_);
  and (_21835_, _11239_, _07953_);
  or (_21836_, _21835_, _21780_);
  and (_21837_, _21836_, _06524_);
  or (_21838_, _21837_, _21834_);
  and (_21839_, _21838_, _07219_);
  or (_21840_, _21780_, _08128_);
  and (_21841_, _21829_, _06426_);
  and (_21842_, _21841_, _21840_);
  or (_21843_, _21842_, _21839_);
  and (_21845_, _21843_, _07217_);
  and (_21846_, _21788_, _06532_);
  and (_21847_, _21846_, _21840_);
  or (_21848_, _21847_, _06437_);
  or (_21849_, _21848_, _21845_);
  and (_21850_, _15514_, _08261_);
  or (_21851_, _21780_, _07229_);
  or (_21852_, _21851_, _21850_);
  and (_21853_, _21852_, _07231_);
  and (_21854_, _21853_, _21849_);
  nor (_21856_, _11238_, _11689_);
  or (_21857_, _21856_, _21780_);
  and (_21858_, _21857_, _06535_);
  or (_21859_, _21858_, _06559_);
  or (_21860_, _21859_, _21854_);
  or (_21861_, _21785_, _07240_);
  and (_21862_, _21861_, _06570_);
  and (_21863_, _21862_, _21860_);
  and (_21864_, _15695_, _08261_);
  or (_21865_, _21864_, _21780_);
  and (_21867_, _21865_, _06566_);
  or (_21868_, _21867_, _01324_);
  or (_21869_, _21868_, _21863_);
  or (_21870_, _01320_, \oc8051_golden_model_1.DPH [6]);
  and (_21871_, _21870_, _42355_);
  and (_42939_, _21871_, _21869_);
  not (_21872_, \oc8051_golden_model_1.TL1 [0]);
  nor (_21873_, _01320_, _21872_);
  nand (_21874_, _11254_, _07958_);
  nor (_21875_, _07958_, _21872_);
  nor (_21877_, _21875_, _07217_);
  nand (_21878_, _21877_, _21874_);
  and (_21879_, _07958_, _07135_);
  or (_21880_, _21879_, _21875_);
  or (_21881_, _21880_, _06260_);
  nor (_21882_, _08374_, _11705_);
  or (_21883_, _21882_, _21875_);
  or (_21884_, _21883_, _06286_);
  and (_21885_, _07958_, \oc8051_golden_model_1.ACC [0]);
  or (_21886_, _21885_, _21875_);
  and (_21888_, _21886_, _07143_);
  nor (_21889_, _07143_, _21872_);
  or (_21890_, _21889_, _06285_);
  or (_21891_, _21890_, _21888_);
  and (_21892_, _21891_, _07169_);
  and (_21893_, _21892_, _21884_);
  and (_21894_, _21880_, _06354_);
  or (_21895_, _21894_, _21893_);
  and (_21896_, _21895_, _06346_);
  and (_21897_, _21886_, _06345_);
  or (_21899_, _21897_, _06259_);
  or (_21900_, _21899_, _21896_);
  and (_21901_, _21900_, _21881_);
  or (_21902_, _21901_, _09486_);
  and (_21903_, _09384_, _07958_);
  or (_21904_, _21875_, _06258_);
  or (_21905_, _21904_, _21903_);
  and (_21906_, _21905_, _21902_);
  or (_21907_, _21906_, _05972_);
  and (_21908_, _14413_, _07958_);
  or (_21910_, _21875_, _06251_);
  or (_21911_, _21910_, _21908_);
  and (_21912_, _21911_, _06216_);
  and (_21913_, _21912_, _21907_);
  and (_21914_, _07958_, _08929_);
  or (_21915_, _21914_, _21875_);
  and (_21916_, _21915_, _06215_);
  or (_21917_, _21916_, _06398_);
  or (_21918_, _21917_, _21913_);
  and (_21919_, _14311_, _07958_);
  or (_21921_, _21919_, _21875_);
  or (_21922_, _21921_, _09025_);
  and (_21923_, _21922_, _09030_);
  and (_21924_, _21923_, _21918_);
  nor (_21925_, _12532_, _11705_);
  or (_21926_, _21925_, _21875_);
  and (_21927_, _21874_, _06524_);
  and (_21928_, _21927_, _21926_);
  or (_21929_, _21928_, _21924_);
  and (_21930_, _21929_, _07219_);
  nand (_21932_, _21915_, _06426_);
  nor (_21933_, _21932_, _21882_);
  or (_21934_, _21933_, _06532_);
  or (_21935_, _21934_, _21930_);
  and (_21936_, _21935_, _21878_);
  or (_21937_, _21936_, _06437_);
  and (_21938_, _14307_, _07958_);
  or (_21939_, _21938_, _21875_);
  or (_21940_, _21939_, _07229_);
  and (_21941_, _21940_, _07231_);
  and (_21943_, _21941_, _21937_);
  and (_21944_, _21926_, _06535_);
  or (_21945_, _21944_, _19480_);
  or (_21946_, _21945_, _21943_);
  or (_21947_, _21883_, _06651_);
  and (_21948_, _21947_, _01320_);
  and (_21949_, _21948_, _21946_);
  or (_21950_, _21949_, _21873_);
  and (_42940_, _21950_, _42355_);
  and (_21951_, _11705_, \oc8051_golden_model_1.TL1 [1]);
  nor (_21953_, _11252_, _11705_);
  or (_21954_, _21953_, _21951_);
  or (_21955_, _21954_, _07231_);
  and (_21956_, _07958_, _09422_);
  or (_21957_, _21956_, _21951_);
  or (_21958_, _21957_, _06260_);
  or (_21959_, _07958_, \oc8051_golden_model_1.TL1 [1]);
  and (_21960_, _14520_, _07958_);
  not (_21961_, _21960_);
  and (_21962_, _21961_, _21959_);
  or (_21964_, _21962_, _06286_);
  and (_21965_, _07958_, \oc8051_golden_model_1.ACC [1]);
  or (_21966_, _21965_, _21951_);
  and (_21967_, _21966_, _07143_);
  and (_21968_, _07144_, \oc8051_golden_model_1.TL1 [1]);
  or (_21969_, _21968_, _06285_);
  or (_21970_, _21969_, _21967_);
  and (_21971_, _21970_, _07169_);
  and (_21972_, _21971_, _21964_);
  and (_21973_, _21957_, _06354_);
  or (_21975_, _21973_, _21972_);
  and (_21976_, _21975_, _06346_);
  and (_21977_, _21966_, _06345_);
  or (_21978_, _21977_, _06259_);
  or (_21979_, _21978_, _21976_);
  and (_21980_, _21979_, _21958_);
  or (_21981_, _21980_, _09486_);
  and (_21982_, _09339_, _07958_);
  or (_21983_, _21951_, _06258_);
  or (_21984_, _21983_, _21982_);
  and (_21986_, _21984_, _06251_);
  and (_21987_, _21986_, _21981_);
  or (_21988_, _14607_, _11705_);
  and (_21989_, _21959_, _05972_);
  and (_21990_, _21989_, _21988_);
  or (_21991_, _21990_, _21987_);
  and (_21992_, _21991_, _06399_);
  or (_21993_, _14505_, _11705_);
  and (_21994_, _21993_, _06398_);
  nand (_21995_, _07958_, _07031_);
  and (_21997_, _21995_, _06215_);
  or (_21998_, _21997_, _21994_);
  and (_21999_, _21998_, _21959_);
  or (_22000_, _21999_, _06524_);
  or (_22001_, _22000_, _21992_);
  nand (_22002_, _11251_, _07958_);
  and (_22003_, _22002_, _21954_);
  or (_22004_, _22003_, _09030_);
  and (_22005_, _22004_, _07219_);
  and (_22006_, _22005_, _22001_);
  or (_22008_, _14503_, _11705_);
  and (_22009_, _21959_, _06426_);
  and (_22010_, _22009_, _22008_);
  or (_22011_, _22010_, _06532_);
  or (_22012_, _22011_, _22006_);
  nor (_22013_, _21951_, _07217_);
  nand (_22014_, _22013_, _22002_);
  and (_22015_, _22014_, _07229_);
  and (_22016_, _22015_, _22012_);
  or (_22017_, _21995_, _08325_);
  and (_22019_, _21959_, _06437_);
  and (_22020_, _22019_, _22017_);
  or (_22021_, _22020_, _06535_);
  or (_22022_, _22021_, _22016_);
  and (_22023_, _22022_, _21955_);
  or (_22024_, _22023_, _06559_);
  or (_22025_, _21962_, _07240_);
  and (_22026_, _22025_, _06570_);
  and (_22027_, _22026_, _22024_);
  or (_22028_, _21960_, _21951_);
  and (_22030_, _22028_, _06566_);
  or (_22031_, _22030_, _01324_);
  or (_22032_, _22031_, _22027_);
  or (_22033_, _01320_, \oc8051_golden_model_1.TL1 [1]);
  and (_22034_, _22033_, _42355_);
  and (_42942_, _22034_, _22032_);
  and (_22035_, _01324_, \oc8051_golden_model_1.TL1 [2]);
  and (_22036_, _11705_, \oc8051_golden_model_1.TL1 [2]);
  and (_22037_, _09293_, _07958_);
  or (_22038_, _22037_, _22036_);
  and (_22040_, _22038_, _09486_);
  and (_22041_, _14703_, _07958_);
  or (_22042_, _22041_, _22036_);
  or (_22043_, _22042_, _06286_);
  and (_22044_, _07958_, \oc8051_golden_model_1.ACC [2]);
  or (_22045_, _22044_, _22036_);
  and (_22046_, _22045_, _07143_);
  and (_22047_, _07144_, \oc8051_golden_model_1.TL1 [2]);
  or (_22048_, _22047_, _06285_);
  or (_22049_, _22048_, _22046_);
  and (_22051_, _22049_, _07169_);
  and (_22052_, _22051_, _22043_);
  and (_22053_, _07958_, _08662_);
  or (_22054_, _22053_, _22036_);
  and (_22055_, _22054_, _06354_);
  or (_22056_, _22055_, _22052_);
  and (_22057_, _22056_, _06346_);
  and (_22058_, _22045_, _06345_);
  or (_22059_, _22058_, _06259_);
  or (_22060_, _22059_, _22057_);
  or (_22062_, _22054_, _06260_);
  and (_22063_, _22062_, _06258_);
  and (_22064_, _22063_, _22060_);
  or (_22065_, _22064_, _05972_);
  or (_22066_, _22065_, _22040_);
  and (_22067_, _14804_, _07958_);
  or (_22068_, _22036_, _06251_);
  or (_22069_, _22068_, _22067_);
  and (_22070_, _22069_, _06216_);
  and (_22071_, _22070_, _22066_);
  and (_22073_, _07958_, _08980_);
  or (_22074_, _22073_, _22036_);
  and (_22075_, _22074_, _06215_);
  or (_22076_, _22075_, _06398_);
  or (_22077_, _22076_, _22071_);
  and (_22078_, _14697_, _07958_);
  or (_22079_, _22078_, _22036_);
  or (_22080_, _22079_, _09025_);
  and (_22081_, _22080_, _09030_);
  and (_22082_, _22081_, _22077_);
  and (_22084_, _11250_, _07958_);
  or (_22085_, _22084_, _22036_);
  and (_22086_, _22085_, _06524_);
  or (_22087_, _22086_, _22082_);
  and (_22088_, _22087_, _07219_);
  or (_22089_, _22036_, _08424_);
  and (_22090_, _22074_, _06426_);
  and (_22091_, _22090_, _22089_);
  or (_22092_, _22091_, _22088_);
  and (_22093_, _22092_, _07217_);
  and (_22095_, _22045_, _06532_);
  and (_22096_, _22095_, _22089_);
  or (_22097_, _22096_, _06437_);
  or (_22098_, _22097_, _22093_);
  and (_22099_, _14694_, _07958_);
  or (_22100_, _22036_, _07229_);
  or (_22101_, _22100_, _22099_);
  and (_22102_, _22101_, _07231_);
  and (_22103_, _22102_, _22098_);
  nor (_22104_, _11249_, _11705_);
  or (_22106_, _22104_, _22036_);
  and (_22107_, _22106_, _06535_);
  or (_22108_, _22107_, _22103_);
  and (_22109_, _22108_, _07240_);
  and (_22110_, _22042_, _06559_);
  or (_22111_, _22110_, _06566_);
  or (_22112_, _22111_, _22109_);
  and (_22113_, _14873_, _07958_);
  or (_22114_, _22036_, _06570_);
  or (_22115_, _22114_, _22113_);
  and (_22117_, _22115_, _01320_);
  and (_22118_, _22117_, _22112_);
  or (_22119_, _22118_, _22035_);
  and (_42943_, _22119_, _42355_);
  and (_22120_, _11705_, \oc8051_golden_model_1.TL1 [3]);
  and (_22121_, _14900_, _07958_);
  or (_22122_, _22121_, _22120_);
  or (_22123_, _22122_, _06286_);
  and (_22124_, _07958_, \oc8051_golden_model_1.ACC [3]);
  or (_22125_, _22124_, _22120_);
  and (_22128_, _22125_, _07143_);
  and (_22129_, _07144_, \oc8051_golden_model_1.TL1 [3]);
  or (_22130_, _22129_, _06285_);
  or (_22131_, _22130_, _22128_);
  and (_22132_, _22131_, _07169_);
  and (_22133_, _22132_, _22123_);
  and (_22134_, _07958_, _09421_);
  or (_22135_, _22134_, _22120_);
  and (_22136_, _22135_, _06354_);
  or (_22137_, _22136_, _22133_);
  and (_22139_, _22137_, _06346_);
  and (_22140_, _22125_, _06345_);
  or (_22141_, _22140_, _06259_);
  or (_22142_, _22141_, _22139_);
  or (_22143_, _22135_, _06260_);
  and (_22144_, _22143_, _06258_);
  and (_22145_, _22144_, _22142_);
  and (_22146_, _09247_, _07958_);
  or (_22147_, _22146_, _22120_);
  and (_22148_, _22147_, _09486_);
  or (_22150_, _22148_, _05972_);
  or (_22151_, _22150_, _22145_);
  and (_22152_, _14998_, _07958_);
  or (_22153_, _22120_, _06251_);
  or (_22154_, _22153_, _22152_);
  and (_22155_, _22154_, _06216_);
  and (_22156_, _22155_, _22151_);
  and (_22157_, _07958_, _08809_);
  or (_22158_, _22157_, _22120_);
  and (_22159_, _22158_, _06215_);
  or (_22161_, _22159_, _06398_);
  or (_22162_, _22161_, _22156_);
  and (_22163_, _14893_, _07958_);
  or (_22164_, _22163_, _22120_);
  or (_22165_, _22164_, _09025_);
  and (_22166_, _22165_, _09030_);
  and (_22167_, _22166_, _22162_);
  and (_22168_, _12529_, _07958_);
  or (_22169_, _22168_, _22120_);
  and (_22170_, _22169_, _06524_);
  or (_22172_, _22170_, _22167_);
  and (_22173_, _22172_, _07219_);
  or (_22174_, _22120_, _08280_);
  and (_22175_, _22158_, _06426_);
  and (_22176_, _22175_, _22174_);
  or (_22177_, _22176_, _22173_);
  and (_22178_, _22177_, _07217_);
  and (_22179_, _22125_, _06532_);
  and (_22180_, _22179_, _22174_);
  or (_22181_, _22180_, _06437_);
  or (_22183_, _22181_, _22178_);
  and (_22184_, _14890_, _07958_);
  or (_22185_, _22120_, _07229_);
  or (_22186_, _22185_, _22184_);
  and (_22187_, _22186_, _07231_);
  and (_22188_, _22187_, _22183_);
  nor (_22189_, _11247_, _11705_);
  or (_22190_, _22189_, _22120_);
  and (_22191_, _22190_, _06535_);
  or (_22192_, _22191_, _06559_);
  or (_22194_, _22192_, _22188_);
  or (_22195_, _22122_, _07240_);
  and (_22196_, _22195_, _06570_);
  and (_22197_, _22196_, _22194_);
  and (_22198_, _15068_, _07958_);
  or (_22199_, _22198_, _22120_);
  and (_22200_, _22199_, _06566_);
  or (_22201_, _22200_, _01324_);
  or (_22202_, _22201_, _22197_);
  or (_22203_, _01320_, \oc8051_golden_model_1.TL1 [3]);
  and (_22205_, _22203_, _42355_);
  and (_42944_, _22205_, _22202_);
  and (_22206_, _11705_, \oc8051_golden_model_1.TL1 [4]);
  and (_22207_, _09420_, _07958_);
  or (_22208_, _22207_, _22206_);
  or (_22209_, _22208_, _06260_);
  and (_22210_, _15133_, _07958_);
  or (_22211_, _22210_, _22206_);
  or (_22212_, _22211_, _06286_);
  and (_22213_, _07958_, \oc8051_golden_model_1.ACC [4]);
  or (_22214_, _22213_, _22206_);
  and (_22215_, _22214_, _07143_);
  and (_22216_, _07144_, \oc8051_golden_model_1.TL1 [4]);
  or (_22217_, _22216_, _06285_);
  or (_22218_, _22217_, _22215_);
  and (_22219_, _22218_, _07169_);
  and (_22220_, _22219_, _22212_);
  and (_22221_, _22208_, _06354_);
  or (_22222_, _22221_, _22220_);
  and (_22223_, _22222_, _06346_);
  and (_22226_, _22214_, _06345_);
  or (_22227_, _22226_, _06259_);
  or (_22228_, _22227_, _22223_);
  and (_22229_, _22228_, _22209_);
  or (_22230_, _22229_, _09486_);
  and (_22231_, _09437_, _07958_);
  or (_22232_, _22206_, _06258_);
  or (_22233_, _22232_, _22231_);
  and (_22234_, _22233_, _06251_);
  and (_22235_, _22234_, _22230_);
  and (_22237_, _15226_, _07958_);
  or (_22238_, _22237_, _22206_);
  and (_22239_, _22238_, _05972_);
  or (_22240_, _22239_, _22235_);
  or (_22241_, _22240_, _10080_);
  and (_22242_, _15114_, _07958_);
  or (_22243_, _22206_, _09025_);
  or (_22244_, _22243_, _22242_);
  and (_22245_, _08919_, _07958_);
  or (_22246_, _22245_, _22206_);
  or (_22248_, _22246_, _06216_);
  and (_22249_, _22248_, _09030_);
  and (_22250_, _22249_, _22244_);
  and (_22251_, _22250_, _22241_);
  and (_22252_, _11245_, _07958_);
  or (_22253_, _22252_, _22206_);
  and (_22254_, _22253_, _06524_);
  or (_22255_, _22254_, _22251_);
  and (_22256_, _22255_, _07219_);
  or (_22257_, _22206_, _08528_);
  and (_22259_, _22246_, _06426_);
  and (_22260_, _22259_, _22257_);
  or (_22261_, _22260_, _22256_);
  and (_22262_, _22261_, _07217_);
  and (_22263_, _22214_, _06532_);
  and (_22264_, _22263_, _22257_);
  or (_22265_, _22264_, _06437_);
  or (_22266_, _22265_, _22262_);
  and (_22267_, _15111_, _07958_);
  or (_22268_, _22206_, _07229_);
  or (_22270_, _22268_, _22267_);
  and (_22271_, _22270_, _07231_);
  and (_22272_, _22271_, _22266_);
  nor (_22273_, _11244_, _11705_);
  or (_22274_, _22273_, _22206_);
  and (_22275_, _22274_, _06535_);
  or (_22276_, _22275_, _06559_);
  or (_22277_, _22276_, _22272_);
  or (_22278_, _22211_, _07240_);
  and (_22279_, _22278_, _06570_);
  and (_22281_, _22279_, _22277_);
  and (_22282_, _15296_, _07958_);
  or (_22283_, _22282_, _22206_);
  and (_22284_, _22283_, _06566_);
  or (_22285_, _22284_, _01324_);
  or (_22286_, _22285_, _22281_);
  or (_22287_, _01320_, \oc8051_golden_model_1.TL1 [4]);
  and (_22288_, _22287_, _42355_);
  and (_42945_, _22288_, _22286_);
  and (_22289_, _11705_, \oc8051_golden_model_1.TL1 [5]);
  and (_22291_, _15330_, _07958_);
  or (_22292_, _22291_, _22289_);
  or (_22293_, _22292_, _06286_);
  and (_22294_, _07958_, \oc8051_golden_model_1.ACC [5]);
  or (_22295_, _22294_, _22289_);
  and (_22296_, _22295_, _07143_);
  and (_22297_, _07144_, \oc8051_golden_model_1.TL1 [5]);
  or (_22298_, _22297_, _06285_);
  or (_22299_, _22298_, _22296_);
  and (_22300_, _22299_, _07169_);
  and (_22302_, _22300_, _22293_);
  and (_22303_, _09419_, _07958_);
  or (_22304_, _22303_, _22289_);
  and (_22305_, _22304_, _06354_);
  or (_22306_, _22305_, _22302_);
  and (_22307_, _22306_, _06346_);
  and (_22308_, _22295_, _06345_);
  or (_22309_, _22308_, _06259_);
  or (_22310_, _22309_, _22307_);
  or (_22311_, _22304_, _06260_);
  and (_22313_, _22311_, _22310_);
  or (_22314_, _22313_, _09486_);
  and (_22315_, _09436_, _07958_);
  or (_22316_, _22289_, _06258_);
  or (_22317_, _22316_, _22315_);
  and (_22318_, _22317_, _06251_);
  and (_22319_, _22318_, _22314_);
  and (_22320_, _15421_, _07958_);
  or (_22321_, _22320_, _22289_);
  and (_22322_, _22321_, _05972_);
  or (_22324_, _22322_, _10080_);
  or (_22325_, _22324_, _22319_);
  and (_22326_, _15313_, _07958_);
  or (_22327_, _22289_, _09025_);
  or (_22328_, _22327_, _22326_);
  and (_22329_, _08913_, _07958_);
  or (_22330_, _22329_, _22289_);
  or (_22331_, _22330_, _06216_);
  and (_22332_, _22331_, _09030_);
  and (_22333_, _22332_, _22328_);
  and (_22335_, _22333_, _22325_);
  and (_22336_, _12536_, _07958_);
  or (_22337_, _22336_, _22289_);
  and (_22338_, _22337_, _06524_);
  or (_22339_, _22338_, _22335_);
  and (_22340_, _22339_, _07219_);
  or (_22341_, _22289_, _08231_);
  and (_22342_, _22330_, _06426_);
  and (_22343_, _22342_, _22341_);
  or (_22344_, _22343_, _22340_);
  and (_22346_, _22344_, _07217_);
  and (_22347_, _22295_, _06532_);
  and (_22348_, _22347_, _22341_);
  or (_22349_, _22348_, _06437_);
  or (_22350_, _22349_, _22346_);
  and (_22351_, _15310_, _07958_);
  or (_22352_, _22289_, _07229_);
  or (_22353_, _22352_, _22351_);
  and (_22354_, _22353_, _07231_);
  and (_22355_, _22354_, _22350_);
  nor (_22357_, _11241_, _11705_);
  or (_22358_, _22357_, _22289_);
  and (_22359_, _22358_, _06535_);
  or (_22360_, _22359_, _06559_);
  or (_22361_, _22360_, _22355_);
  or (_22362_, _22292_, _07240_);
  and (_22363_, _22362_, _06570_);
  and (_22364_, _22363_, _22361_);
  and (_22365_, _15493_, _07958_);
  or (_22366_, _22365_, _22289_);
  and (_22368_, _22366_, _06566_);
  or (_22369_, _22368_, _01324_);
  or (_22370_, _22369_, _22364_);
  or (_22371_, _01320_, \oc8051_golden_model_1.TL1 [5]);
  and (_22372_, _22371_, _42355_);
  and (_42946_, _22372_, _22370_);
  and (_22373_, _11705_, \oc8051_golden_model_1.TL1 [6]);
  and (_22374_, _15521_, _07958_);
  or (_22375_, _22374_, _22373_);
  or (_22376_, _22375_, _06286_);
  and (_22378_, _07958_, \oc8051_golden_model_1.ACC [6]);
  or (_22379_, _22378_, _22373_);
  and (_22380_, _22379_, _07143_);
  and (_22381_, _07144_, \oc8051_golden_model_1.TL1 [6]);
  or (_22382_, _22381_, _06285_);
  or (_22383_, _22382_, _22380_);
  and (_22384_, _22383_, _07169_);
  and (_22385_, _22384_, _22376_);
  and (_22386_, _09418_, _07958_);
  or (_22387_, _22386_, _22373_);
  and (_22389_, _22387_, _06354_);
  or (_22390_, _22389_, _22385_);
  and (_22391_, _22390_, _06346_);
  and (_22392_, _22379_, _06345_);
  or (_22393_, _22392_, _06259_);
  or (_22394_, _22393_, _22391_);
  or (_22395_, _22387_, _06260_);
  and (_22396_, _22395_, _22394_);
  or (_22397_, _22396_, _09486_);
  and (_22398_, _09435_, _07958_);
  or (_22400_, _22373_, _06258_);
  or (_22401_, _22400_, _22398_);
  and (_22402_, _22401_, _06251_);
  and (_22403_, _22402_, _22397_);
  and (_22404_, _15623_, _07958_);
  or (_22405_, _22404_, _22373_);
  and (_22406_, _22405_, _05972_);
  or (_22407_, _22406_, _10080_);
  or (_22408_, _22407_, _22403_);
  and (_22409_, _15517_, _07958_);
  or (_22411_, _22373_, _09025_);
  or (_22412_, _22411_, _22409_);
  and (_22413_, _08845_, _07958_);
  or (_22414_, _22413_, _22373_);
  or (_22415_, _22414_, _06216_);
  and (_22416_, _22415_, _09030_);
  and (_22417_, _22416_, _22412_);
  and (_22418_, _22417_, _22408_);
  and (_22419_, _11239_, _07958_);
  or (_22420_, _22419_, _22373_);
  and (_22422_, _22420_, _06524_);
  or (_22423_, _22422_, _22418_);
  and (_22424_, _22423_, _07219_);
  or (_22425_, _22373_, _08128_);
  and (_22426_, _22414_, _06426_);
  and (_22427_, _22426_, _22425_);
  or (_22428_, _22427_, _22424_);
  and (_22429_, _22428_, _07217_);
  and (_22430_, _22379_, _06532_);
  and (_22431_, _22430_, _22425_);
  or (_22433_, _22431_, _06437_);
  or (_22434_, _22433_, _22429_);
  and (_22435_, _15514_, _07958_);
  or (_22436_, _22373_, _07229_);
  or (_22437_, _22436_, _22435_);
  and (_22438_, _22437_, _07231_);
  and (_22439_, _22438_, _22434_);
  nor (_22440_, _11238_, _11705_);
  or (_22441_, _22440_, _22373_);
  and (_22442_, _22441_, _06535_);
  or (_22444_, _22442_, _06559_);
  or (_22445_, _22444_, _22439_);
  or (_22446_, _22375_, _07240_);
  and (_22447_, _22446_, _06570_);
  and (_22448_, _22447_, _22445_);
  and (_22449_, _15695_, _07958_);
  or (_22450_, _22449_, _22373_);
  and (_22451_, _22450_, _06566_);
  or (_22452_, _22451_, _01324_);
  or (_22453_, _22452_, _22448_);
  or (_22455_, _01320_, \oc8051_golden_model_1.TL1 [6]);
  and (_22456_, _22455_, _42355_);
  and (_42947_, _22456_, _22453_);
  not (_22457_, \oc8051_golden_model_1.TL0 [0]);
  nor (_22458_, _01320_, _22457_);
  nand (_22459_, _11254_, _07912_);
  nor (_22460_, _07912_, _22457_);
  nor (_22461_, _22460_, _07217_);
  nand (_22462_, _22461_, _22459_);
  and (_22463_, _07912_, \oc8051_golden_model_1.ACC [0]);
  or (_22465_, _22463_, _22460_);
  and (_22466_, _22465_, _06345_);
  or (_22467_, _22466_, _06259_);
  nor (_22468_, _08374_, _11782_);
  or (_22469_, _22468_, _22460_);
  and (_22470_, _22469_, _06285_);
  nor (_22471_, _07143_, _22457_);
  and (_22472_, _22465_, _07143_);
  or (_22473_, _22472_, _22471_);
  and (_22474_, _22473_, _06286_);
  or (_22476_, _22474_, _06354_);
  or (_22477_, _22476_, _22470_);
  and (_22478_, _22477_, _06346_);
  or (_22479_, _22478_, _22467_);
  and (_22480_, _07912_, _07135_);
  or (_22481_, _22460_, _19434_);
  or (_22482_, _22481_, _22480_);
  and (_22483_, _22482_, _22479_);
  or (_22484_, _22483_, _09486_);
  and (_22485_, _09384_, _07912_);
  or (_22487_, _22460_, _06258_);
  or (_22488_, _22487_, _22485_);
  and (_22489_, _22488_, _22484_);
  or (_22490_, _22489_, _05972_);
  and (_22491_, _14413_, _07912_);
  or (_22492_, _22460_, _06251_);
  or (_22493_, _22492_, _22491_);
  and (_22494_, _22493_, _06216_);
  and (_22495_, _22494_, _22490_);
  and (_22496_, _07912_, _08929_);
  or (_22498_, _22496_, _22460_);
  and (_22499_, _22498_, _06215_);
  or (_22500_, _22499_, _06398_);
  or (_22501_, _22500_, _22495_);
  and (_22502_, _14311_, _07912_);
  or (_22503_, _22502_, _22460_);
  or (_22504_, _22503_, _09025_);
  and (_22505_, _22504_, _09030_);
  and (_22506_, _22505_, _22501_);
  nor (_22507_, _12532_, _11782_);
  or (_22508_, _22507_, _22460_);
  and (_22509_, _22459_, _06524_);
  and (_22510_, _22509_, _22508_);
  or (_22511_, _22510_, _22506_);
  and (_22512_, _22511_, _07219_);
  nand (_22513_, _22498_, _06426_);
  nor (_22514_, _22513_, _22468_);
  or (_22515_, _22514_, _06532_);
  or (_22516_, _22515_, _22512_);
  and (_22517_, _22516_, _22462_);
  or (_22520_, _22517_, _06437_);
  and (_22521_, _14307_, _07912_);
  or (_22522_, _22460_, _07229_);
  or (_22523_, _22522_, _22521_);
  and (_22524_, _22523_, _07231_);
  and (_22525_, _22524_, _22520_);
  and (_22526_, _22508_, _06535_);
  or (_22527_, _22526_, _19480_);
  or (_22528_, _22527_, _22525_);
  or (_22529_, _22469_, _06651_);
  and (_22531_, _22529_, _01320_);
  and (_22532_, _22531_, _22528_);
  or (_22533_, _22532_, _22458_);
  and (_42949_, _22533_, _42355_);
  and (_22534_, _11782_, \oc8051_golden_model_1.TL0 [1]);
  nor (_22535_, _11252_, _11782_);
  or (_22536_, _22535_, _22534_);
  or (_22537_, _22536_, _07231_);
  or (_22538_, _07912_, \oc8051_golden_model_1.TL0 [1]);
  and (_22539_, _14520_, _07912_);
  not (_22541_, _22539_);
  and (_22542_, _22541_, _22538_);
  or (_22543_, _22542_, _06286_);
  and (_22544_, _07912_, \oc8051_golden_model_1.ACC [1]);
  or (_22545_, _22544_, _22534_);
  and (_22546_, _22545_, _07143_);
  and (_22547_, _07144_, \oc8051_golden_model_1.TL0 [1]);
  or (_22548_, _22547_, _06285_);
  or (_22549_, _22548_, _22546_);
  and (_22550_, _22549_, _07169_);
  and (_22552_, _22550_, _22543_);
  and (_22553_, _07912_, _09422_);
  or (_22554_, _22553_, _22534_);
  and (_22555_, _22554_, _06354_);
  or (_22556_, _22555_, _22552_);
  and (_22557_, _22556_, _06346_);
  and (_22558_, _22545_, _06345_);
  or (_22559_, _22558_, _06259_);
  or (_22560_, _22559_, _22557_);
  or (_22561_, _22554_, _06260_);
  and (_22563_, _22561_, _22560_);
  or (_22564_, _22563_, _09486_);
  and (_22565_, _09339_, _07912_);
  or (_22566_, _22534_, _06258_);
  or (_22567_, _22566_, _22565_);
  and (_22568_, _22567_, _06251_);
  and (_22569_, _22568_, _22564_);
  or (_22570_, _14607_, _11782_);
  and (_22571_, _22538_, _05972_);
  and (_22572_, _22571_, _22570_);
  or (_22574_, _22572_, _22569_);
  and (_22575_, _22574_, _06399_);
  or (_22576_, _14505_, _11782_);
  and (_22577_, _22576_, _06398_);
  nand (_22578_, _07912_, _07031_);
  and (_22579_, _22578_, _06215_);
  or (_22580_, _22579_, _22577_);
  and (_22581_, _22580_, _22538_);
  or (_22582_, _22581_, _06524_);
  or (_22583_, _22582_, _22575_);
  nand (_22585_, _11251_, _07912_);
  and (_22586_, _22585_, _22536_);
  or (_22587_, _22586_, _09030_);
  and (_22588_, _22587_, _07219_);
  and (_22589_, _22588_, _22583_);
  or (_22590_, _14503_, _11782_);
  and (_22591_, _22538_, _06426_);
  and (_22592_, _22591_, _22590_);
  or (_22593_, _22592_, _06532_);
  or (_22594_, _22593_, _22589_);
  nor (_22596_, _22534_, _07217_);
  nand (_22597_, _22596_, _22585_);
  and (_22598_, _22597_, _07229_);
  and (_22599_, _22598_, _22594_);
  or (_22600_, _22578_, _08325_);
  and (_22601_, _22538_, _06437_);
  and (_22602_, _22601_, _22600_);
  or (_22603_, _22602_, _06535_);
  or (_22604_, _22603_, _22599_);
  and (_22605_, _22604_, _22537_);
  or (_22607_, _22605_, _06559_);
  or (_22608_, _22542_, _07240_);
  and (_22609_, _22608_, _06570_);
  and (_22610_, _22609_, _22607_);
  or (_22611_, _22539_, _22534_);
  and (_22612_, _22611_, _06566_);
  or (_22613_, _22612_, _01324_);
  or (_22614_, _22613_, _22610_);
  or (_22615_, _01320_, \oc8051_golden_model_1.TL0 [1]);
  and (_22616_, _22615_, _42355_);
  and (_42950_, _22616_, _22614_);
  and (_22617_, _01324_, \oc8051_golden_model_1.TL0 [2]);
  and (_22618_, _11782_, \oc8051_golden_model_1.TL0 [2]);
  and (_22619_, _09293_, _07912_);
  or (_22620_, _22619_, _22618_);
  and (_22621_, _22620_, _09486_);
  and (_22622_, _14703_, _07912_);
  or (_22623_, _22622_, _22618_);
  or (_22624_, _22623_, _06286_);
  and (_22625_, _07912_, \oc8051_golden_model_1.ACC [2]);
  or (_22628_, _22625_, _22618_);
  and (_22629_, _22628_, _07143_);
  and (_22630_, _07144_, \oc8051_golden_model_1.TL0 [2]);
  or (_22631_, _22630_, _06285_);
  or (_22632_, _22631_, _22629_);
  and (_22633_, _22632_, _07169_);
  and (_22634_, _22633_, _22624_);
  and (_22635_, _07912_, _08662_);
  or (_22636_, _22635_, _22618_);
  and (_22637_, _22636_, _06354_);
  or (_22639_, _22637_, _22634_);
  and (_22640_, _22639_, _06346_);
  and (_22641_, _22628_, _06345_);
  or (_22642_, _22641_, _06259_);
  or (_22643_, _22642_, _22640_);
  or (_22644_, _22636_, _06260_);
  and (_22645_, _22644_, _06258_);
  and (_22646_, _22645_, _22643_);
  or (_22647_, _22646_, _05972_);
  or (_22648_, _22647_, _22621_);
  and (_22650_, _14804_, _07912_);
  or (_22651_, _22618_, _06251_);
  or (_22652_, _22651_, _22650_);
  and (_22653_, _22652_, _06216_);
  and (_22654_, _22653_, _22648_);
  and (_22655_, _07912_, _08980_);
  or (_22656_, _22655_, _22618_);
  and (_22657_, _22656_, _06215_);
  or (_22658_, _22657_, _06398_);
  or (_22659_, _22658_, _22654_);
  and (_22661_, _14697_, _07912_);
  or (_22662_, _22661_, _22618_);
  or (_22663_, _22662_, _09025_);
  and (_22664_, _22663_, _09030_);
  and (_22665_, _22664_, _22659_);
  and (_22666_, _11250_, _07912_);
  or (_22667_, _22666_, _22618_);
  and (_22668_, _22667_, _06524_);
  or (_22669_, _22668_, _22665_);
  and (_22670_, _22669_, _07219_);
  or (_22672_, _22618_, _08424_);
  and (_22673_, _22656_, _06426_);
  and (_22674_, _22673_, _22672_);
  or (_22675_, _22674_, _22670_);
  and (_22676_, _22675_, _07217_);
  and (_22677_, _22628_, _06532_);
  and (_22678_, _22677_, _22672_);
  or (_22679_, _22678_, _06437_);
  or (_22680_, _22679_, _22676_);
  and (_22681_, _14694_, _07912_);
  or (_22683_, _22618_, _07229_);
  or (_22684_, _22683_, _22681_);
  and (_22685_, _22684_, _07231_);
  and (_22686_, _22685_, _22680_);
  nor (_22687_, _11249_, _11782_);
  or (_22688_, _22687_, _22618_);
  and (_22689_, _22688_, _06535_);
  or (_22690_, _22689_, _22686_);
  and (_22691_, _22690_, _07240_);
  and (_22692_, _22623_, _06559_);
  or (_22694_, _22692_, _06566_);
  or (_22695_, _22694_, _22691_);
  and (_22696_, _14873_, _07912_);
  or (_22697_, _22618_, _06570_);
  or (_22698_, _22697_, _22696_);
  and (_22699_, _22698_, _01320_);
  and (_22700_, _22699_, _22695_);
  or (_22701_, _22700_, _22617_);
  and (_42951_, _22701_, _42355_);
  and (_22702_, _11782_, \oc8051_golden_model_1.TL0 [3]);
  and (_22704_, _14900_, _07912_);
  or (_22705_, _22704_, _22702_);
  or (_22706_, _22705_, _06286_);
  and (_22707_, _07912_, \oc8051_golden_model_1.ACC [3]);
  or (_22708_, _22707_, _22702_);
  and (_22709_, _22708_, _07143_);
  and (_22710_, _07144_, \oc8051_golden_model_1.TL0 [3]);
  or (_22711_, _22710_, _06285_);
  or (_22712_, _22711_, _22709_);
  and (_22713_, _22712_, _07169_);
  and (_22715_, _22713_, _22706_);
  and (_22716_, _07912_, _09421_);
  or (_22717_, _22716_, _22702_);
  and (_22718_, _22717_, _06354_);
  or (_22719_, _22718_, _22715_);
  and (_22720_, _22719_, _06346_);
  and (_22721_, _22708_, _06345_);
  or (_22722_, _22721_, _06259_);
  or (_22723_, _22722_, _22720_);
  or (_22724_, _22717_, _06260_);
  and (_22726_, _22724_, _22723_);
  or (_22727_, _22726_, _09486_);
  and (_22728_, _09247_, _07912_);
  or (_22729_, _22702_, _06258_);
  or (_22730_, _22729_, _22728_);
  and (_22731_, _22730_, _06251_);
  and (_22732_, _22731_, _22727_);
  and (_22733_, _14998_, _07912_);
  or (_22734_, _22733_, _22702_);
  and (_22735_, _22734_, _05972_);
  or (_22737_, _22735_, _10080_);
  or (_22738_, _22737_, _22732_);
  and (_22739_, _14893_, _07912_);
  or (_22740_, _22702_, _09025_);
  or (_22741_, _22740_, _22739_);
  and (_22742_, _07912_, _08809_);
  or (_22743_, _22742_, _22702_);
  or (_22744_, _22743_, _06216_);
  and (_22745_, _22744_, _09030_);
  and (_22746_, _22745_, _22741_);
  and (_22748_, _22746_, _22738_);
  and (_22749_, _12529_, _07912_);
  or (_22750_, _22749_, _22702_);
  and (_22751_, _22750_, _06524_);
  or (_22752_, _22751_, _22748_);
  and (_22753_, _22752_, _07219_);
  or (_22754_, _22702_, _08280_);
  and (_22755_, _22743_, _06426_);
  and (_22756_, _22755_, _22754_);
  or (_22757_, _22756_, _22753_);
  and (_22759_, _22757_, _07217_);
  and (_22760_, _22708_, _06532_);
  and (_22761_, _22760_, _22754_);
  or (_22762_, _22761_, _06437_);
  or (_22763_, _22762_, _22759_);
  and (_22764_, _14890_, _07912_);
  or (_22765_, _22702_, _07229_);
  or (_22766_, _22765_, _22764_);
  and (_22767_, _22766_, _07231_);
  and (_22768_, _22767_, _22763_);
  nor (_22770_, _11247_, _11782_);
  or (_22771_, _22770_, _22702_);
  and (_22772_, _22771_, _06535_);
  or (_22773_, _22772_, _06559_);
  or (_22774_, _22773_, _22768_);
  or (_22775_, _22705_, _07240_);
  and (_22776_, _22775_, _06570_);
  and (_22777_, _22776_, _22774_);
  and (_22778_, _15068_, _07912_);
  or (_22779_, _22778_, _22702_);
  and (_22781_, _22779_, _06566_);
  or (_22782_, _22781_, _01324_);
  or (_22783_, _22782_, _22777_);
  or (_22784_, _01320_, \oc8051_golden_model_1.TL0 [3]);
  and (_22785_, _22784_, _42355_);
  and (_42952_, _22785_, _22783_);
  and (_22786_, _11782_, \oc8051_golden_model_1.TL0 [4]);
  and (_22787_, _15133_, _07912_);
  or (_22788_, _22787_, _22786_);
  or (_22789_, _22788_, _06286_);
  and (_22791_, _07912_, \oc8051_golden_model_1.ACC [4]);
  or (_22792_, _22791_, _22786_);
  and (_22793_, _22792_, _07143_);
  and (_22794_, _07144_, \oc8051_golden_model_1.TL0 [4]);
  or (_22795_, _22794_, _06285_);
  or (_22796_, _22795_, _22793_);
  and (_22797_, _22796_, _07169_);
  and (_22798_, _22797_, _22789_);
  and (_22799_, _09420_, _07912_);
  or (_22800_, _22799_, _22786_);
  and (_22802_, _22800_, _06354_);
  or (_22803_, _22802_, _22798_);
  and (_22804_, _22803_, _06346_);
  and (_22805_, _22792_, _06345_);
  or (_22806_, _22805_, _06259_);
  or (_22807_, _22806_, _22804_);
  or (_22808_, _22800_, _06260_);
  and (_22809_, _22808_, _22807_);
  or (_22810_, _22809_, _09486_);
  and (_22811_, _09437_, _07912_);
  or (_22813_, _22786_, _06258_);
  or (_22814_, _22813_, _22811_);
  and (_22815_, _22814_, _06251_);
  and (_22816_, _22815_, _22810_);
  and (_22817_, _15226_, _07912_);
  or (_22818_, _22817_, _22786_);
  and (_22819_, _22818_, _05972_);
  or (_22820_, _22819_, _22816_);
  or (_22821_, _22820_, _10080_);
  and (_22822_, _15114_, _07912_);
  or (_22824_, _22786_, _09025_);
  or (_22825_, _22824_, _22822_);
  and (_22826_, _08919_, _07912_);
  or (_22827_, _22826_, _22786_);
  or (_22828_, _22827_, _06216_);
  and (_22829_, _22828_, _09030_);
  and (_22830_, _22829_, _22825_);
  and (_22831_, _22830_, _22821_);
  and (_22832_, _11245_, _07912_);
  or (_22833_, _22832_, _22786_);
  and (_22834_, _22833_, _06524_);
  or (_22835_, _22834_, _22831_);
  and (_22836_, _22835_, _07219_);
  or (_22837_, _22786_, _08528_);
  and (_22838_, _22827_, _06426_);
  and (_22839_, _22838_, _22837_);
  or (_22840_, _22839_, _22836_);
  and (_22841_, _22840_, _07217_);
  and (_22842_, _22792_, _06532_);
  and (_22843_, _22842_, _22837_);
  or (_22846_, _22843_, _06437_);
  or (_22847_, _22846_, _22841_);
  and (_22848_, _15111_, _07912_);
  or (_22849_, _22786_, _07229_);
  or (_22850_, _22849_, _22848_);
  and (_22851_, _22850_, _07231_);
  and (_22852_, _22851_, _22847_);
  nor (_22853_, _11244_, _11782_);
  or (_22854_, _22853_, _22786_);
  and (_22855_, _22854_, _06535_);
  or (_22857_, _22855_, _06559_);
  or (_22858_, _22857_, _22852_);
  or (_22859_, _22788_, _07240_);
  and (_22860_, _22859_, _06570_);
  and (_22861_, _22860_, _22858_);
  and (_22862_, _15296_, _07912_);
  or (_22863_, _22862_, _22786_);
  and (_22864_, _22863_, _06566_);
  or (_22865_, _22864_, _01324_);
  or (_22866_, _22865_, _22861_);
  or (_22868_, _01320_, \oc8051_golden_model_1.TL0 [4]);
  and (_22869_, _22868_, _42355_);
  and (_42953_, _22869_, _22866_);
  and (_22870_, _11782_, \oc8051_golden_model_1.TL0 [5]);
  and (_22871_, _15330_, _07912_);
  or (_22872_, _22871_, _22870_);
  or (_22873_, _22872_, _06286_);
  and (_22874_, _07912_, \oc8051_golden_model_1.ACC [5]);
  or (_22875_, _22874_, _22870_);
  and (_22876_, _22875_, _07143_);
  and (_22878_, _07144_, \oc8051_golden_model_1.TL0 [5]);
  or (_22879_, _22878_, _06285_);
  or (_22880_, _22879_, _22876_);
  and (_22881_, _22880_, _07169_);
  and (_22882_, _22881_, _22873_);
  and (_22883_, _09419_, _07912_);
  or (_22884_, _22883_, _22870_);
  and (_22885_, _22884_, _06354_);
  or (_22886_, _22885_, _22882_);
  and (_22887_, _22886_, _06346_);
  and (_22889_, _22875_, _06345_);
  or (_22890_, _22889_, _06259_);
  or (_22891_, _22890_, _22887_);
  or (_22892_, _22884_, _06260_);
  and (_22893_, _22892_, _22891_);
  or (_22894_, _22893_, _09486_);
  and (_22895_, _09436_, _07912_);
  or (_22896_, _22870_, _06258_);
  or (_22897_, _22896_, _22895_);
  and (_22898_, _22897_, _06251_);
  and (_22900_, _22898_, _22894_);
  and (_22901_, _15421_, _07912_);
  or (_22902_, _22901_, _22870_);
  and (_22903_, _22902_, _05972_);
  or (_22904_, _22903_, _10080_);
  or (_22905_, _22904_, _22900_);
  and (_22906_, _15313_, _07912_);
  or (_22907_, _22870_, _09025_);
  or (_22908_, _22907_, _22906_);
  and (_22909_, _08913_, _07912_);
  or (_22911_, _22909_, _22870_);
  or (_22912_, _22911_, _06216_);
  and (_22913_, _22912_, _09030_);
  and (_22914_, _22913_, _22908_);
  and (_22915_, _22914_, _22905_);
  and (_22916_, _12536_, _07912_);
  or (_22917_, _22916_, _22870_);
  and (_22918_, _22917_, _06524_);
  or (_22919_, _22918_, _22915_);
  and (_22920_, _22919_, _07219_);
  or (_22922_, _22870_, _08231_);
  and (_22923_, _22911_, _06426_);
  and (_22924_, _22923_, _22922_);
  or (_22925_, _22924_, _22920_);
  and (_22926_, _22925_, _07217_);
  and (_22927_, _22875_, _06532_);
  and (_22928_, _22927_, _22922_);
  or (_22929_, _22928_, _06437_);
  or (_22930_, _22929_, _22926_);
  and (_22931_, _15310_, _07912_);
  or (_22933_, _22870_, _07229_);
  or (_22934_, _22933_, _22931_);
  and (_22935_, _22934_, _07231_);
  and (_22936_, _22935_, _22930_);
  nor (_22937_, _11241_, _11782_);
  or (_22938_, _22937_, _22870_);
  and (_22939_, _22938_, _06535_);
  or (_22940_, _22939_, _06559_);
  or (_22941_, _22940_, _22936_);
  or (_22942_, _22872_, _07240_);
  and (_22944_, _22942_, _06570_);
  and (_22945_, _22944_, _22941_);
  and (_22946_, _15493_, _07912_);
  or (_22947_, _22946_, _22870_);
  and (_22948_, _22947_, _06566_);
  or (_22949_, _22948_, _01324_);
  or (_22950_, _22949_, _22945_);
  or (_22951_, _01320_, \oc8051_golden_model_1.TL0 [5]);
  and (_22952_, _22951_, _42355_);
  and (_42954_, _22952_, _22950_);
  and (_22954_, _11782_, \oc8051_golden_model_1.TL0 [6]);
  and (_22955_, _15521_, _07912_);
  or (_22956_, _22955_, _22954_);
  or (_22957_, _22956_, _06286_);
  and (_22958_, _07912_, \oc8051_golden_model_1.ACC [6]);
  or (_22959_, _22958_, _22954_);
  and (_22960_, _22959_, _07143_);
  and (_22961_, _07144_, \oc8051_golden_model_1.TL0 [6]);
  or (_22962_, _22961_, _06285_);
  or (_22963_, _22962_, _22960_);
  and (_22965_, _22963_, _07169_);
  and (_22966_, _22965_, _22957_);
  and (_22967_, _09418_, _07912_);
  or (_22968_, _22967_, _22954_);
  and (_22969_, _22968_, _06354_);
  or (_22970_, _22969_, _22966_);
  and (_22971_, _22970_, _06346_);
  and (_22972_, _22959_, _06345_);
  or (_22973_, _22972_, _06259_);
  or (_22974_, _22973_, _22971_);
  or (_22976_, _22968_, _06260_);
  and (_22977_, _22976_, _22974_);
  or (_22978_, _22977_, _09486_);
  and (_22979_, _09435_, _07912_);
  or (_22980_, _22954_, _06258_);
  or (_22981_, _22980_, _22979_);
  and (_22982_, _22981_, _06251_);
  and (_22983_, _22982_, _22978_);
  and (_22984_, _15623_, _07912_);
  or (_22985_, _22984_, _22954_);
  and (_22987_, _22985_, _05972_);
  or (_22988_, _22987_, _10080_);
  or (_22989_, _22988_, _22983_);
  and (_22990_, _15517_, _07912_);
  or (_22991_, _22954_, _09025_);
  or (_22992_, _22991_, _22990_);
  and (_22993_, _08845_, _07912_);
  or (_22994_, _22993_, _22954_);
  or (_22995_, _22994_, _06216_);
  and (_22996_, _22995_, _09030_);
  and (_22998_, _22996_, _22992_);
  and (_22999_, _22998_, _22989_);
  and (_23000_, _11239_, _07912_);
  or (_23001_, _23000_, _22954_);
  and (_23002_, _23001_, _06524_);
  or (_23003_, _23002_, _22999_);
  and (_23004_, _23003_, _07219_);
  or (_23005_, _22954_, _08128_);
  and (_23006_, _22994_, _06426_);
  and (_23007_, _23006_, _23005_);
  or (_23009_, _23007_, _23004_);
  and (_23010_, _23009_, _07217_);
  and (_23011_, _22959_, _06532_);
  and (_23012_, _23011_, _23005_);
  or (_23013_, _23012_, _06437_);
  or (_23014_, _23013_, _23010_);
  and (_23015_, _15514_, _07912_);
  or (_23016_, _22954_, _07229_);
  or (_23017_, _23016_, _23015_);
  and (_23018_, _23017_, _07231_);
  and (_23020_, _23018_, _23014_);
  nor (_23021_, _11238_, _11782_);
  or (_23022_, _23021_, _22954_);
  and (_23023_, _23022_, _06535_);
  or (_23024_, _23023_, _06559_);
  or (_23025_, _23024_, _23020_);
  or (_23026_, _22956_, _07240_);
  and (_23027_, _23026_, _06570_);
  and (_23028_, _23027_, _23025_);
  and (_23029_, _15695_, _07912_);
  or (_23031_, _23029_, _22954_);
  and (_23032_, _23031_, _06566_);
  or (_23033_, _23032_, _01324_);
  or (_23034_, _23033_, _23028_);
  or (_23035_, _01320_, \oc8051_golden_model_1.TL0 [6]);
  and (_23036_, _23035_, _42355_);
  and (_42955_, _23036_, _23034_);
  not (_23037_, \oc8051_golden_model_1.TCON [0]);
  nor (_23038_, _01320_, _23037_);
  nand (_23039_, _11254_, _07916_);
  nor (_23041_, _07916_, _23037_);
  nor (_23042_, _23041_, _07217_);
  nand (_23043_, _23042_, _23039_);
  and (_23044_, _07916_, _07135_);
  or (_23045_, _23044_, _23041_);
  or (_23046_, _23045_, _06260_);
  nor (_23047_, _08374_, _11860_);
  or (_23048_, _23047_, _23041_);
  or (_23049_, _23048_, _06286_);
  and (_23050_, _07916_, \oc8051_golden_model_1.ACC [0]);
  or (_23052_, _23050_, _23041_);
  and (_23053_, _23052_, _07143_);
  nor (_23054_, _07143_, _23037_);
  or (_23055_, _23054_, _06285_);
  or (_23056_, _23055_, _23053_);
  and (_23057_, _23056_, _06282_);
  and (_23058_, _23057_, _23049_);
  nor (_23059_, _08600_, _23037_);
  and (_23060_, _14326_, _08600_);
  or (_23061_, _23060_, _23059_);
  and (_23063_, _23061_, _06281_);
  or (_23064_, _23063_, _23058_);
  and (_23065_, _23064_, _07169_);
  and (_23066_, _23045_, _06354_);
  or (_23067_, _23066_, _06345_);
  or (_23068_, _23067_, _23065_);
  or (_23069_, _23052_, _06346_);
  and (_23070_, _23069_, _06278_);
  and (_23071_, _23070_, _23068_);
  and (_23072_, _23041_, _06277_);
  or (_23074_, _23072_, _06270_);
  or (_23075_, _23074_, _23071_);
  or (_23076_, _23048_, _06271_);
  and (_23077_, _23076_, _06267_);
  and (_23078_, _23077_, _23075_);
  and (_23079_, _14358_, _08600_);
  or (_23080_, _23079_, _23059_);
  and (_23081_, _23080_, _06266_);
  or (_23082_, _23081_, _06259_);
  or (_23083_, _23082_, _23078_);
  and (_23085_, _23083_, _23046_);
  or (_23086_, _23085_, _09486_);
  and (_23087_, _09384_, _07916_);
  or (_23088_, _23041_, _06258_);
  or (_23089_, _23088_, _23087_);
  and (_23090_, _23089_, _06251_);
  and (_23091_, _23090_, _23086_);
  and (_23092_, _14413_, _07916_);
  or (_23093_, _23092_, _23041_);
  and (_23094_, _23093_, _05972_);
  or (_23095_, _23094_, _23091_);
  or (_23096_, _23095_, _10080_);
  and (_23097_, _14311_, _07916_);
  or (_23098_, _23041_, _09025_);
  or (_23099_, _23098_, _23097_);
  and (_23100_, _07916_, _08929_);
  or (_23101_, _23100_, _23041_);
  or (_23102_, _23101_, _06216_);
  and (_23103_, _23102_, _09030_);
  and (_23104_, _23103_, _23099_);
  and (_23107_, _23104_, _23096_);
  nor (_23108_, _12532_, _11860_);
  or (_23109_, _23108_, _23041_);
  and (_23110_, _23039_, _06524_);
  and (_23111_, _23110_, _23109_);
  or (_23112_, _23111_, _23107_);
  and (_23113_, _23112_, _07219_);
  nand (_23114_, _23101_, _06426_);
  nor (_23115_, _23114_, _23047_);
  or (_23116_, _23115_, _06532_);
  or (_23118_, _23116_, _23113_);
  and (_23119_, _23118_, _23043_);
  or (_23120_, _23119_, _06437_);
  and (_23121_, _14307_, _07916_);
  or (_23122_, _23041_, _07229_);
  or (_23123_, _23122_, _23121_);
  and (_23124_, _23123_, _07231_);
  and (_23125_, _23124_, _23120_);
  and (_23126_, _23109_, _06535_);
  or (_23127_, _23126_, _06559_);
  or (_23129_, _23127_, _23125_);
  or (_23130_, _23048_, _07240_);
  and (_23131_, _23130_, _23129_);
  or (_23132_, _23131_, _05932_);
  or (_23133_, _23041_, _05933_);
  and (_23134_, _23133_, _23132_);
  or (_23135_, _23134_, _06566_);
  or (_23136_, _23048_, _06570_);
  and (_23137_, _23136_, _01320_);
  and (_23138_, _23137_, _23135_);
  or (_23140_, _23138_, _23038_);
  and (_42957_, _23140_, _42355_);
  not (_23141_, \oc8051_golden_model_1.TCON [1]);
  nor (_23142_, _01320_, _23141_);
  nor (_23143_, _07916_, _23141_);
  nor (_23144_, _11252_, _11860_);
  or (_23145_, _23144_, _23143_);
  or (_23146_, _23145_, _07231_);
  and (_23147_, _07916_, _09422_);
  or (_23148_, _23147_, _23143_);
  or (_23150_, _23148_, _07169_);
  or (_23151_, _07916_, \oc8051_golden_model_1.TCON [1]);
  and (_23152_, _14520_, _07916_);
  not (_23153_, _23152_);
  and (_23154_, _23153_, _23151_);
  or (_23155_, _23154_, _06286_);
  and (_23156_, _07916_, \oc8051_golden_model_1.ACC [1]);
  or (_23157_, _23156_, _23143_);
  and (_23158_, _23157_, _07143_);
  nor (_23159_, _07143_, _23141_);
  or (_23161_, _23159_, _06285_);
  or (_23162_, _23161_, _23158_);
  and (_23163_, _23162_, _06282_);
  and (_23164_, _23163_, _23155_);
  nor (_23165_, _08600_, _23141_);
  and (_23166_, _14508_, _08600_);
  or (_23167_, _23166_, _23165_);
  and (_23168_, _23167_, _06281_);
  or (_23169_, _23168_, _06354_);
  or (_23170_, _23169_, _23164_);
  and (_23172_, _23170_, _23150_);
  or (_23173_, _23172_, _06345_);
  or (_23174_, _23157_, _06346_);
  and (_23175_, _23174_, _06278_);
  and (_23176_, _23175_, _23173_);
  and (_23177_, _14511_, _08600_);
  or (_23178_, _23177_, _23165_);
  and (_23179_, _23178_, _06277_);
  or (_23180_, _23179_, _06270_);
  or (_23181_, _23180_, _23176_);
  and (_23183_, _23166_, _14507_);
  or (_23184_, _23165_, _06271_);
  or (_23185_, _23184_, _23183_);
  and (_23186_, _23185_, _06267_);
  and (_23187_, _23186_, _23181_);
  or (_23188_, _23165_, _14551_);
  and (_23189_, _23188_, _06266_);
  and (_23190_, _23189_, _23167_);
  or (_23191_, _23190_, _06259_);
  or (_23192_, _23191_, _23187_);
  or (_23194_, _23148_, _06260_);
  and (_23195_, _23194_, _23192_);
  or (_23196_, _23195_, _09486_);
  and (_23197_, _09339_, _07916_);
  or (_23198_, _23143_, _06258_);
  or (_23199_, _23198_, _23197_);
  and (_23200_, _23199_, _06251_);
  and (_23201_, _23200_, _23196_);
  and (_23202_, _14607_, _07916_);
  or (_23203_, _23202_, _23143_);
  and (_23205_, _23203_, _05972_);
  or (_23206_, _23205_, _23201_);
  and (_23207_, _23206_, _06399_);
  or (_23208_, _14505_, _11860_);
  and (_23209_, _23208_, _06398_);
  nand (_23210_, _07916_, _07031_);
  and (_23211_, _23210_, _06215_);
  or (_23212_, _23211_, _23209_);
  and (_23213_, _23212_, _23151_);
  or (_23214_, _23213_, _06524_);
  or (_23216_, _23214_, _23207_);
  nand (_23217_, _11251_, _07916_);
  and (_23218_, _23217_, _23145_);
  or (_23219_, _23218_, _09030_);
  and (_23220_, _23219_, _07219_);
  and (_23221_, _23220_, _23216_);
  or (_23222_, _14503_, _11860_);
  and (_23223_, _23151_, _06426_);
  and (_23224_, _23223_, _23222_);
  or (_23225_, _23224_, _06532_);
  or (_23227_, _23225_, _23221_);
  nor (_23228_, _23143_, _07217_);
  nand (_23229_, _23228_, _23217_);
  and (_23230_, _23229_, _07229_);
  and (_23231_, _23230_, _23227_);
  or (_23232_, _23210_, _08325_);
  and (_23233_, _23151_, _06437_);
  and (_23234_, _23233_, _23232_);
  or (_23235_, _23234_, _06535_);
  or (_23236_, _23235_, _23231_);
  and (_23238_, _23236_, _23146_);
  or (_23239_, _23238_, _06559_);
  or (_23240_, _23154_, _07240_);
  and (_23241_, _23240_, _05933_);
  and (_23242_, _23241_, _23239_);
  and (_23243_, _23178_, _05932_);
  or (_23244_, _23243_, _06566_);
  or (_23245_, _23244_, _23242_);
  or (_23246_, _23143_, _06570_);
  or (_23247_, _23246_, _23152_);
  and (_23249_, _23247_, _01320_);
  and (_23250_, _23249_, _23245_);
  or (_23251_, _23250_, _23142_);
  and (_42958_, _23251_, _42355_);
  and (_23252_, _01324_, \oc8051_golden_model_1.TCON [2]);
  and (_23253_, _11860_, \oc8051_golden_model_1.TCON [2]);
  and (_23254_, _07916_, _08662_);
  or (_23255_, _23254_, _23253_);
  or (_23256_, _23255_, _06260_);
  and (_23257_, _23255_, _06354_);
  and (_23259_, _11865_, \oc8051_golden_model_1.TCON [2]);
  and (_23260_, _14716_, _08600_);
  or (_23261_, _23260_, _23259_);
  or (_23262_, _23261_, _06282_);
  and (_23263_, _14703_, _07916_);
  or (_23264_, _23263_, _23253_);
  and (_23265_, _23264_, _06285_);
  and (_23266_, _07144_, \oc8051_golden_model_1.TCON [2]);
  and (_23267_, _07916_, \oc8051_golden_model_1.ACC [2]);
  or (_23268_, _23267_, _23253_);
  and (_23270_, _23268_, _07143_);
  or (_23271_, _23270_, _23266_);
  and (_23272_, _23271_, _06286_);
  or (_23273_, _23272_, _06281_);
  or (_23274_, _23273_, _23265_);
  and (_23275_, _23274_, _23262_);
  and (_23276_, _23275_, _07169_);
  or (_23277_, _23276_, _23257_);
  or (_23278_, _23277_, _06345_);
  or (_23279_, _23268_, _06346_);
  and (_23281_, _23279_, _06278_);
  and (_23282_, _23281_, _23278_);
  and (_23283_, _14699_, _08600_);
  or (_23284_, _23283_, _23259_);
  and (_23285_, _23284_, _06277_);
  or (_23286_, _23285_, _06270_);
  or (_23287_, _23286_, _23282_);
  or (_23288_, _23259_, _14731_);
  and (_23289_, _23288_, _23261_);
  or (_23290_, _23289_, _06271_);
  and (_23292_, _23290_, _06267_);
  and (_23293_, _23292_, _23287_);
  and (_23294_, _14749_, _08600_);
  or (_23295_, _23294_, _23259_);
  and (_23296_, _23295_, _06266_);
  or (_23297_, _23296_, _06259_);
  or (_23298_, _23297_, _23293_);
  and (_23299_, _23298_, _23256_);
  or (_23300_, _23299_, _09486_);
  and (_23301_, _09293_, _07916_);
  or (_23303_, _23253_, _06258_);
  or (_23304_, _23303_, _23301_);
  and (_23305_, _23304_, _06251_);
  and (_23306_, _23305_, _23300_);
  and (_23307_, _14804_, _07916_);
  or (_23308_, _23253_, _23307_);
  and (_23309_, _23308_, _05972_);
  or (_23310_, _23309_, _23306_);
  or (_23311_, _23310_, _10080_);
  and (_23312_, _14697_, _07916_);
  or (_23314_, _23253_, _09025_);
  or (_23315_, _23314_, _23312_);
  and (_23316_, _07916_, _08980_);
  or (_23317_, _23316_, _23253_);
  or (_23318_, _23317_, _06216_);
  and (_23319_, _23318_, _09030_);
  and (_23320_, _23319_, _23315_);
  and (_23321_, _23320_, _23311_);
  and (_23322_, _11250_, _07916_);
  or (_23323_, _23322_, _23253_);
  and (_23325_, _23323_, _06524_);
  or (_23326_, _23325_, _23321_);
  and (_23327_, _23326_, _07219_);
  or (_23328_, _23253_, _08424_);
  and (_23329_, _23317_, _06426_);
  and (_23330_, _23329_, _23328_);
  or (_23331_, _23330_, _23327_);
  and (_23332_, _23331_, _07217_);
  and (_23333_, _23268_, _06532_);
  and (_23334_, _23333_, _23328_);
  or (_23336_, _23334_, _06437_);
  or (_23337_, _23336_, _23332_);
  and (_23338_, _14694_, _07916_);
  or (_23339_, _23253_, _07229_);
  or (_23340_, _23339_, _23338_);
  and (_23341_, _23340_, _07231_);
  and (_23342_, _23341_, _23337_);
  nor (_23343_, _11249_, _11860_);
  or (_23344_, _23343_, _23253_);
  and (_23345_, _23344_, _06535_);
  or (_23347_, _23345_, _06559_);
  or (_23348_, _23347_, _23342_);
  or (_23349_, _23264_, _07240_);
  and (_23350_, _23349_, _05933_);
  and (_23351_, _23350_, _23348_);
  and (_23352_, _23284_, _05932_);
  or (_23353_, _23352_, _06566_);
  or (_23354_, _23353_, _23351_);
  and (_23355_, _14873_, _07916_);
  or (_23356_, _23253_, _06570_);
  or (_23358_, _23356_, _23355_);
  and (_23359_, _23358_, _01320_);
  and (_23360_, _23359_, _23354_);
  or (_23361_, _23360_, _23252_);
  and (_42959_, _23361_, _42355_);
  and (_23362_, _01324_, \oc8051_golden_model_1.TCON [3]);
  and (_23363_, _11860_, \oc8051_golden_model_1.TCON [3]);
  and (_23364_, _07916_, _09421_);
  or (_23365_, _23364_, _23363_);
  or (_23366_, _23365_, _06260_);
  and (_23368_, _14900_, _07916_);
  or (_23369_, _23368_, _23363_);
  or (_23370_, _23369_, _06286_);
  and (_23371_, _07916_, \oc8051_golden_model_1.ACC [3]);
  or (_23372_, _23371_, _23363_);
  and (_23373_, _23372_, _07143_);
  and (_23374_, _07144_, \oc8051_golden_model_1.TCON [3]);
  or (_23375_, _23374_, _06285_);
  or (_23376_, _23375_, _23373_);
  and (_23377_, _23376_, _06282_);
  and (_23378_, _23377_, _23370_);
  and (_23379_, _11865_, \oc8051_golden_model_1.TCON [3]);
  and (_23380_, _14897_, _08600_);
  or (_23381_, _23380_, _23379_);
  and (_23382_, _23381_, _06281_);
  or (_23383_, _23382_, _06354_);
  or (_23384_, _23383_, _23378_);
  or (_23385_, _23365_, _07169_);
  and (_23386_, _23385_, _23384_);
  or (_23387_, _23386_, _06345_);
  or (_23390_, _23372_, _06346_);
  and (_23391_, _23390_, _06278_);
  and (_23392_, _23391_, _23387_);
  and (_23393_, _14895_, _08600_);
  or (_23394_, _23393_, _23379_);
  and (_23395_, _23394_, _06277_);
  or (_23396_, _23395_, _06270_);
  or (_23397_, _23396_, _23392_);
  or (_23398_, _23379_, _14926_);
  and (_23399_, _23398_, _23381_);
  or (_23401_, _23399_, _06271_);
  and (_23402_, _23401_, _06267_);
  and (_23403_, _23402_, _23397_);
  and (_23404_, _14943_, _08600_);
  or (_23405_, _23404_, _23379_);
  and (_23406_, _23405_, _06266_);
  or (_23407_, _23406_, _06259_);
  or (_23408_, _23407_, _23403_);
  and (_23409_, _23408_, _23366_);
  or (_23410_, _23409_, _09486_);
  and (_23412_, _09247_, _07916_);
  or (_23413_, _23363_, _06258_);
  or (_23414_, _23413_, _23412_);
  and (_23415_, _23414_, _06251_);
  and (_23416_, _23415_, _23410_);
  and (_23417_, _14998_, _07916_);
  or (_23418_, _23363_, _23417_);
  and (_23419_, _23418_, _05972_);
  or (_23420_, _23419_, _23416_);
  or (_23421_, _23420_, _10080_);
  and (_23423_, _14893_, _07916_);
  or (_23424_, _23363_, _09025_);
  or (_23425_, _23424_, _23423_);
  and (_23426_, _07916_, _08809_);
  or (_23427_, _23426_, _23363_);
  or (_23428_, _23427_, _06216_);
  and (_23429_, _23428_, _09030_);
  and (_23430_, _23429_, _23425_);
  and (_23431_, _23430_, _23421_);
  and (_23432_, _12529_, _07916_);
  or (_23434_, _23432_, _23363_);
  and (_23435_, _23434_, _06524_);
  or (_23436_, _23435_, _23431_);
  and (_23437_, _23436_, _07219_);
  or (_23438_, _23363_, _08280_);
  and (_23439_, _23427_, _06426_);
  and (_23440_, _23439_, _23438_);
  or (_23441_, _23440_, _23437_);
  and (_23442_, _23441_, _07217_);
  and (_23443_, _23372_, _06532_);
  and (_23445_, _23443_, _23438_);
  or (_23446_, _23445_, _06437_);
  or (_23447_, _23446_, _23442_);
  and (_23448_, _14890_, _07916_);
  or (_23449_, _23363_, _07229_);
  or (_23450_, _23449_, _23448_);
  and (_23451_, _23450_, _07231_);
  and (_23452_, _23451_, _23447_);
  nor (_23453_, _11247_, _11860_);
  or (_23454_, _23453_, _23363_);
  and (_23456_, _23454_, _06535_);
  or (_23457_, _23456_, _06559_);
  or (_23458_, _23457_, _23452_);
  or (_23459_, _23369_, _07240_);
  and (_23460_, _23459_, _05933_);
  and (_23461_, _23460_, _23458_);
  and (_23462_, _23394_, _05932_);
  or (_23463_, _23462_, _06566_);
  or (_23464_, _23463_, _23461_);
  and (_23465_, _15068_, _07916_);
  or (_23467_, _23363_, _06570_);
  or (_23468_, _23467_, _23465_);
  and (_23469_, _23468_, _01320_);
  and (_23470_, _23469_, _23464_);
  or (_23471_, _23470_, _23362_);
  and (_42961_, _23471_, _42355_);
  and (_23472_, _01324_, \oc8051_golden_model_1.TCON [4]);
  and (_23473_, _11860_, \oc8051_golden_model_1.TCON [4]);
  and (_23474_, _09420_, _07916_);
  or (_23475_, _23474_, _23473_);
  or (_23477_, _23475_, _06260_);
  and (_23478_, _11865_, \oc8051_golden_model_1.TCON [4]);
  and (_23479_, _15145_, _08600_);
  or (_23480_, _23479_, _23478_);
  and (_23481_, _23480_, _06277_);
  and (_23482_, _15133_, _07916_);
  or (_23483_, _23482_, _23473_);
  or (_23484_, _23483_, _06286_);
  and (_23485_, _07916_, \oc8051_golden_model_1.ACC [4]);
  or (_23486_, _23485_, _23473_);
  and (_23488_, _23486_, _07143_);
  and (_23489_, _07144_, \oc8051_golden_model_1.TCON [4]);
  or (_23490_, _23489_, _06285_);
  or (_23491_, _23490_, _23488_);
  and (_23492_, _23491_, _06282_);
  and (_23493_, _23492_, _23484_);
  and (_23494_, _15116_, _08600_);
  or (_23495_, _23494_, _23478_);
  and (_23496_, _23495_, _06281_);
  or (_23497_, _23496_, _06354_);
  or (_23499_, _23497_, _23493_);
  or (_23500_, _23475_, _07169_);
  and (_23501_, _23500_, _23499_);
  or (_23502_, _23501_, _06345_);
  or (_23503_, _23486_, _06346_);
  and (_23504_, _23503_, _06278_);
  and (_23505_, _23504_, _23502_);
  or (_23506_, _23505_, _23481_);
  and (_23507_, _23506_, _06271_);
  or (_23508_, _23478_, _15152_);
  and (_23510_, _23508_, _06270_);
  and (_23511_, _23510_, _23495_);
  or (_23512_, _23511_, _23507_);
  and (_23513_, _23512_, _06267_);
  and (_23514_, _15170_, _08600_);
  or (_23515_, _23514_, _23478_);
  and (_23516_, _23515_, _06266_);
  or (_23517_, _23516_, _06259_);
  or (_23518_, _23517_, _23513_);
  and (_23519_, _23518_, _23477_);
  or (_23521_, _23519_, _09486_);
  and (_23522_, _09437_, _07916_);
  or (_23523_, _23473_, _06258_);
  or (_23524_, _23523_, _23522_);
  and (_23525_, _23524_, _06251_);
  and (_23526_, _23525_, _23521_);
  and (_23527_, _15226_, _07916_);
  or (_23528_, _23527_, _23473_);
  and (_23529_, _23528_, _05972_);
  or (_23530_, _23529_, _10080_);
  or (_23532_, _23530_, _23526_);
  and (_23533_, _15114_, _07916_);
  or (_23534_, _23473_, _09025_);
  or (_23535_, _23534_, _23533_);
  and (_23536_, _08919_, _07916_);
  or (_23537_, _23536_, _23473_);
  or (_23538_, _23537_, _06216_);
  and (_23539_, _23538_, _09030_);
  and (_23540_, _23539_, _23535_);
  and (_23541_, _23540_, _23532_);
  and (_23543_, _11245_, _07916_);
  or (_23544_, _23543_, _23473_);
  and (_23545_, _23544_, _06524_);
  or (_23546_, _23545_, _23541_);
  and (_23547_, _23546_, _07219_);
  or (_23548_, _23473_, _08528_);
  and (_23549_, _23537_, _06426_);
  and (_23550_, _23549_, _23548_);
  or (_23551_, _23550_, _23547_);
  and (_23552_, _23551_, _07217_);
  and (_23554_, _23486_, _06532_);
  and (_23555_, _23554_, _23548_);
  or (_23556_, _23555_, _06437_);
  or (_23557_, _23556_, _23552_);
  and (_23558_, _15111_, _07916_);
  or (_23559_, _23473_, _07229_);
  or (_23560_, _23559_, _23558_);
  and (_23561_, _23560_, _07231_);
  and (_23562_, _23561_, _23557_);
  nor (_23563_, _11244_, _11860_);
  or (_23565_, _23563_, _23473_);
  and (_23566_, _23565_, _06535_);
  or (_23567_, _23566_, _06559_);
  or (_23568_, _23567_, _23562_);
  or (_23569_, _23483_, _07240_);
  and (_23570_, _23569_, _05933_);
  and (_23571_, _23570_, _23568_);
  and (_23572_, _23480_, _05932_);
  or (_23573_, _23572_, _06566_);
  or (_23574_, _23573_, _23571_);
  and (_23576_, _15296_, _07916_);
  or (_23577_, _23473_, _06570_);
  or (_23578_, _23577_, _23576_);
  and (_23579_, _23578_, _01320_);
  and (_23580_, _23579_, _23574_);
  or (_23581_, _23580_, _23472_);
  and (_42962_, _23581_, _42355_);
  and (_23582_, _01324_, \oc8051_golden_model_1.TCON [5]);
  and (_23583_, _11860_, \oc8051_golden_model_1.TCON [5]);
  and (_23584_, _15330_, _07916_);
  or (_23586_, _23584_, _23583_);
  or (_23587_, _23586_, _06286_);
  and (_23588_, _07916_, \oc8051_golden_model_1.ACC [5]);
  or (_23589_, _23588_, _23583_);
  and (_23590_, _23589_, _07143_);
  and (_23591_, _07144_, \oc8051_golden_model_1.TCON [5]);
  or (_23592_, _23591_, _06285_);
  or (_23593_, _23592_, _23590_);
  and (_23594_, _23593_, _06282_);
  and (_23595_, _23594_, _23587_);
  and (_23597_, _11865_, \oc8051_golden_model_1.TCON [5]);
  and (_23598_, _15315_, _08600_);
  or (_23599_, _23598_, _23597_);
  and (_23600_, _23599_, _06281_);
  or (_23601_, _23600_, _06354_);
  or (_23602_, _23601_, _23595_);
  and (_23603_, _09419_, _07916_);
  or (_23604_, _23603_, _23583_);
  or (_23605_, _23604_, _07169_);
  and (_23606_, _23605_, _23602_);
  or (_23608_, _23606_, _06345_);
  or (_23609_, _23589_, _06346_);
  and (_23610_, _23609_, _06278_);
  and (_23611_, _23610_, _23608_);
  and (_23612_, _15342_, _08600_);
  or (_23613_, _23612_, _23597_);
  and (_23614_, _23613_, _06277_);
  or (_23615_, _23614_, _06270_);
  or (_23616_, _23615_, _23611_);
  or (_23617_, _23597_, _15349_);
  and (_23619_, _23617_, _23599_);
  or (_23620_, _23619_, _06271_);
  and (_23621_, _23620_, _06267_);
  and (_23622_, _23621_, _23616_);
  or (_23623_, _23597_, _15365_);
  and (_23624_, _23623_, _06266_);
  and (_23625_, _23624_, _23599_);
  or (_23626_, _23625_, _06259_);
  or (_23627_, _23626_, _23622_);
  or (_23628_, _23604_, _06260_);
  and (_23629_, _23628_, _23627_);
  or (_23630_, _23629_, _09486_);
  and (_23631_, _09436_, _07916_);
  or (_23632_, _23583_, _06258_);
  or (_23633_, _23632_, _23631_);
  and (_23634_, _23633_, _06251_);
  and (_23635_, _23634_, _23630_);
  and (_23636_, _15421_, _07916_);
  or (_23637_, _23636_, _23583_);
  and (_23638_, _23637_, _05972_);
  or (_23640_, _23638_, _10080_);
  or (_23641_, _23640_, _23635_);
  and (_23642_, _15313_, _07916_);
  or (_23643_, _23583_, _09025_);
  or (_23644_, _23643_, _23642_);
  and (_23645_, _08913_, _07916_);
  or (_23646_, _23645_, _23583_);
  or (_23647_, _23646_, _06216_);
  and (_23648_, _23647_, _09030_);
  and (_23649_, _23648_, _23644_);
  and (_23651_, _23649_, _23641_);
  and (_23652_, _12536_, _07916_);
  or (_23653_, _23652_, _23583_);
  and (_23654_, _23653_, _06524_);
  or (_23655_, _23654_, _23651_);
  and (_23656_, _23655_, _07219_);
  or (_23657_, _23583_, _08231_);
  and (_23658_, _23646_, _06426_);
  and (_23659_, _23658_, _23657_);
  or (_23660_, _23659_, _23656_);
  and (_23662_, _23660_, _07217_);
  and (_23663_, _23589_, _06532_);
  and (_23664_, _23663_, _23657_);
  or (_23665_, _23664_, _06437_);
  or (_23666_, _23665_, _23662_);
  and (_23667_, _15310_, _07916_);
  or (_23668_, _23583_, _07229_);
  or (_23669_, _23668_, _23667_);
  and (_23670_, _23669_, _07231_);
  and (_23671_, _23670_, _23666_);
  nor (_23672_, _11241_, _11860_);
  or (_23673_, _23672_, _23583_);
  and (_23674_, _23673_, _06535_);
  or (_23675_, _23674_, _06559_);
  or (_23676_, _23675_, _23671_);
  or (_23677_, _23586_, _07240_);
  and (_23678_, _23677_, _05933_);
  and (_23679_, _23678_, _23676_);
  and (_23680_, _23613_, _05932_);
  or (_23681_, _23680_, _06566_);
  or (_23683_, _23681_, _23679_);
  and (_23684_, _15493_, _07916_);
  or (_23685_, _23583_, _06570_);
  or (_23686_, _23685_, _23684_);
  and (_23687_, _23686_, _01320_);
  and (_23688_, _23687_, _23683_);
  or (_23689_, _23688_, _23582_);
  and (_42963_, _23689_, _42355_);
  and (_23690_, _01324_, \oc8051_golden_model_1.TCON [6]);
  and (_23691_, _11860_, \oc8051_golden_model_1.TCON [6]);
  and (_23692_, _15521_, _07916_);
  or (_23693_, _23692_, _23691_);
  or (_23694_, _23693_, _06286_);
  and (_23695_, _07916_, \oc8051_golden_model_1.ACC [6]);
  or (_23696_, _23695_, _23691_);
  and (_23697_, _23696_, _07143_);
  and (_23698_, _07144_, \oc8051_golden_model_1.TCON [6]);
  or (_23699_, _23698_, _06285_);
  or (_23700_, _23699_, _23697_);
  and (_23701_, _23700_, _06282_);
  and (_23703_, _23701_, _23694_);
  and (_23704_, _11865_, \oc8051_golden_model_1.TCON [6]);
  and (_23705_, _15535_, _08600_);
  or (_23706_, _23705_, _23704_);
  and (_23707_, _23706_, _06281_);
  or (_23708_, _23707_, _06354_);
  or (_23709_, _23708_, _23703_);
  and (_23710_, _09418_, _07916_);
  or (_23711_, _23710_, _23691_);
  or (_23712_, _23711_, _07169_);
  and (_23714_, _23712_, _23709_);
  or (_23715_, _23714_, _06345_);
  or (_23716_, _23696_, _06346_);
  and (_23717_, _23716_, _06278_);
  and (_23718_, _23717_, _23715_);
  and (_23719_, _15544_, _08600_);
  or (_23720_, _23719_, _23704_);
  and (_23721_, _23720_, _06277_);
  or (_23722_, _23721_, _06270_);
  or (_23723_, _23722_, _23718_);
  or (_23724_, _23704_, _15551_);
  and (_23725_, _23724_, _23706_);
  or (_23726_, _23725_, _06271_);
  and (_23727_, _23726_, _06267_);
  and (_23728_, _23727_, _23723_);
  and (_23729_, _15568_, _08600_);
  or (_23730_, _23729_, _23704_);
  and (_23731_, _23730_, _06266_);
  or (_23732_, _23731_, _06259_);
  or (_23733_, _23732_, _23728_);
  or (_23735_, _23711_, _06260_);
  and (_23736_, _23735_, _23733_);
  or (_23737_, _23736_, _09486_);
  and (_23738_, _09435_, _07916_);
  or (_23739_, _23691_, _06258_);
  or (_23740_, _23739_, _23738_);
  and (_23741_, _23740_, _06251_);
  and (_23742_, _23741_, _23737_);
  and (_23743_, _15623_, _07916_);
  or (_23744_, _23743_, _23691_);
  and (_23746_, _23744_, _05972_);
  or (_23747_, _23746_, _10080_);
  or (_23748_, _23747_, _23742_);
  and (_23749_, _15517_, _07916_);
  or (_23750_, _23691_, _09025_);
  or (_23751_, _23750_, _23749_);
  and (_23752_, _08845_, _07916_);
  or (_23753_, _23752_, _23691_);
  or (_23754_, _23753_, _06216_);
  and (_23755_, _23754_, _09030_);
  and (_23756_, _23755_, _23751_);
  and (_23757_, _23756_, _23748_);
  and (_23758_, _11239_, _07916_);
  or (_23759_, _23758_, _23691_);
  and (_23760_, _23759_, _06524_);
  or (_23761_, _23760_, _23757_);
  and (_23762_, _23761_, _07219_);
  or (_23763_, _23691_, _08128_);
  and (_23764_, _23753_, _06426_);
  and (_23765_, _23764_, _23763_);
  or (_23767_, _23765_, _23762_);
  and (_23768_, _23767_, _07217_);
  and (_23769_, _23696_, _06532_);
  and (_23770_, _23769_, _23763_);
  or (_23771_, _23770_, _06437_);
  or (_23772_, _23771_, _23768_);
  and (_23773_, _15514_, _07916_);
  or (_23774_, _23691_, _07229_);
  or (_23775_, _23774_, _23773_);
  and (_23776_, _23775_, _07231_);
  and (_23778_, _23776_, _23772_);
  nor (_23779_, _11238_, _11860_);
  or (_23780_, _23779_, _23691_);
  and (_23781_, _23780_, _06535_);
  or (_23782_, _23781_, _06559_);
  or (_23783_, _23782_, _23778_);
  or (_23784_, _23693_, _07240_);
  and (_23785_, _23784_, _05933_);
  and (_23786_, _23785_, _23783_);
  and (_23787_, _23720_, _05932_);
  or (_23788_, _23787_, _06566_);
  or (_23789_, _23788_, _23786_);
  and (_23790_, _15695_, _07916_);
  or (_23791_, _23691_, _06570_);
  or (_23792_, _23791_, _23790_);
  and (_23793_, _23792_, _01320_);
  and (_23794_, _23793_, _23789_);
  or (_23795_, _23794_, _23690_);
  and (_42964_, _23795_, _42355_);
  and (_23796_, _01324_, \oc8051_golden_model_1.TH1 [0]);
  and (_23798_, _07900_, \oc8051_golden_model_1.ACC [0]);
  and (_23799_, _23798_, _08374_);
  and (_23800_, _11961_, \oc8051_golden_model_1.TH1 [0]);
  or (_23801_, _23800_, _07217_);
  or (_23802_, _23801_, _23799_);
  or (_23803_, _23800_, _23798_);
  and (_23804_, _23803_, _06345_);
  or (_23805_, _23804_, _06259_);
  nor (_23806_, _08374_, _11961_);
  or (_23807_, _23806_, _23800_);
  and (_23808_, _23807_, _06285_);
  and (_23809_, _07144_, \oc8051_golden_model_1.TH1 [0]);
  and (_23810_, _23803_, _07143_);
  or (_23811_, _23810_, _23809_);
  and (_23812_, _23811_, _06286_);
  or (_23813_, _23812_, _06354_);
  or (_23814_, _23813_, _23808_);
  and (_23815_, _23814_, _06346_);
  or (_23816_, _23815_, _23805_);
  and (_23817_, _07900_, _07135_);
  or (_23819_, _23800_, _19434_);
  or (_23820_, _23819_, _23817_);
  and (_23821_, _23820_, _23816_);
  or (_23822_, _23821_, _09486_);
  and (_23823_, _09384_, _07900_);
  or (_23824_, _23800_, _06258_);
  or (_23825_, _23824_, _23823_);
  and (_23826_, _23825_, _23822_);
  or (_23827_, _23826_, _05972_);
  and (_23828_, _14413_, _07900_);
  or (_23830_, _23800_, _06251_);
  or (_23831_, _23830_, _23828_);
  and (_23832_, _23831_, _06216_);
  and (_23833_, _23832_, _23827_);
  and (_23834_, _07900_, _08929_);
  or (_23835_, _23834_, _23800_);
  and (_23836_, _23835_, _06215_);
  or (_23837_, _23836_, _06398_);
  or (_23838_, _23837_, _23833_);
  and (_23839_, _14311_, _07900_);
  or (_23841_, _23839_, _23800_);
  or (_23842_, _23841_, _09025_);
  and (_23843_, _23842_, _09030_);
  and (_23844_, _23843_, _23838_);
  nor (_23845_, _12532_, _11961_);
  or (_23846_, _23845_, _23800_);
  nor (_23847_, _23799_, _09030_);
  and (_23848_, _23847_, _23846_);
  or (_23849_, _23848_, _23844_);
  and (_23850_, _23849_, _07219_);
  nand (_23851_, _23835_, _06426_);
  nor (_23852_, _23851_, _23806_);
  or (_23853_, _23852_, _06532_);
  or (_23854_, _23853_, _23850_);
  and (_23855_, _23854_, _23802_);
  or (_23856_, _23855_, _06437_);
  and (_23857_, _14307_, _07900_);
  or (_23858_, _23800_, _07229_);
  or (_23859_, _23858_, _23857_);
  and (_23860_, _23859_, _07231_);
  and (_23862_, _23860_, _23856_);
  and (_23863_, _23846_, _06535_);
  or (_23864_, _23863_, _19480_);
  or (_23865_, _23864_, _23862_);
  or (_23866_, _23807_, _06651_);
  and (_23867_, _23866_, _01320_);
  and (_23868_, _23867_, _23865_);
  or (_23869_, _23868_, _23796_);
  and (_42966_, _23869_, _42355_);
  and (_23870_, _01324_, \oc8051_golden_model_1.TH1 [1]);
  and (_23872_, _11961_, \oc8051_golden_model_1.TH1 [1]);
  and (_23873_, _07900_, _09422_);
  or (_23874_, _23873_, _23872_);
  or (_23875_, _23874_, _06260_);
  and (_23876_, _07900_, \oc8051_golden_model_1.ACC [1]);
  or (_23877_, _23876_, _23872_);
  and (_23878_, _23877_, _06345_);
  or (_23879_, _23878_, _06259_);
  or (_23880_, _07900_, \oc8051_golden_model_1.TH1 [1]);
  and (_23881_, _14520_, _07900_);
  not (_23882_, _23881_);
  and (_23883_, _23882_, _23880_);
  and (_23884_, _23883_, _06285_);
  and (_23885_, _07144_, \oc8051_golden_model_1.TH1 [1]);
  and (_23886_, _23877_, _07143_);
  or (_23887_, _23886_, _23885_);
  and (_23888_, _23887_, _06286_);
  or (_23889_, _23888_, _06354_);
  or (_23890_, _23889_, _23884_);
  or (_23891_, _23874_, _07169_);
  and (_23893_, _23891_, _06346_);
  and (_23894_, _23893_, _23890_);
  or (_23895_, _23894_, _23879_);
  and (_23896_, _23895_, _23875_);
  or (_23897_, _23896_, _09486_);
  and (_23898_, _23897_, _06251_);
  and (_23899_, _09339_, _07900_);
  or (_23900_, _23872_, _06258_);
  or (_23901_, _23900_, _23899_);
  and (_23902_, _23901_, _23898_);
  or (_23904_, _14607_, _11961_);
  and (_23905_, _23880_, _05972_);
  and (_23906_, _23905_, _23904_);
  or (_23907_, _23906_, _23902_);
  and (_23908_, _23907_, _06399_);
  or (_23909_, _14505_, _11961_);
  and (_23910_, _23909_, _06398_);
  nand (_23911_, _07900_, _07031_);
  and (_23912_, _23911_, _06215_);
  or (_23913_, _23912_, _23910_);
  and (_23914_, _23913_, _23880_);
  or (_23915_, _23914_, _06524_);
  or (_23916_, _23915_, _23908_);
  and (_23917_, _11253_, _07900_);
  or (_23918_, _23917_, _23872_);
  or (_23919_, _23918_, _09030_);
  and (_23920_, _23919_, _07219_);
  and (_23921_, _23920_, _23916_);
  or (_23922_, _14503_, _11961_);
  and (_23923_, _23880_, _06426_);
  and (_23925_, _23923_, _23922_);
  or (_23926_, _23925_, _06532_);
  or (_23927_, _23926_, _23921_);
  and (_23928_, _23876_, _08325_);
  or (_23929_, _23872_, _07217_);
  or (_23930_, _23929_, _23928_);
  and (_23931_, _23930_, _07229_);
  and (_23932_, _23931_, _23927_);
  or (_23933_, _23911_, _08325_);
  and (_23934_, _23880_, _06437_);
  and (_23936_, _23934_, _23933_);
  or (_23937_, _23936_, _06535_);
  or (_23938_, _23937_, _23932_);
  nor (_23939_, _11252_, _11961_);
  or (_23940_, _23939_, _23872_);
  or (_23941_, _23940_, _07231_);
  and (_23942_, _23941_, _07240_);
  and (_23943_, _23942_, _23938_);
  and (_23944_, _23883_, _06559_);
  or (_23945_, _23944_, _06566_);
  or (_23946_, _23945_, _23943_);
  or (_23947_, _23872_, _06570_);
  or (_23948_, _23947_, _23881_);
  and (_23949_, _23948_, _01320_);
  and (_23950_, _23949_, _23946_);
  or (_23951_, _23950_, _23870_);
  and (_42967_, _23951_, _42355_);
  and (_23952_, _01324_, \oc8051_golden_model_1.TH1 [2]);
  and (_23953_, _11961_, \oc8051_golden_model_1.TH1 [2]);
  and (_23954_, _07900_, _08662_);
  or (_23956_, _23954_, _23953_);
  or (_23957_, _23956_, _06260_);
  and (_23958_, _14703_, _07900_);
  or (_23959_, _23958_, _23953_);
  and (_23960_, _23959_, _06285_);
  and (_23961_, _07144_, \oc8051_golden_model_1.TH1 [2]);
  and (_23962_, _07900_, \oc8051_golden_model_1.ACC [2]);
  or (_23963_, _23962_, _23953_);
  and (_23964_, _23963_, _07143_);
  or (_23965_, _23964_, _23961_);
  and (_23967_, _23965_, _06286_);
  or (_23968_, _23967_, _06354_);
  or (_23969_, _23968_, _23960_);
  or (_23970_, _23956_, _07169_);
  and (_23971_, _23970_, _06346_);
  and (_23972_, _23971_, _23969_);
  and (_23973_, _23963_, _06345_);
  or (_23974_, _23973_, _06259_);
  or (_23975_, _23974_, _23972_);
  and (_23976_, _23975_, _23957_);
  or (_23977_, _23976_, _09486_);
  and (_23978_, _09293_, _07900_);
  or (_23979_, _23953_, _06258_);
  or (_23980_, _23979_, _23978_);
  and (_23981_, _23980_, _23977_);
  or (_23982_, _23981_, _05972_);
  and (_23983_, _14804_, _07900_);
  or (_23984_, _23953_, _06251_);
  or (_23985_, _23984_, _23983_);
  and (_23986_, _23985_, _06216_);
  and (_23987_, _23986_, _23982_);
  nor (_23988_, _11961_, _06689_);
  or (_23989_, _23988_, _23953_);
  and (_23990_, _23989_, _06215_);
  or (_23991_, _23990_, _06398_);
  or (_23992_, _23991_, _23987_);
  and (_23993_, _14697_, _07900_);
  or (_23994_, _23993_, _23953_);
  or (_23995_, _23994_, _09025_);
  and (_23996_, _23995_, _09030_);
  and (_23999_, _23996_, _23992_);
  and (_24000_, _11250_, _07900_);
  or (_24001_, _24000_, _23953_);
  and (_24002_, _24001_, _06524_);
  or (_24003_, _24002_, _23999_);
  and (_24004_, _24003_, _07219_);
  or (_24005_, _23953_, _08424_);
  and (_24006_, _23989_, _06426_);
  and (_24007_, _24006_, _24005_);
  or (_24008_, _24007_, _24004_);
  and (_24009_, _24008_, _07217_);
  and (_24010_, _23963_, _06532_);
  and (_24011_, _24010_, _24005_);
  or (_24012_, _24011_, _06437_);
  or (_24013_, _24012_, _24009_);
  and (_24014_, _14694_, _07900_);
  or (_24015_, _23953_, _07229_);
  or (_24016_, _24015_, _24014_);
  and (_24017_, _24016_, _07231_);
  and (_24018_, _24017_, _24013_);
  nor (_24020_, _11249_, _11961_);
  or (_24021_, _24020_, _23953_);
  and (_24022_, _24021_, _06535_);
  or (_24023_, _24022_, _24018_);
  and (_24024_, _24023_, _07240_);
  and (_24025_, _23959_, _06559_);
  or (_24026_, _24025_, _06566_);
  or (_24027_, _24026_, _24024_);
  and (_24028_, _14873_, _07900_);
  or (_24029_, _23953_, _06570_);
  or (_24031_, _24029_, _24028_);
  and (_24032_, _24031_, _01320_);
  and (_24033_, _24032_, _24027_);
  or (_24034_, _24033_, _23952_);
  and (_42968_, _24034_, _42355_);
  and (_24035_, _11961_, \oc8051_golden_model_1.TH1 [3]);
  and (_24036_, _14900_, _07900_);
  or (_24037_, _24036_, _24035_);
  or (_24038_, _24037_, _06286_);
  and (_24039_, _07900_, \oc8051_golden_model_1.ACC [3]);
  or (_24041_, _24039_, _24035_);
  and (_24042_, _24041_, _07143_);
  and (_24043_, _07144_, \oc8051_golden_model_1.TH1 [3]);
  or (_24044_, _24043_, _06285_);
  or (_24045_, _24044_, _24042_);
  and (_24046_, _24045_, _07169_);
  and (_24047_, _24046_, _24038_);
  and (_24048_, _07900_, _09421_);
  or (_24049_, _24048_, _24035_);
  and (_24050_, _24049_, _06354_);
  or (_24051_, _24050_, _24047_);
  and (_24052_, _24051_, _06346_);
  and (_24053_, _24041_, _06345_);
  or (_24054_, _24053_, _06259_);
  or (_24055_, _24054_, _24052_);
  or (_24056_, _24049_, _06260_);
  and (_24057_, _24056_, _06258_);
  and (_24058_, _24057_, _24055_);
  and (_24059_, _09247_, _07900_);
  or (_24060_, _24059_, _24035_);
  and (_24062_, _24060_, _09486_);
  or (_24063_, _24062_, _05972_);
  or (_24064_, _24063_, _24058_);
  and (_24065_, _14998_, _07900_);
  or (_24066_, _24035_, _06251_);
  or (_24067_, _24066_, _24065_);
  and (_24068_, _24067_, _06216_);
  and (_24069_, _24068_, _24064_);
  nor (_24070_, _11961_, _06517_);
  or (_24071_, _24070_, _24035_);
  and (_24073_, _24071_, _06215_);
  or (_24074_, _24073_, _06398_);
  or (_24075_, _24074_, _24069_);
  and (_24076_, _14893_, _07900_);
  or (_24077_, _24076_, _24035_);
  or (_24078_, _24077_, _09025_);
  and (_24079_, _24078_, _09030_);
  and (_24080_, _24079_, _24075_);
  and (_24081_, _12529_, _07900_);
  or (_24082_, _24081_, _24035_);
  and (_24083_, _24082_, _06524_);
  or (_24084_, _24083_, _24080_);
  and (_24085_, _24084_, _07219_);
  or (_24086_, _24035_, _08280_);
  and (_24087_, _24071_, _06426_);
  and (_24088_, _24087_, _24086_);
  or (_24089_, _24088_, _24085_);
  and (_24090_, _24089_, _07217_);
  and (_24091_, _24041_, _06532_);
  and (_24092_, _24091_, _24086_);
  or (_24094_, _24092_, _06437_);
  or (_24095_, _24094_, _24090_);
  and (_24096_, _14890_, _07900_);
  or (_24097_, _24035_, _07229_);
  or (_24098_, _24097_, _24096_);
  and (_24099_, _24098_, _07231_);
  and (_24100_, _24099_, _24095_);
  nor (_24101_, _11247_, _11961_);
  or (_24102_, _24101_, _24035_);
  and (_24103_, _24102_, _06535_);
  or (_24105_, _24103_, _06559_);
  or (_24106_, _24105_, _24100_);
  or (_24107_, _24037_, _07240_);
  and (_24108_, _24107_, _06570_);
  and (_24109_, _24108_, _24106_);
  and (_24110_, _15068_, _07900_);
  or (_24111_, _24110_, _24035_);
  and (_24112_, _24111_, _06566_);
  or (_24113_, _24112_, _01324_);
  or (_24114_, _24113_, _24109_);
  or (_24116_, _01320_, \oc8051_golden_model_1.TH1 [3]);
  and (_24117_, _24116_, _42355_);
  and (_42969_, _24117_, _24114_);
  and (_24118_, _11961_, \oc8051_golden_model_1.TH1 [4]);
  and (_24119_, _15133_, _07900_);
  or (_24120_, _24119_, _24118_);
  or (_24121_, _24120_, _06286_);
  and (_24122_, _07900_, \oc8051_golden_model_1.ACC [4]);
  or (_24123_, _24122_, _24118_);
  and (_24124_, _24123_, _07143_);
  and (_24125_, _07144_, \oc8051_golden_model_1.TH1 [4]);
  or (_24126_, _24125_, _06285_);
  or (_24127_, _24126_, _24124_);
  and (_24128_, _24127_, _07169_);
  and (_24129_, _24128_, _24121_);
  and (_24130_, _09420_, _07900_);
  or (_24131_, _24130_, _24118_);
  and (_24132_, _24131_, _06354_);
  or (_24133_, _24132_, _24129_);
  and (_24134_, _24133_, _06346_);
  and (_24136_, _24123_, _06345_);
  or (_24137_, _24136_, _06259_);
  or (_24138_, _24137_, _24134_);
  or (_24139_, _24131_, _06260_);
  and (_24140_, _24139_, _24138_);
  or (_24141_, _24140_, _09486_);
  and (_24142_, _09437_, _07900_);
  or (_24143_, _24118_, _06258_);
  or (_24144_, _24143_, _24142_);
  and (_24145_, _24144_, _06251_);
  and (_24147_, _24145_, _24141_);
  and (_24148_, _15226_, _07900_);
  or (_24149_, _24148_, _24118_);
  and (_24150_, _24149_, _05972_);
  or (_24151_, _24150_, _24147_);
  or (_24152_, _24151_, _10080_);
  and (_24153_, _15114_, _07900_);
  or (_24154_, _24118_, _09025_);
  or (_24155_, _24154_, _24153_);
  nor (_24156_, _08879_, _11961_);
  or (_24157_, _24156_, _24118_);
  or (_24158_, _24157_, _06216_);
  and (_24159_, _24158_, _09030_);
  and (_24160_, _24159_, _24155_);
  and (_24161_, _24160_, _24152_);
  and (_24162_, _11245_, _07900_);
  or (_24163_, _24162_, _24118_);
  and (_24164_, _24163_, _06524_);
  or (_24165_, _24164_, _24161_);
  and (_24166_, _24165_, _07219_);
  or (_24168_, _24118_, _08528_);
  and (_24169_, _24157_, _06426_);
  and (_24170_, _24169_, _24168_);
  or (_24171_, _24170_, _24166_);
  and (_24172_, _24171_, _07217_);
  and (_24173_, _24123_, _06532_);
  and (_24174_, _24173_, _24168_);
  or (_24175_, _24174_, _06437_);
  or (_24176_, _24175_, _24172_);
  and (_24177_, _15111_, _07900_);
  or (_24179_, _24118_, _07229_);
  or (_24180_, _24179_, _24177_);
  and (_24181_, _24180_, _07231_);
  and (_24182_, _24181_, _24176_);
  nor (_24183_, _11244_, _11961_);
  or (_24184_, _24183_, _24118_);
  and (_24185_, _24184_, _06535_);
  or (_24186_, _24185_, _06559_);
  or (_24187_, _24186_, _24182_);
  or (_24188_, _24120_, _07240_);
  and (_24190_, _24188_, _06570_);
  and (_24191_, _24190_, _24187_);
  and (_24192_, _15296_, _07900_);
  or (_24193_, _24192_, _24118_);
  and (_24194_, _24193_, _06566_);
  or (_24195_, _24194_, _01324_);
  or (_24196_, _24195_, _24191_);
  or (_24197_, _01320_, \oc8051_golden_model_1.TH1 [4]);
  and (_24198_, _24197_, _42355_);
  and (_42970_, _24198_, _24196_);
  and (_24200_, _11961_, \oc8051_golden_model_1.TH1 [5]);
  and (_24201_, _15330_, _07900_);
  or (_24202_, _24201_, _24200_);
  or (_24203_, _24202_, _06286_);
  and (_24204_, _07900_, \oc8051_golden_model_1.ACC [5]);
  or (_24205_, _24204_, _24200_);
  and (_24206_, _24205_, _07143_);
  and (_24207_, _07144_, \oc8051_golden_model_1.TH1 [5]);
  or (_24208_, _24207_, _06285_);
  or (_24209_, _24208_, _24206_);
  and (_24211_, _24209_, _07169_);
  and (_24212_, _24211_, _24203_);
  and (_24213_, _09419_, _07900_);
  or (_24214_, _24213_, _24200_);
  and (_24215_, _24214_, _06354_);
  or (_24216_, _24215_, _24212_);
  and (_24217_, _24216_, _06346_);
  and (_24218_, _24205_, _06345_);
  or (_24219_, _24218_, _06259_);
  or (_24220_, _24219_, _24217_);
  or (_24222_, _24214_, _06260_);
  and (_24223_, _24222_, _24220_);
  or (_24224_, _24223_, _09486_);
  and (_24225_, _09436_, _07900_);
  or (_24226_, _24200_, _06258_);
  or (_24227_, _24226_, _24225_);
  and (_24228_, _24227_, _06251_);
  and (_24229_, _24228_, _24224_);
  and (_24230_, _15421_, _07900_);
  or (_24231_, _24230_, _24200_);
  and (_24233_, _24231_, _05972_);
  or (_24234_, _24233_, _10080_);
  or (_24235_, _24234_, _24229_);
  and (_24236_, _15313_, _07900_);
  or (_24237_, _24200_, _09025_);
  or (_24238_, _24237_, _24236_);
  and (_24239_, _08913_, _07900_);
  or (_24240_, _24239_, _24200_);
  or (_24241_, _24240_, _06216_);
  and (_24242_, _24241_, _09030_);
  and (_24244_, _24242_, _24238_);
  and (_24245_, _24244_, _24235_);
  and (_24246_, _12536_, _07900_);
  or (_24247_, _24246_, _24200_);
  and (_24248_, _24247_, _06524_);
  or (_24249_, _24248_, _24245_);
  and (_24250_, _24249_, _07219_);
  or (_24251_, _24200_, _08231_);
  and (_24252_, _24240_, _06426_);
  and (_24253_, _24252_, _24251_);
  or (_24255_, _24253_, _24250_);
  and (_24256_, _24255_, _07217_);
  and (_24257_, _24205_, _06532_);
  and (_24258_, _24257_, _24251_);
  or (_24259_, _24258_, _06437_);
  or (_24260_, _24259_, _24256_);
  and (_24261_, _15310_, _07900_);
  or (_24262_, _24200_, _07229_);
  or (_24263_, _24262_, _24261_);
  and (_24264_, _24263_, _07231_);
  and (_24265_, _24264_, _24260_);
  nor (_24266_, _11241_, _11961_);
  or (_24267_, _24266_, _24200_);
  and (_24268_, _24267_, _06535_);
  or (_24269_, _24268_, _06559_);
  or (_24270_, _24269_, _24265_);
  or (_24271_, _24202_, _07240_);
  and (_24272_, _24271_, _06570_);
  and (_24273_, _24272_, _24270_);
  and (_24274_, _15493_, _07900_);
  or (_24275_, _24274_, _24200_);
  and (_24276_, _24275_, _06566_);
  or (_24277_, _24276_, _01324_);
  or (_24278_, _24277_, _24273_);
  or (_24279_, _01320_, \oc8051_golden_model_1.TH1 [5]);
  and (_24280_, _24279_, _42355_);
  and (_42971_, _24280_, _24278_);
  and (_24281_, _11961_, \oc8051_golden_model_1.TH1 [6]);
  and (_24282_, _15521_, _07900_);
  or (_24283_, _24282_, _24281_);
  or (_24286_, _24283_, _06286_);
  and (_24287_, _07900_, \oc8051_golden_model_1.ACC [6]);
  or (_24288_, _24287_, _24281_);
  and (_24289_, _24288_, _07143_);
  and (_24290_, _07144_, \oc8051_golden_model_1.TH1 [6]);
  or (_24291_, _24290_, _06285_);
  or (_24292_, _24291_, _24289_);
  and (_24293_, _24292_, _07169_);
  and (_24294_, _24293_, _24286_);
  and (_24295_, _09418_, _07900_);
  or (_24297_, _24295_, _24281_);
  and (_24298_, _24297_, _06354_);
  or (_24299_, _24298_, _24294_);
  and (_24300_, _24299_, _06346_);
  and (_24301_, _24288_, _06345_);
  or (_24302_, _24301_, _06259_);
  or (_24303_, _24302_, _24300_);
  or (_24304_, _24297_, _06260_);
  and (_24305_, _24304_, _24303_);
  or (_24306_, _24305_, _09486_);
  and (_24308_, _09435_, _07900_);
  or (_24309_, _24281_, _06258_);
  or (_24310_, _24309_, _24308_);
  and (_24311_, _24310_, _06251_);
  and (_24312_, _24311_, _24306_);
  and (_24313_, _15623_, _07900_);
  or (_24314_, _24313_, _24281_);
  and (_24315_, _24314_, _05972_);
  or (_24316_, _24315_, _10080_);
  or (_24317_, _24316_, _24312_);
  and (_24319_, _15517_, _07900_);
  or (_24320_, _24281_, _09025_);
  or (_24321_, _24320_, _24319_);
  nor (_24322_, _08844_, _11961_);
  or (_24323_, _24322_, _24281_);
  or (_24324_, _24323_, _06216_);
  and (_24325_, _24324_, _09030_);
  and (_24326_, _24325_, _24321_);
  and (_24327_, _24326_, _24317_);
  and (_24328_, _11239_, _07900_);
  or (_24330_, _24328_, _24281_);
  and (_24331_, _24330_, _06524_);
  or (_24332_, _24331_, _24327_);
  and (_24333_, _24332_, _07219_);
  or (_24334_, _24281_, _08128_);
  and (_24335_, _24323_, _06426_);
  and (_24336_, _24335_, _24334_);
  or (_24337_, _24336_, _24333_);
  and (_24338_, _24337_, _07217_);
  and (_24339_, _24288_, _06532_);
  and (_24341_, _24339_, _24334_);
  or (_24342_, _24341_, _06437_);
  or (_24343_, _24342_, _24338_);
  and (_24344_, _15514_, _07900_);
  or (_24345_, _24281_, _07229_);
  or (_24346_, _24345_, _24344_);
  and (_24347_, _24346_, _07231_);
  and (_24348_, _24347_, _24343_);
  nor (_24349_, _11238_, _11961_);
  or (_24350_, _24349_, _24281_);
  and (_24352_, _24350_, _06535_);
  or (_24353_, _24352_, _06559_);
  or (_24354_, _24353_, _24348_);
  or (_24355_, _24283_, _07240_);
  and (_24356_, _24355_, _06570_);
  and (_24357_, _24356_, _24354_);
  and (_24358_, _15695_, _07900_);
  or (_24359_, _24358_, _24281_);
  and (_24360_, _24359_, _06566_);
  or (_24361_, _24360_, _01324_);
  or (_24363_, _24361_, _24357_);
  or (_24364_, _01320_, \oc8051_golden_model_1.TH1 [6]);
  and (_24365_, _24364_, _42355_);
  and (_42972_, _24365_, _24363_);
  and (_24366_, _01324_, \oc8051_golden_model_1.TH0 [0]);
  and (_24367_, _07908_, \oc8051_golden_model_1.ACC [0]);
  and (_24368_, _24367_, _08374_);
  and (_24369_, _12038_, \oc8051_golden_model_1.TH0 [0]);
  or (_24370_, _24369_, _07217_);
  or (_24371_, _24370_, _24368_);
  and (_24373_, _07908_, _07135_);
  or (_24374_, _24373_, _24369_);
  or (_24375_, _24374_, _06260_);
  nor (_24376_, _08374_, _12038_);
  or (_24377_, _24376_, _24369_);
  or (_24378_, _24377_, _06286_);
  or (_24379_, _24369_, _24367_);
  and (_24380_, _24379_, _07143_);
  and (_24381_, _07144_, \oc8051_golden_model_1.TH0 [0]);
  or (_24382_, _24381_, _06285_);
  or (_24384_, _24382_, _24380_);
  and (_24385_, _24384_, _07169_);
  and (_24386_, _24385_, _24378_);
  and (_24387_, _24374_, _06354_);
  or (_24388_, _24387_, _24386_);
  and (_24389_, _24388_, _06346_);
  and (_24390_, _24379_, _06345_);
  or (_24391_, _24390_, _06259_);
  or (_24392_, _24391_, _24389_);
  and (_24393_, _24392_, _24375_);
  or (_24395_, _24393_, _09486_);
  and (_24396_, _09384_, _07908_);
  or (_24397_, _24369_, _06258_);
  or (_24398_, _24397_, _24396_);
  and (_24399_, _24398_, _24395_);
  or (_24400_, _24399_, _05972_);
  and (_24401_, _14413_, _07908_);
  or (_24402_, _24369_, _06251_);
  or (_24403_, _24402_, _24401_);
  and (_24404_, _24403_, _06216_);
  and (_24406_, _24404_, _24400_);
  and (_24407_, _07908_, _08929_);
  or (_24408_, _24407_, _24369_);
  and (_24409_, _24408_, _06215_);
  or (_24410_, _24409_, _06398_);
  or (_24411_, _24410_, _24406_);
  and (_24412_, _14311_, _07908_);
  or (_24413_, _24412_, _24369_);
  or (_24414_, _24413_, _09025_);
  and (_24415_, _24414_, _09030_);
  and (_24417_, _24415_, _24411_);
  nor (_24418_, _12532_, _12038_);
  or (_24419_, _24418_, _24369_);
  nor (_24420_, _24368_, _09030_);
  and (_24421_, _24420_, _24419_);
  or (_24422_, _24421_, _24417_);
  and (_24423_, _24422_, _07219_);
  nand (_24424_, _24408_, _06426_);
  nor (_24425_, _24424_, _24376_);
  or (_24426_, _24425_, _06532_);
  or (_24428_, _24426_, _24423_);
  and (_24429_, _24428_, _24371_);
  or (_24430_, _24429_, _06437_);
  and (_24431_, _14307_, _07908_);
  or (_24432_, _24369_, _07229_);
  or (_24433_, _24432_, _24431_);
  and (_24434_, _24433_, _07231_);
  and (_24435_, _24434_, _24430_);
  and (_24436_, _24419_, _06535_);
  or (_24437_, _24436_, _19480_);
  or (_24439_, _24437_, _24435_);
  or (_24440_, _24377_, _06651_);
  and (_24441_, _24440_, _01320_);
  and (_24442_, _24441_, _24439_);
  or (_24443_, _24442_, _24366_);
  and (_42974_, _24443_, _42355_);
  not (_24444_, \oc8051_golden_model_1.TH0 [1]);
  nor (_24445_, _01320_, _24444_);
  nor (_24446_, _07908_, _24444_);
  and (_24447_, _07908_, _09422_);
  or (_24449_, _24447_, _24446_);
  or (_24450_, _24449_, _06260_);
  or (_24451_, _07908_, \oc8051_golden_model_1.TH0 [1]);
  and (_24452_, _14520_, _07908_);
  not (_24453_, _24452_);
  and (_24454_, _24453_, _24451_);
  or (_24455_, _24454_, _06286_);
  and (_24456_, _07908_, \oc8051_golden_model_1.ACC [1]);
  or (_24457_, _24456_, _24446_);
  and (_24458_, _24457_, _07143_);
  nor (_24460_, _07143_, _24444_);
  or (_24461_, _24460_, _06285_);
  or (_24462_, _24461_, _24458_);
  and (_24463_, _24462_, _07169_);
  and (_24464_, _24463_, _24455_);
  and (_24465_, _24449_, _06354_);
  or (_24466_, _24465_, _24464_);
  and (_24467_, _24466_, _06346_);
  and (_24468_, _24457_, _06345_);
  or (_24469_, _24468_, _06259_);
  or (_24471_, _24469_, _24467_);
  and (_24472_, _24471_, _24450_);
  or (_24473_, _24472_, _09486_);
  and (_24474_, _09339_, _07908_);
  or (_24475_, _24446_, _06258_);
  or (_24476_, _24475_, _24474_);
  and (_24477_, _24476_, _06251_);
  and (_24478_, _24477_, _24473_);
  or (_24479_, _14607_, _12038_);
  and (_24480_, _24451_, _05972_);
  and (_24482_, _24480_, _24479_);
  or (_24483_, _24482_, _24478_);
  and (_24484_, _24483_, _06399_);
  or (_24485_, _14505_, _12038_);
  and (_24486_, _24485_, _06398_);
  nand (_24487_, _07908_, _07031_);
  and (_24488_, _24487_, _06215_);
  or (_24489_, _24488_, _24486_);
  and (_24490_, _24489_, _24451_);
  or (_24491_, _24490_, _06524_);
  or (_24493_, _24491_, _24484_);
  nor (_24494_, _11252_, _12038_);
  or (_24495_, _24494_, _24446_);
  nand (_24496_, _11251_, _07908_);
  and (_24497_, _24496_, _24495_);
  or (_24498_, _24497_, _09030_);
  and (_24499_, _24498_, _07219_);
  and (_24500_, _24499_, _24493_);
  or (_24501_, _14503_, _12038_);
  and (_24502_, _24451_, _06426_);
  and (_24504_, _24502_, _24501_);
  or (_24505_, _24504_, _06532_);
  or (_24506_, _24505_, _24500_);
  nor (_24507_, _24446_, _07217_);
  nand (_24508_, _24507_, _24496_);
  and (_24509_, _24508_, _07229_);
  and (_24510_, _24509_, _24506_);
  or (_24511_, _24487_, _08325_);
  and (_24512_, _24451_, _06437_);
  and (_24513_, _24512_, _24511_);
  or (_24514_, _24513_, _06535_);
  or (_24515_, _24514_, _24510_);
  or (_24516_, _24495_, _07231_);
  and (_24517_, _24516_, _07240_);
  and (_24518_, _24517_, _24515_);
  and (_24519_, _24454_, _06559_);
  or (_24520_, _24519_, _06566_);
  or (_24521_, _24520_, _24518_);
  or (_24522_, _24446_, _06570_);
  or (_24523_, _24522_, _24452_);
  and (_24526_, _24523_, _01320_);
  and (_24527_, _24526_, _24521_);
  or (_24528_, _24527_, _24445_);
  and (_42975_, _24528_, _42355_);
  and (_24529_, _01324_, \oc8051_golden_model_1.TH0 [2]);
  and (_24530_, _12038_, \oc8051_golden_model_1.TH0 [2]);
  and (_24531_, _09293_, _07908_);
  or (_24532_, _24531_, _24530_);
  and (_24533_, _24532_, _09486_);
  and (_24534_, _14703_, _07908_);
  or (_24536_, _24534_, _24530_);
  or (_24537_, _24536_, _06286_);
  and (_24538_, _07908_, \oc8051_golden_model_1.ACC [2]);
  or (_24539_, _24538_, _24530_);
  and (_24540_, _24539_, _07143_);
  and (_24541_, _07144_, \oc8051_golden_model_1.TH0 [2]);
  or (_24542_, _24541_, _06285_);
  or (_24543_, _24542_, _24540_);
  and (_24544_, _24543_, _07169_);
  and (_24545_, _24544_, _24537_);
  and (_24547_, _07908_, _08662_);
  or (_24548_, _24547_, _24530_);
  and (_24549_, _24548_, _06354_);
  or (_24550_, _24549_, _24545_);
  and (_24551_, _24550_, _06346_);
  and (_24552_, _24539_, _06345_);
  or (_24553_, _24552_, _06259_);
  or (_24554_, _24553_, _24551_);
  or (_24555_, _24548_, _06260_);
  and (_24556_, _24555_, _06258_);
  and (_24558_, _24556_, _24554_);
  or (_24559_, _24558_, _05972_);
  or (_24560_, _24559_, _24533_);
  and (_24561_, _14804_, _07908_);
  or (_24562_, _24530_, _06251_);
  or (_24563_, _24562_, _24561_);
  and (_24564_, _24563_, _06216_);
  and (_24565_, _24564_, _24560_);
  and (_24566_, _07908_, _08980_);
  or (_24567_, _24566_, _24530_);
  and (_24569_, _24567_, _06215_);
  or (_24570_, _24569_, _06398_);
  or (_24571_, _24570_, _24565_);
  and (_24572_, _14697_, _07908_);
  or (_24573_, _24572_, _24530_);
  or (_24574_, _24573_, _09025_);
  and (_24575_, _24574_, _09030_);
  and (_24576_, _24575_, _24571_);
  and (_24577_, _11250_, _07908_);
  or (_24578_, _24577_, _24530_);
  and (_24580_, _24578_, _06524_);
  or (_24581_, _24580_, _24576_);
  and (_24582_, _24581_, _07219_);
  or (_24583_, _24530_, _08424_);
  and (_24584_, _24567_, _06426_);
  and (_24585_, _24584_, _24583_);
  or (_24586_, _24585_, _24582_);
  and (_24587_, _24586_, _07217_);
  and (_24588_, _24539_, _06532_);
  and (_24589_, _24588_, _24583_);
  or (_24591_, _24589_, _06437_);
  or (_24592_, _24591_, _24587_);
  and (_24593_, _14694_, _07908_);
  or (_24594_, _24530_, _07229_);
  or (_24595_, _24594_, _24593_);
  and (_24596_, _24595_, _07231_);
  and (_24597_, _24596_, _24592_);
  nor (_24598_, _11249_, _12038_);
  or (_24599_, _24598_, _24530_);
  and (_24600_, _24599_, _06535_);
  or (_24602_, _24600_, _24597_);
  and (_24603_, _24602_, _07240_);
  and (_24604_, _24536_, _06559_);
  or (_24605_, _24604_, _06566_);
  or (_24606_, _24605_, _24603_);
  and (_24607_, _14873_, _07908_);
  or (_24608_, _24530_, _06570_);
  or (_24609_, _24608_, _24607_);
  and (_24610_, _24609_, _01320_);
  and (_24611_, _24610_, _24606_);
  or (_24613_, _24611_, _24529_);
  and (_42976_, _24613_, _42355_);
  and (_24614_, _12038_, \oc8051_golden_model_1.TH0 [3]);
  and (_24615_, _14900_, _07908_);
  or (_24616_, _24615_, _24614_);
  or (_24617_, _24616_, _06286_);
  and (_24618_, _07908_, \oc8051_golden_model_1.ACC [3]);
  or (_24619_, _24618_, _24614_);
  and (_24620_, _24619_, _07143_);
  and (_24621_, _07144_, \oc8051_golden_model_1.TH0 [3]);
  or (_24623_, _24621_, _06285_);
  or (_24624_, _24623_, _24620_);
  and (_24625_, _24624_, _07169_);
  and (_24626_, _24625_, _24617_);
  and (_24627_, _07908_, _09421_);
  or (_24628_, _24627_, _24614_);
  and (_24629_, _24628_, _06354_);
  or (_24630_, _24629_, _24626_);
  and (_24631_, _24630_, _06346_);
  and (_24632_, _24619_, _06345_);
  or (_24634_, _24632_, _06259_);
  or (_24635_, _24634_, _24631_);
  or (_24636_, _24628_, _06260_);
  and (_24637_, _24636_, _24635_);
  or (_24638_, _24637_, _09486_);
  and (_24639_, _09247_, _07908_);
  or (_24640_, _24614_, _06258_);
  or (_24641_, _24640_, _24639_);
  and (_24642_, _24641_, _06251_);
  and (_24643_, _24642_, _24638_);
  and (_24645_, _14998_, _07908_);
  or (_24646_, _24645_, _24614_);
  and (_24647_, _24646_, _05972_);
  or (_24648_, _24647_, _10080_);
  or (_24649_, _24648_, _24643_);
  and (_24650_, _14893_, _07908_);
  or (_24651_, _24614_, _09025_);
  or (_24652_, _24651_, _24650_);
  and (_24653_, _07908_, _08809_);
  or (_24654_, _24653_, _24614_);
  or (_24656_, _24654_, _06216_);
  and (_24657_, _24656_, _09030_);
  and (_24658_, _24657_, _24652_);
  and (_24659_, _24658_, _24649_);
  and (_24660_, _12529_, _07908_);
  or (_24661_, _24660_, _24614_);
  and (_24662_, _24661_, _06524_);
  or (_24663_, _24662_, _24659_);
  and (_24664_, _24663_, _07219_);
  or (_24665_, _24614_, _08280_);
  and (_24667_, _24654_, _06426_);
  and (_24668_, _24667_, _24665_);
  or (_24669_, _24668_, _24664_);
  and (_24670_, _24669_, _07217_);
  and (_24671_, _24619_, _06532_);
  and (_24672_, _24671_, _24665_);
  or (_24673_, _24672_, _06437_);
  or (_24674_, _24673_, _24670_);
  and (_24675_, _14890_, _07908_);
  or (_24676_, _24614_, _07229_);
  or (_24678_, _24676_, _24675_);
  and (_24679_, _24678_, _07231_);
  and (_24680_, _24679_, _24674_);
  nor (_24681_, _11247_, _12038_);
  or (_24682_, _24681_, _24614_);
  and (_24683_, _24682_, _06535_);
  or (_24684_, _24683_, _06559_);
  or (_24685_, _24684_, _24680_);
  or (_24686_, _24616_, _07240_);
  and (_24687_, _24686_, _06570_);
  and (_24689_, _24687_, _24685_);
  and (_24690_, _15068_, _07908_);
  or (_24691_, _24690_, _24614_);
  and (_24692_, _24691_, _06566_);
  or (_24693_, _24692_, _01324_);
  or (_24694_, _24693_, _24689_);
  or (_24695_, _01320_, \oc8051_golden_model_1.TH0 [3]);
  and (_24696_, _24695_, _42355_);
  and (_42977_, _24696_, _24694_);
  and (_24697_, _12038_, \oc8051_golden_model_1.TH0 [4]);
  and (_24699_, _09420_, _07908_);
  or (_24700_, _24699_, _24697_);
  or (_24701_, _24700_, _06260_);
  and (_24702_, _15133_, _07908_);
  or (_24703_, _24702_, _24697_);
  or (_24704_, _24703_, _06286_);
  and (_24705_, _07908_, \oc8051_golden_model_1.ACC [4]);
  or (_24706_, _24705_, _24697_);
  and (_24707_, _24706_, _07143_);
  and (_24708_, _07144_, \oc8051_golden_model_1.TH0 [4]);
  or (_24710_, _24708_, _06285_);
  or (_24711_, _24710_, _24707_);
  and (_24712_, _24711_, _07169_);
  and (_24713_, _24712_, _24704_);
  and (_24714_, _24700_, _06354_);
  or (_24715_, _24714_, _24713_);
  and (_24716_, _24715_, _06346_);
  and (_24717_, _24706_, _06345_);
  or (_24718_, _24717_, _06259_);
  or (_24719_, _24718_, _24716_);
  and (_24721_, _24719_, _24701_);
  or (_24722_, _24721_, _09486_);
  and (_24723_, _09437_, _07908_);
  or (_24724_, _24697_, _06258_);
  or (_24725_, _24724_, _24723_);
  and (_24726_, _24725_, _06251_);
  and (_24727_, _24726_, _24722_);
  and (_24728_, _15226_, _07908_);
  or (_24729_, _24728_, _24697_);
  and (_24730_, _24729_, _05972_);
  or (_24732_, _24730_, _24727_);
  or (_24733_, _24732_, _10080_);
  and (_24734_, _15114_, _07908_);
  or (_24735_, _24697_, _09025_);
  or (_24736_, _24735_, _24734_);
  and (_24737_, _08919_, _07908_);
  or (_24738_, _24737_, _24697_);
  or (_24739_, _24738_, _06216_);
  and (_24740_, _24739_, _09030_);
  and (_24741_, _24740_, _24736_);
  and (_24743_, _24741_, _24733_);
  and (_24744_, _11245_, _07908_);
  or (_24745_, _24744_, _24697_);
  and (_24746_, _24745_, _06524_);
  or (_24747_, _24746_, _24743_);
  and (_24748_, _24747_, _07219_);
  or (_24749_, _24697_, _08528_);
  and (_24750_, _24738_, _06426_);
  and (_24751_, _24750_, _24749_);
  or (_24752_, _24751_, _24748_);
  and (_24754_, _24752_, _07217_);
  and (_24755_, _24706_, _06532_);
  and (_24756_, _24755_, _24749_);
  or (_24757_, _24756_, _06437_);
  or (_24758_, _24757_, _24754_);
  and (_24759_, _15111_, _07908_);
  or (_24760_, _24697_, _07229_);
  or (_24761_, _24760_, _24759_);
  and (_24762_, _24761_, _07231_);
  and (_24763_, _24762_, _24758_);
  nor (_24765_, _11244_, _12038_);
  or (_24766_, _24765_, _24697_);
  and (_24767_, _24766_, _06535_);
  or (_24768_, _24767_, _06559_);
  or (_24769_, _24768_, _24763_);
  or (_24770_, _24703_, _07240_);
  and (_24771_, _24770_, _06570_);
  and (_24772_, _24771_, _24769_);
  and (_24773_, _15296_, _07908_);
  or (_24774_, _24773_, _24697_);
  and (_24776_, _24774_, _06566_);
  or (_24777_, _24776_, _01324_);
  or (_24778_, _24777_, _24772_);
  or (_24779_, _01320_, \oc8051_golden_model_1.TH0 [4]);
  and (_24780_, _24779_, _42355_);
  and (_42978_, _24780_, _24778_);
  and (_24781_, _12038_, \oc8051_golden_model_1.TH0 [5]);
  and (_24782_, _15330_, _07908_);
  or (_24783_, _24782_, _24781_);
  or (_24784_, _24783_, _06286_);
  and (_24786_, _07908_, \oc8051_golden_model_1.ACC [5]);
  or (_24787_, _24786_, _24781_);
  and (_24788_, _24787_, _07143_);
  and (_24789_, _07144_, \oc8051_golden_model_1.TH0 [5]);
  or (_24790_, _24789_, _06285_);
  or (_24791_, _24790_, _24788_);
  and (_24792_, _24791_, _07169_);
  and (_24793_, _24792_, _24784_);
  and (_24794_, _09419_, _07908_);
  or (_24795_, _24794_, _24781_);
  and (_24797_, _24795_, _06354_);
  or (_24798_, _24797_, _24793_);
  and (_24799_, _24798_, _06346_);
  and (_24800_, _24787_, _06345_);
  or (_24801_, _24800_, _06259_);
  or (_24802_, _24801_, _24799_);
  or (_24803_, _24795_, _06260_);
  and (_24804_, _24803_, _24802_);
  or (_24805_, _24804_, _09486_);
  and (_24806_, _09436_, _07908_);
  or (_24808_, _24781_, _06258_);
  or (_24809_, _24808_, _24806_);
  and (_24810_, _24809_, _06251_);
  and (_24811_, _24810_, _24805_);
  and (_24812_, _15421_, _07908_);
  or (_24813_, _24812_, _24781_);
  and (_24814_, _24813_, _05972_);
  or (_24815_, _24814_, _10080_);
  or (_24816_, _24815_, _24811_);
  and (_24817_, _15313_, _07908_);
  or (_24819_, _24781_, _09025_);
  or (_24820_, _24819_, _24817_);
  and (_24821_, _08913_, _07908_);
  or (_24822_, _24821_, _24781_);
  or (_24823_, _24822_, _06216_);
  and (_24824_, _24823_, _09030_);
  and (_24825_, _24824_, _24820_);
  and (_24826_, _24825_, _24816_);
  and (_24827_, _12536_, _07908_);
  or (_24828_, _24827_, _24781_);
  and (_24830_, _24828_, _06524_);
  or (_24831_, _24830_, _24826_);
  and (_24832_, _24831_, _07219_);
  or (_24833_, _24781_, _08231_);
  and (_24834_, _24822_, _06426_);
  and (_24835_, _24834_, _24833_);
  or (_24836_, _24835_, _24832_);
  and (_24837_, _24836_, _07217_);
  and (_24838_, _24787_, _06532_);
  and (_24839_, _24838_, _24833_);
  or (_24841_, _24839_, _06437_);
  or (_24842_, _24841_, _24837_);
  and (_24843_, _15310_, _07908_);
  or (_24844_, _24781_, _07229_);
  or (_24845_, _24844_, _24843_);
  and (_24846_, _24845_, _07231_);
  and (_24847_, _24846_, _24842_);
  nor (_24848_, _11241_, _12038_);
  or (_24849_, _24848_, _24781_);
  and (_24850_, _24849_, _06535_);
  or (_24852_, _24850_, _06559_);
  or (_24853_, _24852_, _24847_);
  or (_24854_, _24783_, _07240_);
  and (_24855_, _24854_, _06570_);
  and (_24856_, _24855_, _24853_);
  and (_24857_, _15493_, _07908_);
  or (_24858_, _24857_, _24781_);
  and (_24859_, _24858_, _06566_);
  or (_24860_, _24859_, _01324_);
  or (_24861_, _24860_, _24856_);
  or (_24863_, _01320_, \oc8051_golden_model_1.TH0 [5]);
  and (_24864_, _24863_, _42355_);
  and (_42980_, _24864_, _24861_);
  and (_24865_, _12038_, \oc8051_golden_model_1.TH0 [6]);
  and (_24866_, _15521_, _07908_);
  or (_24867_, _24866_, _24865_);
  or (_24868_, _24867_, _06286_);
  and (_24869_, _07908_, \oc8051_golden_model_1.ACC [6]);
  or (_24870_, _24869_, _24865_);
  and (_24871_, _24870_, _07143_);
  and (_24873_, _07144_, \oc8051_golden_model_1.TH0 [6]);
  or (_24874_, _24873_, _06285_);
  or (_24875_, _24874_, _24871_);
  and (_24876_, _24875_, _07169_);
  and (_24877_, _24876_, _24868_);
  and (_24878_, _09418_, _07908_);
  or (_24879_, _24878_, _24865_);
  and (_24880_, _24879_, _06354_);
  or (_24881_, _24880_, _24877_);
  and (_24882_, _24881_, _06346_);
  and (_24884_, _24870_, _06345_);
  or (_24885_, _24884_, _06259_);
  or (_24886_, _24885_, _24882_);
  or (_24887_, _24879_, _06260_);
  and (_24888_, _24887_, _24886_);
  or (_24889_, _24888_, _09486_);
  and (_24890_, _09435_, _07908_);
  or (_24891_, _24865_, _06258_);
  or (_24892_, _24891_, _24890_);
  and (_24893_, _24892_, _06251_);
  and (_24895_, _24893_, _24889_);
  and (_24896_, _15623_, _07908_);
  or (_24897_, _24896_, _24865_);
  and (_24898_, _24897_, _05972_);
  or (_24899_, _24898_, _10080_);
  or (_24900_, _24899_, _24895_);
  and (_24901_, _15517_, _07908_);
  or (_24902_, _24865_, _09025_);
  or (_24903_, _24902_, _24901_);
  and (_24904_, _08845_, _07908_);
  or (_24906_, _24904_, _24865_);
  or (_24907_, _24906_, _06216_);
  and (_24908_, _24907_, _09030_);
  and (_24909_, _24908_, _24903_);
  and (_24910_, _24909_, _24900_);
  and (_24911_, _11239_, _07908_);
  or (_24912_, _24911_, _24865_);
  and (_24913_, _24912_, _06524_);
  or (_24914_, _24913_, _24910_);
  and (_24915_, _24914_, _07219_);
  or (_24917_, _24865_, _08128_);
  and (_24918_, _24906_, _06426_);
  and (_24919_, _24918_, _24917_);
  or (_24920_, _24919_, _24915_);
  and (_24921_, _24920_, _07217_);
  and (_24922_, _24870_, _06532_);
  and (_24923_, _24922_, _24917_);
  or (_24924_, _24923_, _06437_);
  or (_24925_, _24924_, _24921_);
  and (_24926_, _15514_, _07908_);
  or (_24928_, _24865_, _07229_);
  or (_24929_, _24928_, _24926_);
  and (_24930_, _24929_, _07231_);
  and (_24931_, _24930_, _24925_);
  nor (_24932_, _11238_, _12038_);
  or (_24933_, _24932_, _24865_);
  and (_24934_, _24933_, _06535_);
  or (_24935_, _24934_, _06559_);
  or (_24936_, _24935_, _24931_);
  or (_24937_, _24867_, _07240_);
  and (_24939_, _24937_, _06570_);
  and (_24940_, _24939_, _24936_);
  and (_24941_, _15695_, _07908_);
  or (_24942_, _24941_, _24865_);
  and (_24943_, _24942_, _06566_);
  or (_24944_, _24943_, _01324_);
  or (_24945_, _24944_, _24940_);
  or (_24946_, _01320_, \oc8051_golden_model_1.TH0 [6]);
  and (_24947_, _24946_, _42355_);
  and (_42981_, _24947_, _24945_);
  and (_24949_, _13027_, _13019_);
  or (_24950_, _24949_, _05619_);
  and (_24951_, _12998_, _13005_);
  or (_24952_, _24951_, _05619_);
  and (_24953_, _12129_, _12981_);
  or (_24954_, _24953_, _05619_);
  and (_24955_, _12749_, _07229_);
  or (_24956_, _24955_, _05619_);
  and (_24957_, _12244_, _07219_);
  or (_24958_, _24957_, _05619_);
  and (_24960_, _12695_, _09025_);
  or (_24961_, _24960_, _05619_);
  nand (_24962_, _12540_, \oc8051_golden_model_1.PC [0]);
  and (_24963_, _06850_, \oc8051_golden_model_1.PC [0]);
  nor (_24964_, _24963_, _12319_);
  or (_24965_, _24964_, _12540_);
  and (_24966_, _24965_, _06347_);
  and (_24967_, _24966_, _24962_);
  and (_24968_, _12400_, _05619_);
  and (_24969_, _24964_, _12398_);
  or (_24971_, _24969_, _06424_);
  or (_24972_, _24971_, _24968_);
  nand (_24973_, _06850_, _07152_);
  nand (_24974_, _12448_, \oc8051_golden_model_1.PC [0]);
  and (_24975_, _07454_, _06756_);
  or (_24976_, _24975_, _05619_);
  nand (_24977_, _24975_, _05619_);
  nand (_24978_, _24977_, _24976_);
  nor (_24979_, _12448_, _07152_);
  nand (_24980_, _24979_, _24978_);
  and (_24982_, _24980_, _24974_);
  and (_24983_, _24982_, _24973_);
  or (_24984_, _24983_, _08734_);
  and (_24985_, _12430_, \oc8051_golden_model_1.PC [0]);
  nor (_24986_, _06248_, \oc8051_golden_model_1.PC [0]);
  nor (_24987_, _24986_, _12189_);
  and (_24988_, _24987_, _12432_);
  or (_24989_, _24988_, _24985_);
  or (_24990_, _24989_, _08736_);
  and (_24991_, _24990_, _24984_);
  or (_24993_, _24991_, _07159_);
  nand (_24994_, _07159_, \oc8051_golden_model_1.PC [0]);
  and (_24995_, _24994_, _06286_);
  and (_24996_, _24995_, _24993_);
  or (_24997_, _12420_, _05619_);
  or (_24998_, _24964_, _12418_);
  and (_24999_, _24998_, _06285_);
  and (_25000_, _24999_, _24997_);
  or (_25001_, _25000_, _12410_);
  or (_25002_, _25001_, _24996_);
  or (_25004_, _12409_, _05619_);
  and (_25005_, _25004_, _05949_);
  and (_25006_, _25005_, _25002_);
  or (_25007_, _06850_, _05949_);
  and (_25008_, _12468_, _12404_);
  nand (_25009_, _25008_, _25007_);
  or (_25010_, _25009_, _25006_);
  or (_25011_, _25008_, _05619_);
  and (_25012_, _25011_, _05955_);
  and (_25013_, _25012_, _25010_);
  nor (_25015_, _06850_, _05955_);
  or (_25016_, _25015_, _12485_);
  or (_25017_, _25016_, _25013_);
  and (_25018_, _12519_, _05619_);
  not (_25019_, _12519_);
  and (_25020_, _24964_, _25019_);
  or (_25021_, _25020_, _12484_);
  or (_25022_, _25021_, _25018_);
  and (_25023_, _25022_, _25017_);
  or (_25024_, _25023_, _06423_);
  and (_25026_, _25024_, _14105_);
  and (_25027_, _25026_, _24972_);
  or (_25028_, _25027_, _24967_);
  and (_25029_, _25028_, _12528_);
  nand (_25030_, _12559_, \oc8051_golden_model_1.PC [0]);
  or (_25031_, _24964_, _12559_);
  and (_25032_, _25031_, _06419_);
  and (_25033_, _25032_, _25030_);
  or (_25034_, _25033_, _12254_);
  or (_25035_, _25034_, _25029_);
  nand (_25037_, _12254_, \oc8051_golden_model_1.PC [0]);
  and (_25038_, _25037_, _05946_);
  and (_25039_, _25038_, _25035_);
  nor (_25040_, _06850_, _05946_);
  or (_25041_, _25040_, _12589_);
  or (_25042_, _25041_, _25039_);
  or (_25043_, _12585_, _05619_);
  and (_25044_, _25043_, _05953_);
  and (_25045_, _25044_, _25042_);
  or (_25046_, _06850_, _05953_);
  and (_25048_, _12595_, _05940_);
  nand (_25049_, _25048_, _25046_);
  or (_25050_, _25049_, _25045_);
  or (_25051_, _25048_, _05619_);
  and (_25052_, _25051_, _15174_);
  and (_25053_, _25052_, _25050_);
  or (_25054_, _06850_, _15174_);
  nor (_25055_, _06395_, _05972_);
  and (_25056_, _25055_, _12252_);
  nand (_25057_, _25056_, _25054_);
  or (_25058_, _25057_, _25053_);
  or (_25059_, _25056_, _05619_);
  and (_25060_, _25059_, _05998_);
  and (_25061_, _25060_, _25058_);
  nor (_25062_, _06850_, _05998_);
  or (_25063_, _25062_, _12630_);
  or (_25064_, _25063_, _25061_);
  or (_25065_, _24987_, _12631_);
  and (_25066_, _25065_, _25064_);
  or (_25067_, _25066_, _06215_);
  and (_25070_, _06215_, \oc8051_golden_model_1.PC [0]);
  nor (_25071_, _12644_, _25070_);
  and (_25072_, _25071_, _25067_);
  and (_25073_, _12644_, _05979_);
  or (_25074_, _25073_, _06004_);
  or (_25075_, _25074_, _25072_);
  nand (_25076_, _06850_, _06004_);
  and (_25077_, _25076_, _12685_);
  and (_25078_, _25077_, _25075_);
  or (_25079_, _24987_, _11327_);
  nand (_25081_, _11327_, _05619_);
  and (_25082_, _25081_, _12247_);
  nand (_25083_, _25082_, _25079_);
  nand (_25084_, _25083_, _24960_);
  or (_25085_, _25084_, _25078_);
  and (_25086_, _25085_, _24961_);
  or (_25087_, _25086_, _06001_);
  nand (_25088_, _06850_, _06001_);
  and (_25089_, _25088_, _12712_);
  and (_25090_, _25089_, _25087_);
  or (_25092_, _24987_, _12248_);
  or (_25093_, _11327_, \oc8051_golden_model_1.PC [0]);
  and (_25094_, _25093_, _12711_);
  nand (_25095_, _25094_, _25092_);
  nand (_25096_, _25095_, _24957_);
  or (_25097_, _25096_, _25090_);
  and (_25098_, _25097_, _24958_);
  or (_25099_, _25098_, _06013_);
  nand (_25100_, _06850_, _06013_);
  and (_25101_, _25100_, _12733_);
  and (_25103_, _25101_, _25099_);
  or (_25104_, _24987_, \oc8051_golden_model_1.PSW [7]);
  or (_25105_, _10774_, \oc8051_golden_model_1.PC [0]);
  and (_25106_, _25105_, _12732_);
  nand (_25107_, _25106_, _25104_);
  nand (_25108_, _25107_, _24955_);
  or (_25109_, _25108_, _25103_);
  and (_25110_, _25109_, _24956_);
  or (_25111_, _25110_, _06008_);
  nand (_25112_, _06850_, _06008_);
  and (_25114_, _25112_, _12762_);
  and (_25115_, _25114_, _25111_);
  nor (_25116_, _08786_, _05619_);
  and (_25117_, _08786_, _05619_);
  or (_25118_, _25117_, _25116_);
  nand (_25119_, _25118_, _12239_);
  and (_25120_, _12767_, _12775_);
  nand (_25121_, _25120_, _25119_);
  or (_25122_, _25121_, _25115_);
  or (_25123_, _25120_, _05619_);
  and (_25125_, _25123_, _12782_);
  and (_25126_, _25125_, _25122_);
  and (_25127_, _09384_, _06543_);
  or (_25128_, _25127_, _06011_);
  or (_25129_, _25128_, _25126_);
  nand (_25130_, _06850_, _06011_);
  and (_25131_, _25130_, _12786_);
  and (_25132_, _25131_, _25129_);
  not (_25133_, _12970_);
  or (_25134_, _24964_, _25133_);
  or (_25136_, _12970_, _05619_);
  and (_25137_, _25136_, _06436_);
  nand (_25138_, _25137_, _25134_);
  nand (_25139_, _25138_, _24953_);
  or (_25140_, _25139_, _25132_);
  and (_25141_, _25140_, _24954_);
  or (_25142_, _25141_, _06290_);
  not (_25143_, _05994_);
  or (_25144_, _09384_, _06291_);
  and (_25145_, _25144_, _25143_);
  and (_25147_, _25145_, _25142_);
  nor (_25148_, _06850_, _25143_);
  or (_25149_, _25148_, _25147_);
  and (_25150_, _25149_, _06435_);
  nand (_25151_, _12970_, \oc8051_golden_model_1.PC [0]);
  or (_25152_, _24964_, _12970_);
  and (_25153_, _25152_, _25151_);
  nand (_25154_, _25153_, _06434_);
  nand (_25155_, _25154_, _24951_);
  or (_25156_, _25155_, _25150_);
  and (_25158_, _25156_, _24952_);
  or (_25159_, _25158_, _07678_);
  nand (_25160_, _07678_, _06850_);
  and (_25161_, _25160_, _05933_);
  and (_25162_, _25161_, _25159_);
  nand (_25163_, _25153_, _05932_);
  nand (_25164_, _25163_, _24949_);
  or (_25165_, _25164_, _25162_);
  and (_25166_, _25165_, _24950_);
  nor (_25167_, _06393_, _05989_);
  not (_25169_, _25167_);
  or (_25170_, _25169_, _25166_);
  nand (_25171_, _25169_, _06850_);
  and (_25172_, _25171_, _13039_);
  and (_25173_, _25172_, _25170_);
  and (_25174_, _13035_, _05619_);
  or (_25175_, _25174_, _01324_);
  or (_25176_, _25175_, _25173_);
  or (_25177_, _01320_, \oc8051_golden_model_1.PC [0]);
  and (_25178_, _25177_, _42355_);
  and (_42983_, _25178_, _25176_);
  and (_25180_, _06566_, _05585_);
  and (_25181_, _06559_, _05585_);
  or (_25182_, _08547_, _06035_);
  or (_25183_, _12129_, _06035_);
  or (_25184_, _12767_, _06035_);
  nand (_25185_, _12745_, _06034_);
  or (_25186_, _12244_, _06035_);
  or (_25187_, _12695_, _06035_);
  or (_25188_, _09015_, _05585_);
  or (_25190_, _12595_, _06035_);
  nand (_25191_, _12254_, _06034_);
  or (_25192_, _12321_, _12319_);
  and (_25193_, _25192_, _12322_);
  or (_25194_, _25193_, _12519_);
  nand (_25195_, _12519_, _06035_);
  and (_25196_, _25195_, _25194_);
  or (_25197_, _25196_, _12484_);
  nor (_25198_, _07031_, _05955_);
  or (_25199_, _12468_, _06035_);
  or (_25201_, _12425_, _12428_);
  or (_25202_, _12427_, _12424_);
  or (_25203_, _25202_, _25201_);
  nor (_25204_, _12191_, _12189_);
  nor (_25205_, _25204_, _12192_);
  and (_25206_, _25205_, _25203_);
  and (_25207_, _12430_, _05585_);
  or (_25208_, _25207_, _25206_);
  or (_25209_, _25208_, _08736_);
  nand (_25210_, _07031_, _07152_);
  nand (_25212_, _12448_, _06034_);
  not (_25213_, _24979_);
  and (_25214_, _06755_, _05619_);
  nor (_25215_, _07454_, _05619_);
  nor (_25216_, _25215_, _07143_);
  and (_25217_, _25216_, _06756_);
  nor (_25218_, _25217_, _25214_);
  nand (_25219_, _25218_, \oc8051_golden_model_1.PC [1]);
  or (_25220_, _25218_, \oc8051_golden_model_1.PC [1]);
  and (_25221_, _25220_, _25219_);
  or (_25223_, _25221_, _25213_);
  and (_25224_, _25223_, _25212_);
  and (_25225_, _25224_, _25210_);
  or (_25226_, _25225_, _08734_);
  and (_25227_, _25226_, _08639_);
  and (_25228_, _25227_, _25209_);
  and (_25229_, _07159_, _06035_);
  or (_25230_, _25229_, _06285_);
  or (_25231_, _25230_, _25228_);
  and (_25232_, _25193_, _12420_);
  and (_25234_, _12418_, _06034_);
  or (_25235_, _25234_, _06286_);
  or (_25236_, _25235_, _25232_);
  and (_25237_, _25236_, _25231_);
  or (_25238_, _25237_, _12410_);
  or (_25239_, _12409_, _06035_);
  and (_25240_, _25239_, _06282_);
  and (_25241_, _25240_, _25238_);
  and (_25242_, _06281_, _05585_);
  or (_25243_, _25242_, _07460_);
  or (_25245_, _25243_, _25241_);
  nand (_25246_, _07031_, _07460_);
  and (_25247_, _25246_, _07169_);
  and (_25248_, _25247_, _25245_);
  nand (_25249_, _06354_, _05585_);
  nand (_25250_, _25249_, _12404_);
  or (_25251_, _25250_, _25248_);
  or (_25252_, _12404_, _06035_);
  and (_25253_, _25252_, _06346_);
  and (_25254_, _25253_, _25251_);
  nand (_25256_, _06345_, _05585_);
  nand (_25257_, _25256_, _12468_);
  or (_25258_, _25257_, _25254_);
  and (_25259_, _25258_, _25199_);
  or (_25260_, _25259_, _06277_);
  nand (_25261_, _06277_, \oc8051_golden_model_1.PC [1]);
  and (_25262_, _25261_, _05955_);
  and (_25263_, _25262_, _25260_);
  or (_25264_, _25263_, _25198_);
  and (_25265_, _25264_, _06778_);
  nand (_25267_, _06276_, _05585_);
  nand (_25268_, _25267_, _12484_);
  or (_25269_, _25268_, _25265_);
  and (_25270_, _25269_, _25197_);
  or (_25271_, _25270_, _06423_);
  and (_25272_, _25193_, _12398_);
  and (_25273_, _12400_, _06034_);
  or (_25274_, _25273_, _06424_);
  or (_25275_, _25274_, _25272_);
  and (_25276_, _25275_, _14105_);
  and (_25278_, _25276_, _25271_);
  not (_25279_, _12540_);
  and (_25280_, _25193_, _25279_);
  and (_25281_, _12540_, _06034_);
  or (_25282_, _25281_, _25280_);
  and (_25283_, _25282_, _06347_);
  or (_25284_, _25283_, _25278_);
  and (_25285_, _25284_, _12528_);
  or (_25286_, _25193_, _12559_);
  nand (_25287_, _12559_, _06035_);
  and (_25289_, _25287_, _06419_);
  and (_25290_, _25289_, _25286_);
  or (_25291_, _25290_, _12254_);
  or (_25292_, _25291_, _25285_);
  and (_25293_, _25292_, _25191_);
  or (_25294_, _25293_, _06270_);
  nand (_25295_, _06270_, \oc8051_golden_model_1.PC [1]);
  and (_25296_, _25295_, _05946_);
  and (_25297_, _25296_, _25294_);
  nor (_25298_, _07031_, _05946_);
  not (_25300_, _07374_);
  nor (_25301_, _07034_, _05952_);
  not (_25302_, _25301_);
  and (_25303_, _25302_, _12572_);
  and (_25304_, _25303_, _25300_);
  not (_25305_, _25304_);
  or (_25306_, _25305_, _25298_);
  or (_25307_, _25306_, _25297_);
  or (_25308_, _25304_, _05585_);
  and (_25309_, _25308_, _12583_);
  and (_25311_, _25309_, _25307_);
  nand (_25312_, _12582_, _06035_);
  nand (_25313_, _25312_, _12584_);
  or (_25314_, _25313_, _25311_);
  or (_25315_, _12584_, _06035_);
  and (_25316_, _25315_, _14014_);
  and (_25317_, _25316_, _25314_);
  not (_25318_, _05953_);
  and (_25319_, _06371_, _05585_);
  or (_25320_, _25319_, _25318_);
  or (_25321_, _25320_, _25317_);
  nand (_25322_, _07031_, _25318_);
  and (_25323_, _25322_, _14013_);
  and (_25324_, _25323_, _25321_);
  nand (_25325_, _10555_, _06803_);
  and (_25326_, _06370_, _05585_);
  or (_25327_, _25326_, _10718_);
  nor (_25328_, _25327_, _25325_);
  nand (_25329_, _25328_, _14151_);
  or (_25330_, _25329_, _25324_);
  and (_25333_, _25330_, _25190_);
  or (_25334_, _25333_, _12600_);
  or (_25335_, _12599_, _05585_);
  and (_25336_, _25335_, _05940_);
  and (_25337_, _25336_, _25334_);
  nor (_25338_, _06034_, _05940_);
  or (_25339_, _25338_, _06266_);
  or (_25340_, _25339_, _25337_);
  nand (_25341_, _06266_, \oc8051_golden_model_1.PC [1]);
  and (_25342_, _25341_, _25340_);
  or (_25344_, _25342_, _05974_);
  nand (_25345_, _07031_, _05974_);
  and (_25346_, _25345_, _06396_);
  and (_25347_, _25346_, _25344_);
  nand (_25348_, _06395_, _06034_);
  nand (_25349_, _25348_, _06261_);
  or (_25350_, _25349_, _25347_);
  or (_25351_, _06261_, _05585_);
  and (_25352_, _25351_, _06251_);
  and (_25353_, _25352_, _25350_);
  nand (_25355_, _06034_, _05972_);
  nand (_25356_, _25355_, _12252_);
  or (_25357_, _25356_, _25353_);
  or (_25358_, _12252_, _06035_);
  and (_25359_, _25358_, _06854_);
  and (_25360_, _25359_, _25357_);
  and (_25361_, _06330_, _05585_);
  or (_25362_, _25361_, _05997_);
  or (_25363_, _25362_, _25360_);
  nand (_25364_, _07031_, _05997_);
  and (_25366_, _25364_, _12631_);
  and (_25367_, _25366_, _25363_);
  and (_25368_, _25205_, _12630_);
  or (_25369_, _25368_, _09016_);
  or (_25370_, _25369_, _25367_);
  and (_25371_, _25370_, _25188_);
  or (_25372_, _25371_, _06215_);
  nand (_25373_, _06215_, _06035_);
  and (_25374_, _25373_, _10892_);
  and (_25375_, _25374_, _25372_);
  and (_25377_, _10891_, _05585_);
  or (_25378_, _25377_, _12644_);
  or (_25379_, _25378_, _25375_);
  not (_25380_, _12644_);
  or (_25381_, _25380_, _06032_);
  and (_25382_, _25381_, _06860_);
  and (_25383_, _25382_, _25379_);
  and (_25384_, _06329_, _05585_);
  or (_25385_, _25384_, _06004_);
  or (_25386_, _25385_, _25383_);
  nand (_25388_, _07031_, _06004_);
  and (_25389_, _25388_, _12685_);
  and (_25390_, _25389_, _25386_);
  or (_25391_, _25205_, _11327_);
  nand (_25392_, _11327_, \oc8051_golden_model_1.PC [1]);
  and (_25393_, _25392_, _12247_);
  and (_25394_, _25393_, _25391_);
  or (_25395_, _25394_, _12697_);
  or (_25396_, _25395_, _25390_);
  and (_25397_, _25396_, _25187_);
  or (_25399_, _25397_, _12700_);
  or (_25400_, _12699_, _05585_);
  and (_25401_, _25400_, _09025_);
  and (_25402_, _25401_, _25399_);
  and (_25403_, _06398_, _06034_);
  or (_25404_, _25403_, _06524_);
  or (_25405_, _25404_, _25402_);
  nand (_25406_, _06524_, \oc8051_golden_model_1.PC [1]);
  and (_25407_, _25406_, _25405_);
  or (_25408_, _25407_, _06001_);
  nand (_25410_, _07031_, _06001_);
  and (_25411_, _25410_, _12712_);
  and (_25412_, _25411_, _25408_);
  or (_25413_, _25205_, _12248_);
  or (_25414_, _11327_, _05585_);
  and (_25415_, _25414_, _12711_);
  and (_25416_, _25415_, _25413_);
  or (_25417_, _25416_, _12720_);
  or (_25418_, _25417_, _25412_);
  and (_25419_, _25418_, _25186_);
  or (_25421_, _25419_, _10970_);
  or (_25422_, _10969_, _05585_);
  and (_25423_, _25422_, _07219_);
  and (_25424_, _25423_, _25421_);
  and (_25425_, _06426_, _06034_);
  or (_25426_, _25425_, _06532_);
  or (_25427_, _25426_, _25424_);
  nand (_25428_, _06532_, \oc8051_golden_model_1.PC [1]);
  and (_25429_, _25428_, _25427_);
  or (_25430_, _25429_, _06013_);
  nand (_25432_, _07031_, _06013_);
  and (_25433_, _25432_, _12733_);
  and (_25434_, _25433_, _25430_);
  or (_25435_, _25205_, \oc8051_golden_model_1.PSW [7]);
  nand (_25436_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_25437_, _25436_, _12732_);
  and (_25438_, _25437_, _25435_);
  or (_25439_, _25438_, _12745_);
  or (_25440_, _25439_, _25434_);
  and (_25441_, _25440_, _25185_);
  nor (_25443_, _07446_, _07059_);
  or (_25444_, _25443_, _25441_);
  nand (_25445_, _25443_, _06034_);
  nor (_25446_, _09012_, _07059_);
  nor (_25447_, _25446_, _10989_);
  and (_25448_, _25447_, _25445_);
  and (_25449_, _25448_, _25444_);
  nor (_25450_, _25447_, _06034_);
  or (_25451_, _25450_, _11008_);
  or (_25452_, _25451_, _25449_);
  or (_25454_, _11007_, _05585_);
  and (_25455_, _25454_, _07229_);
  and (_25456_, _25455_, _25452_);
  nand (_25457_, _06437_, _06034_);
  nand (_25458_, _25457_, _12759_);
  or (_25459_, _25458_, _25456_);
  nand (_25460_, _07031_, _06008_);
  and (_25461_, _25460_, _12762_);
  or (_25462_, _06008_, _05585_);
  or (_25463_, _25462_, _07231_);
  and (_25465_, _25463_, _25461_);
  and (_25466_, _25465_, _25459_);
  or (_25467_, _25205_, _10774_);
  or (_25468_, \oc8051_golden_model_1.PSW [7], _05585_);
  and (_25469_, _25468_, _12239_);
  and (_25470_, _25469_, _25467_);
  or (_25471_, _25470_, _12771_);
  or (_25472_, _25471_, _25466_);
  and (_25473_, _25472_, _25184_);
  or (_25474_, _25473_, _12770_);
  or (_25476_, _12769_, _05585_);
  and (_25477_, _25476_, _12775_);
  and (_25478_, _25477_, _25474_);
  and (_25479_, _11111_, _06035_);
  or (_25480_, _25479_, _06543_);
  or (_25481_, _25480_, _25478_);
  or (_25482_, _09339_, _12782_);
  and (_25483_, _25482_, _25481_);
  or (_25484_, _25483_, _06011_);
  nand (_25485_, _07031_, _06011_);
  and (_25487_, _25485_, _12786_);
  and (_25488_, _25487_, _25484_);
  or (_25489_, _12970_, _06034_);
  or (_25490_, _25193_, _25133_);
  and (_25491_, _25490_, _06436_);
  and (_25492_, _25491_, _25489_);
  or (_25493_, _25492_, _12790_);
  or (_25494_, _25493_, _25488_);
  and (_25495_, _25494_, _25183_);
  or (_25496_, _25495_, _12979_);
  or (_25498_, _12978_, _05585_);
  and (_25499_, _25498_, _12981_);
  and (_25500_, _25499_, _25496_);
  and (_25501_, _10472_, _06035_);
  or (_25502_, _25501_, _06290_);
  or (_25503_, _25502_, _25500_);
  or (_25504_, _09339_, _06291_);
  and (_25505_, _25504_, _25503_);
  or (_25506_, _25505_, _05994_);
  nand (_25507_, _07031_, _05994_);
  and (_25509_, _25507_, _06435_);
  and (_25510_, _25509_, _25506_);
  or (_25511_, _25193_, _12970_);
  nand (_25512_, _12970_, _06035_);
  and (_25513_, _25512_, _25511_);
  and (_25514_, _25513_, _06434_);
  or (_25515_, _25514_, _14448_);
  or (_25516_, _25515_, _25510_);
  and (_25517_, _25516_, _25182_);
  or (_25518_, _25517_, _07245_);
  or (_25520_, _07244_, _06035_);
  and (_25521_, _25520_, _07240_);
  and (_25522_, _25521_, _25518_);
  or (_25523_, _25522_, _25181_);
  and (_25524_, _25523_, _13005_);
  nor (_25525_, _13005_, _06034_);
  or (_25526_, _25525_, _07678_);
  or (_25527_, _25526_, _25524_);
  nand (_25528_, _07678_, _07031_);
  and (_25529_, _25528_, _05933_);
  and (_25531_, _25529_, _25527_);
  and (_25532_, _25513_, _05932_);
  and (_25533_, _07482_, _10952_);
  or (_25534_, _25533_, _25532_);
  or (_25535_, _25534_, _25531_);
  nor (_25536_, _07472_, _07042_);
  and (_25537_, _25533_, _06034_);
  nor (_25538_, _25537_, _25536_);
  and (_25539_, _25538_, _25535_);
  nand (_25540_, _25536_, _06035_);
  and (_25542_, _17951_, _05766_);
  nor (_25543_, _25542_, _07261_);
  nand (_25544_, _25543_, _25540_);
  or (_25545_, _25544_, _25539_);
  or (_25546_, _25543_, _06035_);
  and (_25547_, _25546_, _06570_);
  and (_25548_, _25547_, _25545_);
  or (_25549_, _25548_, _25180_);
  and (_25550_, _25549_, _13027_);
  nor (_25551_, _13027_, _06034_);
  or (_25553_, _25551_, _25169_);
  or (_25554_, _25553_, _25550_);
  nand (_25555_, _25169_, _07031_);
  and (_25556_, _25555_, _13039_);
  and (_25557_, _25556_, _25554_);
  and (_25558_, _13035_, _06035_);
  or (_25559_, _25558_, _01324_);
  or (_25560_, _25559_, _25557_);
  or (_25561_, _01320_, \oc8051_golden_model_1.PC [1]);
  and (_25562_, _25561_, _42355_);
  and (_42984_, _25562_, _25560_);
  and (_25564_, _06566_, _06060_);
  or (_25565_, _12129_, _06074_);
  or (_25566_, _12767_, _06074_);
  or (_25567_, _12749_, _06074_);
  or (_25568_, _12244_, _06074_);
  or (_25569_, _12695_, _06074_);
  and (_25570_, _06702_, _06003_);
  and (_25571_, _25570_, _06060_);
  nand (_25572_, _07510_, _06451_);
  or (_25574_, _25304_, _06060_);
  nand (_25575_, _12254_, _06075_);
  and (_25576_, _12430_, _06060_);
  nor (_25577_, _12196_, _12194_);
  nor (_25578_, _25577_, _12197_);
  and (_25579_, _25578_, _12432_);
  or (_25580_, _25579_, _08736_);
  or (_25581_, _25580_, _25576_);
  nor (_25582_, _07858_, _06689_);
  nand (_25583_, _07143_, _06451_);
  nor (_25585_, _07143_, \oc8051_golden_model_1.PC [2]);
  nand (_25586_, _25585_, _07454_);
  and (_25587_, _25586_, _25583_);
  or (_25588_, _25587_, _06755_);
  or (_25589_, _24975_, _06074_);
  and (_25590_, _25589_, _25588_);
  or (_25591_, _25590_, _12448_);
  and (_25592_, _25591_, _07858_);
  or (_25593_, _25592_, _25582_);
  nand (_25594_, _12448_, _06075_);
  and (_25596_, _25594_, _25593_);
  or (_25597_, _25596_, _08734_);
  and (_25598_, _25597_, _25581_);
  or (_25599_, _25598_, _07159_);
  nand (_25600_, _07159_, _06075_);
  and (_25601_, _25600_, _06286_);
  and (_25602_, _25601_, _25599_);
  or (_25603_, _12326_, _12324_);
  and (_25604_, _25603_, _12327_);
  or (_25605_, _25604_, _12418_);
  or (_25607_, _12420_, _12314_);
  and (_25608_, _25607_, _06285_);
  and (_25609_, _25608_, _25605_);
  or (_25610_, _25609_, _12410_);
  or (_25611_, _25610_, _25602_);
  or (_25612_, _12409_, _06074_);
  and (_25613_, _25612_, _06282_);
  and (_25614_, _25613_, _25611_);
  and (_25615_, _06281_, _06060_);
  or (_25616_, _25615_, _07460_);
  or (_25618_, _25616_, _25614_);
  nand (_25619_, _06689_, _07460_);
  and (_25620_, _25619_, _07169_);
  and (_25621_, _25620_, _25618_);
  nand (_25622_, _06354_, _06060_);
  nand (_25623_, _25622_, _12404_);
  or (_25624_, _25623_, _25621_);
  or (_25625_, _12404_, _06074_);
  and (_25626_, _25625_, _06346_);
  and (_25627_, _25626_, _25624_);
  nand (_25628_, _06345_, _06060_);
  nand (_25629_, _25628_, _12468_);
  or (_25630_, _25629_, _25627_);
  or (_25631_, _12468_, _06074_);
  and (_25632_, _25631_, _06278_);
  and (_25633_, _25632_, _25630_);
  and (_25634_, _06277_, _06060_);
  or (_25635_, _25634_, _12475_);
  or (_25636_, _25635_, _25633_);
  nand (_25637_, _06689_, _12475_);
  and (_25640_, _25637_, _06778_);
  and (_25641_, _25640_, _25636_);
  nand (_25642_, _06276_, _06060_);
  nand (_25643_, _25642_, _12484_);
  or (_25644_, _25643_, _25641_);
  or (_25645_, _25604_, _12519_);
  or (_25646_, _25019_, _12314_);
  and (_25647_, _25646_, _25645_);
  or (_25648_, _25647_, _12484_);
  and (_25649_, _25648_, _25644_);
  or (_25651_, _25649_, _06423_);
  and (_25652_, _12400_, _12314_);
  and (_25653_, _25604_, _12398_);
  or (_25654_, _25653_, _25652_);
  or (_25655_, _25654_, _06424_);
  and (_25656_, _25655_, _25651_);
  or (_25657_, _25656_, _06347_);
  and (_25658_, _12540_, _12314_);
  and (_25659_, _25604_, _25279_);
  or (_25660_, _25659_, _14105_);
  or (_25662_, _25660_, _25658_);
  and (_25663_, _25662_, _12528_);
  and (_25664_, _25663_, _25657_);
  or (_25665_, _25604_, _12559_);
  or (_25666_, _12560_, _12314_);
  and (_25667_, _25666_, _06419_);
  and (_25668_, _25667_, _25665_);
  or (_25669_, _25668_, _12254_);
  or (_25670_, _25669_, _25664_);
  and (_25671_, _25670_, _25575_);
  or (_25673_, _25671_, _06270_);
  nand (_25674_, _06270_, _06451_);
  and (_25675_, _25674_, _05946_);
  and (_25676_, _25675_, _25673_);
  nor (_25677_, _06689_, _05946_);
  or (_25678_, _25677_, _25305_);
  or (_25679_, _25678_, _25676_);
  and (_25680_, _25679_, _25574_);
  or (_25681_, _25680_, _12589_);
  or (_25682_, _12585_, _06074_);
  and (_25684_, _25682_, _14014_);
  and (_25685_, _25684_, _25681_);
  and (_25686_, _06371_, _06060_);
  or (_25687_, _25686_, _25318_);
  or (_25688_, _25687_, _25685_);
  nand (_25689_, _06689_, _25318_);
  and (_25690_, _25689_, _14013_);
  and (_25691_, _25690_, _25688_);
  nand (_25692_, _06370_, _06060_);
  nand (_25693_, _25692_, _12595_);
  or (_25695_, _25693_, _25691_);
  or (_25696_, _12595_, _06074_);
  and (_25697_, _25696_, _25695_);
  or (_25698_, _25697_, _12600_);
  or (_25699_, _12599_, _06060_);
  and (_25700_, _25699_, _05940_);
  and (_25701_, _25700_, _25698_);
  nor (_25702_, _06075_, _05940_);
  or (_25703_, _25702_, _06266_);
  or (_25704_, _25703_, _25701_);
  nand (_25706_, _06266_, _06451_);
  and (_25707_, _25706_, _25704_);
  or (_25708_, _25707_, _05974_);
  nand (_25709_, _06689_, _05974_);
  and (_25710_, _25709_, _06396_);
  and (_25711_, _25710_, _25708_);
  and (_25712_, _12314_, _06395_);
  or (_25713_, _25712_, _07510_);
  or (_25714_, _25713_, _25711_);
  and (_25715_, _25714_, _25572_);
  nor (_25717_, _07449_, _05983_);
  or (_25718_, _25717_, _25715_);
  nand (_25719_, _25717_, _06451_);
  and (_25720_, _25719_, _06251_);
  and (_25721_, _25720_, _25718_);
  nand (_25722_, _12314_, _05972_);
  nand (_25723_, _25722_, _12252_);
  or (_25724_, _25723_, _25721_);
  or (_25725_, _12252_, _06074_);
  and (_25726_, _25725_, _06854_);
  and (_25728_, _25726_, _25724_);
  and (_25729_, _06330_, _06060_);
  or (_25730_, _25729_, _05997_);
  or (_25731_, _25730_, _25728_);
  nand (_25732_, _06689_, _05997_);
  and (_25733_, _25732_, _25731_);
  or (_25734_, _25733_, _12630_);
  nor (_25735_, _25578_, _12631_);
  nor (_25736_, _25735_, _25570_);
  and (_25737_, _25736_, _25734_);
  nor (_25739_, _25737_, _25571_);
  nor (_25740_, _10954_, _07205_);
  nor (_25741_, _25740_, _25739_);
  and (_25742_, _25740_, _06060_);
  or (_25743_, _25742_, _09013_);
  or (_25744_, _25743_, _25741_);
  nand (_25745_, _09013_, _06451_);
  and (_25746_, _25745_, _06216_);
  and (_25747_, _25746_, _25744_);
  and (_25748_, _12314_, _06215_);
  or (_25750_, _25748_, _10891_);
  or (_25751_, _25750_, _25747_);
  nand (_25752_, _10891_, _06451_);
  and (_25753_, _25752_, _25751_);
  or (_25754_, _25753_, _12644_);
  or (_25755_, _25380_, _06070_);
  and (_25756_, _25755_, _06860_);
  and (_25757_, _25756_, _25754_);
  and (_25758_, _06329_, _06060_);
  or (_25759_, _25758_, _06004_);
  or (_25761_, _25759_, _25757_);
  nand (_25762_, _06689_, _06004_);
  and (_25763_, _25762_, _12685_);
  and (_25764_, _25763_, _25761_);
  or (_25765_, _25578_, _11327_);
  nand (_25766_, _11327_, _06451_);
  and (_25767_, _25766_, _12247_);
  and (_25768_, _25767_, _25765_);
  or (_25769_, _25768_, _12697_);
  or (_25770_, _25769_, _25764_);
  and (_25772_, _25770_, _25569_);
  or (_25773_, _25772_, _12700_);
  or (_25774_, _12699_, _06060_);
  and (_25775_, _25774_, _09025_);
  and (_25776_, _25775_, _25773_);
  and (_25777_, _12314_, _06398_);
  or (_25778_, _25777_, _06524_);
  or (_25779_, _25778_, _25776_);
  nand (_25780_, _06524_, _06451_);
  and (_25781_, _25780_, _25779_);
  or (_25783_, _25781_, _06001_);
  nand (_25784_, _06689_, _06001_);
  and (_25785_, _25784_, _12712_);
  and (_25786_, _25785_, _25783_);
  or (_25787_, _25578_, _12248_);
  or (_25788_, _11327_, _06060_);
  and (_25789_, _25788_, _12711_);
  and (_25790_, _25789_, _25787_);
  or (_25791_, _25790_, _12720_);
  or (_25792_, _25791_, _25786_);
  and (_25794_, _25792_, _25568_);
  or (_25795_, _25794_, _10970_);
  or (_25796_, _10969_, _06060_);
  and (_25797_, _25796_, _07219_);
  and (_25798_, _25797_, _25795_);
  and (_25799_, _12314_, _06426_);
  or (_25800_, _25799_, _06532_);
  or (_25801_, _25800_, _25798_);
  nand (_25802_, _06532_, _06451_);
  and (_25803_, _25802_, _25801_);
  or (_25805_, _25803_, _06013_);
  nand (_25806_, _06689_, _06013_);
  and (_25807_, _25806_, _12733_);
  and (_25808_, _25807_, _25805_);
  or (_25809_, _25578_, \oc8051_golden_model_1.PSW [7]);
  or (_25810_, _06060_, _10774_);
  and (_25811_, _25810_, _12732_);
  and (_25812_, _25811_, _25809_);
  or (_25813_, _25812_, _12751_);
  or (_25814_, _25813_, _25808_);
  and (_25816_, _25814_, _25567_);
  or (_25817_, _25816_, _11008_);
  or (_25818_, _11007_, _06060_);
  and (_25819_, _25818_, _07229_);
  and (_25820_, _25819_, _25817_);
  and (_25821_, _12314_, _06437_);
  or (_25822_, _25821_, _06535_);
  or (_25823_, _25822_, _25820_);
  nand (_25824_, _06535_, _06451_);
  and (_25825_, _25824_, _25823_);
  or (_25827_, _25825_, _06008_);
  nand (_25828_, _06689_, _06008_);
  and (_25829_, _25828_, _12762_);
  and (_25830_, _25829_, _25827_);
  or (_25831_, _25578_, _10774_);
  or (_25832_, _06060_, \oc8051_golden_model_1.PSW [7]);
  and (_25833_, _25832_, _12239_);
  and (_25834_, _25833_, _25831_);
  or (_25835_, _25834_, _12771_);
  or (_25836_, _25835_, _25830_);
  and (_25838_, _25836_, _25566_);
  or (_25839_, _25838_, _12770_);
  or (_25840_, _12769_, _06060_);
  and (_25841_, _25840_, _12775_);
  and (_25842_, _25841_, _25839_);
  and (_25843_, _11111_, _06074_);
  or (_25844_, _25843_, _06543_);
  or (_25845_, _25844_, _25842_);
  or (_25846_, _09293_, _12782_);
  and (_25847_, _25846_, _25845_);
  or (_25849_, _25847_, _06011_);
  nand (_25850_, _06689_, _06011_);
  and (_25851_, _25850_, _12786_);
  and (_25852_, _25851_, _25849_);
  or (_25853_, _25604_, _25133_);
  or (_25854_, _12314_, _12970_);
  and (_25855_, _25854_, _06436_);
  and (_25856_, _25855_, _25853_);
  or (_25857_, _25856_, _12790_);
  or (_25858_, _25857_, _25852_);
  and (_25860_, _25858_, _25565_);
  or (_25861_, _25860_, _12979_);
  or (_25862_, _12978_, _06060_);
  and (_25863_, _25862_, _12981_);
  and (_25864_, _25863_, _25861_);
  and (_25865_, _10472_, _06074_);
  or (_25866_, _25865_, _06290_);
  or (_25867_, _25866_, _25864_);
  or (_25868_, _09293_, _06291_);
  and (_25869_, _25868_, _25867_);
  or (_25871_, _25869_, _05994_);
  nand (_25872_, _06689_, _05994_);
  and (_25873_, _25872_, _06435_);
  and (_25874_, _25873_, _25871_);
  or (_25875_, _25604_, _12970_);
  or (_25876_, _12314_, _25133_);
  and (_25877_, _25876_, _25875_);
  and (_25878_, _25877_, _06434_);
  or (_25879_, _25878_, _12999_);
  or (_25880_, _25879_, _25874_);
  or (_25882_, _12998_, _06074_);
  and (_25883_, _25882_, _07240_);
  and (_25884_, _25883_, _25880_);
  nand (_25885_, _06559_, _06060_);
  nand (_25886_, _25885_, _13005_);
  or (_25887_, _25886_, _25884_);
  or (_25888_, _13005_, _06074_);
  and (_25889_, _25888_, _25887_);
  or (_25890_, _25889_, _07678_);
  nand (_25891_, _07678_, _06689_);
  and (_25893_, _25891_, _05933_);
  and (_25894_, _25893_, _25890_);
  and (_25895_, _25877_, _05932_);
  or (_25896_, _25895_, _13020_);
  or (_25897_, _25896_, _25894_);
  or (_25898_, _13019_, _06074_);
  and (_25899_, _25898_, _06570_);
  and (_25900_, _25899_, _25897_);
  or (_25901_, _25900_, _25564_);
  and (_25902_, _25901_, _13027_);
  nor (_25904_, _13027_, _06075_);
  or (_25905_, _25904_, _25169_);
  or (_25906_, _25905_, _25902_);
  nand (_25907_, _25169_, _06689_);
  and (_25908_, _25907_, _13039_);
  and (_25909_, _25908_, _25906_);
  and (_25910_, _13035_, _06074_);
  or (_25911_, _25910_, _01324_);
  or (_25912_, _25911_, _25909_);
  or (_25913_, _01320_, \oc8051_golden_model_1.PC [2]);
  and (_25915_, _25913_, _42355_);
  and (_42985_, _25915_, _25912_);
  and (_25916_, _06566_, _06095_);
  and (_25917_, _06559_, _06095_);
  or (_25918_, _09247_, _06291_);
  or (_25919_, _12129_, _06458_);
  or (_25920_, _12767_, _06458_);
  or (_25921_, _12749_, _06458_);
  or (_25922_, _12244_, _06458_);
  or (_25923_, _12695_, _06458_);
  or (_25925_, _09015_, _06095_);
  nand (_25926_, _06266_, _06456_);
  or (_25927_, _25304_, _06095_);
  nand (_25928_, _12254_, _06100_);
  nor (_25929_, _07858_, _06517_);
  nand (_25930_, _07143_, _06456_);
  and (_25931_, _25930_, _06756_);
  and (_25932_, _07454_, \oc8051_golden_model_1.PC [3]);
  or (_25933_, _25932_, _07143_);
  and (_25934_, _25933_, _25931_);
  nor (_25936_, _24975_, _06100_);
  or (_25937_, _25936_, _12448_);
  or (_25938_, _25937_, _25934_);
  and (_25939_, _25938_, _07858_);
  or (_25940_, _25939_, _25929_);
  nand (_25941_, _12448_, _06100_);
  and (_25942_, _25941_, _25940_);
  or (_25943_, _25942_, _08734_);
  and (_25944_, _12430_, _06095_);
  or (_25945_, _12186_, _12185_);
  nand (_25947_, _25945_, _12198_);
  or (_25948_, _25945_, _12198_);
  and (_25949_, _25948_, _25947_);
  and (_25950_, _25949_, _12432_);
  or (_25951_, _25950_, _08736_);
  or (_25952_, _25951_, _25944_);
  and (_25953_, _25952_, _25943_);
  or (_25954_, _25953_, _07159_);
  nand (_25955_, _07159_, _06100_);
  and (_25956_, _25955_, _06286_);
  and (_25957_, _25956_, _25954_);
  and (_25958_, _12418_, _12310_);
  or (_25959_, _12312_, _12311_);
  nand (_25960_, _25959_, _12328_);
  or (_25961_, _25959_, _12328_);
  and (_25962_, _25961_, _25960_);
  and (_25963_, _25962_, _12420_);
  or (_25964_, _25963_, _25958_);
  and (_25965_, _25964_, _06285_);
  or (_25966_, _25965_, _12410_);
  or (_25969_, _25966_, _25957_);
  or (_25970_, _12409_, _06458_);
  and (_25971_, _25970_, _06282_);
  and (_25972_, _25971_, _25969_);
  and (_25973_, _06281_, _06095_);
  or (_25974_, _25973_, _07460_);
  or (_25975_, _25974_, _25972_);
  nand (_25976_, _06517_, _07460_);
  and (_25977_, _25976_, _07169_);
  and (_25978_, _25977_, _25975_);
  nand (_25980_, _06354_, _06095_);
  nand (_25981_, _25980_, _12404_);
  or (_25982_, _25981_, _25978_);
  or (_25983_, _12404_, _06458_);
  and (_25984_, _25983_, _06346_);
  and (_25985_, _25984_, _25982_);
  nand (_25986_, _06345_, _06095_);
  nand (_25987_, _25986_, _12468_);
  or (_25988_, _25987_, _25985_);
  or (_25989_, _12468_, _06458_);
  and (_25991_, _25989_, _06278_);
  and (_25992_, _25991_, _25988_);
  and (_25993_, _06277_, _06095_);
  or (_25994_, _25993_, _12475_);
  or (_25995_, _25994_, _25992_);
  nand (_25996_, _06517_, _12475_);
  and (_25997_, _25996_, _06778_);
  and (_25998_, _25997_, _25995_);
  nand (_25999_, _06276_, _06095_);
  nand (_26000_, _25999_, _12484_);
  or (_26002_, _26000_, _25998_);
  and (_26003_, _12519_, _12310_);
  and (_26004_, _25962_, _25019_);
  or (_26005_, _26004_, _26003_);
  or (_26006_, _26005_, _12484_);
  and (_26007_, _26006_, _26002_);
  or (_26008_, _26007_, _06423_);
  and (_26009_, _12400_, _12310_);
  and (_26010_, _25962_, _12398_);
  or (_26011_, _26010_, _26009_);
  or (_26013_, _26011_, _06424_);
  and (_26014_, _26013_, _26008_);
  or (_26015_, _26014_, _06347_);
  and (_26016_, _25962_, _25279_);
  and (_26017_, _12540_, _12310_);
  or (_26018_, _26017_, _14105_);
  or (_26019_, _26018_, _26016_);
  and (_26020_, _26019_, _12528_);
  and (_26021_, _26020_, _26015_);
  or (_26022_, _25962_, _12559_);
  or (_26024_, _12560_, _12310_);
  and (_26025_, _26024_, _06419_);
  and (_26026_, _26025_, _26022_);
  or (_26027_, _26026_, _12254_);
  or (_26028_, _26027_, _26021_);
  and (_26029_, _26028_, _25928_);
  or (_26030_, _26029_, _06270_);
  nand (_26031_, _06270_, _06456_);
  and (_26032_, _26031_, _05946_);
  and (_26033_, _26032_, _26030_);
  nor (_26035_, _06517_, _05946_);
  or (_26036_, _26035_, _25305_);
  or (_26037_, _26036_, _26033_);
  and (_26038_, _26037_, _25927_);
  or (_26039_, _26038_, _12589_);
  or (_26040_, _12585_, _06458_);
  and (_26041_, _26040_, _14014_);
  and (_26042_, _26041_, _26039_);
  and (_26043_, _06371_, _06095_);
  or (_26044_, _26043_, _25318_);
  or (_26046_, _26044_, _26042_);
  nand (_26047_, _06517_, _25318_);
  and (_26048_, _26047_, _14013_);
  and (_26049_, _26048_, _26046_);
  nand (_26050_, _06370_, _06095_);
  nand (_26051_, _26050_, _12595_);
  or (_26052_, _26051_, _26049_);
  or (_26053_, _12595_, _06458_);
  and (_26054_, _26053_, _26052_);
  or (_26055_, _26054_, _12600_);
  or (_26057_, _12599_, _06095_);
  and (_26058_, _26057_, _05940_);
  and (_26059_, _26058_, _26055_);
  nor (_26060_, _05940_, _06100_);
  or (_26061_, _26060_, _06266_);
  or (_26062_, _26061_, _26059_);
  and (_26063_, _26062_, _25926_);
  or (_26064_, _26063_, _05974_);
  nand (_26065_, _06517_, _05974_);
  and (_26066_, _26065_, _06396_);
  and (_26068_, _26066_, _26064_);
  nand (_26069_, _12310_, _06395_);
  nand (_26070_, _26069_, _06261_);
  or (_26071_, _26070_, _26068_);
  or (_26072_, _06261_, _06095_);
  and (_26073_, _26072_, _06251_);
  and (_26074_, _26073_, _26071_);
  nand (_26075_, _12310_, _05972_);
  nand (_26076_, _26075_, _12252_);
  or (_26077_, _26076_, _26074_);
  or (_26079_, _12252_, _06458_);
  and (_26080_, _26079_, _06854_);
  and (_26081_, _26080_, _26077_);
  and (_26082_, _06330_, _06095_);
  or (_26083_, _26082_, _05997_);
  or (_26084_, _26083_, _26081_);
  nand (_26085_, _06517_, _05997_);
  and (_26086_, _26085_, _12631_);
  and (_26087_, _26086_, _26084_);
  and (_26088_, _25949_, _12630_);
  or (_26090_, _26088_, _09016_);
  or (_26091_, _26090_, _26087_);
  and (_26092_, _26091_, _25925_);
  or (_26093_, _26092_, _06215_);
  or (_26094_, _12310_, _06216_);
  and (_26095_, _26094_, _10892_);
  and (_26096_, _26095_, _26093_);
  and (_26097_, _10891_, _06095_);
  or (_26098_, _26097_, _12644_);
  or (_26099_, _26098_, _26096_);
  or (_26101_, _25380_, _06115_);
  and (_26102_, _26101_, _06860_);
  and (_26103_, _26102_, _26099_);
  and (_26104_, _06329_, _06095_);
  or (_26105_, _26104_, _06004_);
  or (_26106_, _26105_, _26103_);
  nand (_26107_, _06517_, _06004_);
  and (_26108_, _26107_, _12685_);
  and (_26109_, _26108_, _26106_);
  or (_26110_, _25949_, _11327_);
  nand (_26112_, _11327_, _06456_);
  and (_26113_, _26112_, _12247_);
  and (_26114_, _26113_, _26110_);
  or (_26115_, _26114_, _12697_);
  or (_26116_, _26115_, _26109_);
  and (_26117_, _26116_, _25923_);
  or (_26118_, _26117_, _12700_);
  or (_26119_, _12699_, _06095_);
  and (_26120_, _26119_, _09025_);
  and (_26121_, _26120_, _26118_);
  and (_26123_, _12310_, _06398_);
  or (_26124_, _26123_, _06524_);
  or (_26125_, _26124_, _26121_);
  nand (_26126_, _06524_, _06456_);
  and (_26127_, _26126_, _26125_);
  or (_26128_, _26127_, _06001_);
  nand (_26129_, _06517_, _06001_);
  and (_26130_, _26129_, _12712_);
  and (_26131_, _26130_, _26128_);
  or (_26132_, _25949_, _12248_);
  or (_26134_, _11327_, _06095_);
  and (_26135_, _26134_, _12711_);
  and (_26136_, _26135_, _26132_);
  or (_26137_, _26136_, _12720_);
  or (_26138_, _26137_, _26131_);
  and (_26139_, _26138_, _25922_);
  or (_26140_, _26139_, _10970_);
  or (_26141_, _10969_, _06095_);
  and (_26142_, _26141_, _07219_);
  and (_26143_, _26142_, _26140_);
  and (_26145_, _12310_, _06426_);
  or (_26146_, _26145_, _06532_);
  or (_26147_, _26146_, _26143_);
  nand (_26148_, _06532_, _06456_);
  and (_26149_, _26148_, _26147_);
  or (_26150_, _26149_, _06013_);
  nand (_26151_, _06517_, _06013_);
  and (_26152_, _26151_, _12733_);
  and (_26153_, _26152_, _26150_);
  or (_26154_, _25949_, \oc8051_golden_model_1.PSW [7]);
  or (_26156_, _06095_, _10774_);
  and (_26157_, _26156_, _12732_);
  and (_26158_, _26157_, _26154_);
  or (_26159_, _26158_, _12751_);
  or (_26160_, _26159_, _26153_);
  and (_26161_, _26160_, _25921_);
  or (_26162_, _26161_, _11008_);
  or (_26163_, _11007_, _06095_);
  and (_26164_, _26163_, _07229_);
  and (_26165_, _26164_, _26162_);
  and (_26167_, _12310_, _06437_);
  or (_26168_, _26167_, _06535_);
  or (_26169_, _26168_, _26165_);
  nand (_26170_, _06535_, _06456_);
  and (_26171_, _26170_, _26169_);
  or (_26172_, _26171_, _06008_);
  nand (_26173_, _06517_, _06008_);
  and (_26174_, _26173_, _12762_);
  and (_26175_, _26174_, _26172_);
  or (_26176_, _25949_, _10774_);
  or (_26178_, _06095_, \oc8051_golden_model_1.PSW [7]);
  and (_26179_, _26178_, _12239_);
  and (_26180_, _26179_, _26176_);
  or (_26181_, _26180_, _12771_);
  or (_26182_, _26181_, _26175_);
  and (_26183_, _26182_, _25920_);
  or (_26184_, _26183_, _12770_);
  or (_26185_, _12769_, _06095_);
  and (_26186_, _26185_, _12775_);
  and (_26187_, _26186_, _26184_);
  and (_26189_, _11111_, _06458_);
  or (_26190_, _26189_, _06543_);
  or (_26191_, _26190_, _26187_);
  or (_26192_, _09247_, _12782_);
  and (_26193_, _26192_, _26191_);
  or (_26194_, _26193_, _06011_);
  nand (_26195_, _06517_, _06011_);
  and (_26196_, _26195_, _12786_);
  and (_26197_, _26196_, _26194_);
  or (_26198_, _25962_, _25133_);
  or (_26200_, _12310_, _12970_);
  and (_26201_, _26200_, _06436_);
  and (_26202_, _26201_, _26198_);
  or (_26203_, _26202_, _12790_);
  or (_26204_, _26203_, _26197_);
  and (_26205_, _26204_, _25919_);
  or (_26206_, _26205_, _12979_);
  or (_26207_, _12978_, _06095_);
  and (_26208_, _26207_, _12981_);
  and (_26209_, _26208_, _26206_);
  and (_26211_, _10472_, _06458_);
  or (_26212_, _26211_, _06290_);
  or (_26213_, _26212_, _26209_);
  and (_26214_, _26213_, _25918_);
  or (_26215_, _26214_, _05994_);
  nand (_26216_, _06517_, _05994_);
  and (_26217_, _26216_, _06435_);
  and (_26218_, _26217_, _26215_);
  or (_26219_, _25962_, _12970_);
  or (_26220_, _12310_, _25133_);
  and (_26222_, _26220_, _26219_);
  and (_26223_, _26222_, _06434_);
  or (_26224_, _26223_, _12999_);
  or (_26225_, _26224_, _26218_);
  or (_26226_, _12998_, _06458_);
  and (_26227_, _26226_, _07240_);
  and (_26228_, _26227_, _26225_);
  or (_26229_, _26228_, _25917_);
  and (_26230_, _26229_, _13005_);
  nor (_26231_, _13005_, _06100_);
  or (_26233_, _26231_, _07678_);
  or (_26234_, _26233_, _26230_);
  nand (_26235_, _07678_, _06517_);
  and (_26236_, _26235_, _05933_);
  and (_26237_, _26236_, _26234_);
  and (_26238_, _26222_, _05932_);
  or (_26239_, _26238_, _13020_);
  or (_26240_, _26239_, _26237_);
  or (_26241_, _13019_, _06458_);
  and (_26242_, _26241_, _06570_);
  and (_26244_, _26242_, _26240_);
  or (_26245_, _26244_, _25916_);
  and (_26246_, _26245_, _13027_);
  nor (_26247_, _13027_, _06100_);
  or (_26248_, _26247_, _25169_);
  or (_26249_, _26248_, _26246_);
  nand (_26250_, _25169_, _06517_);
  and (_26251_, _26250_, _13039_);
  and (_26252_, _26251_, _26249_);
  and (_26253_, _13035_, _06458_);
  or (_26255_, _26253_, _01324_);
  or (_26256_, _26255_, _26252_);
  or (_26257_, _01320_, \oc8051_golden_model_1.PC [3]);
  and (_26258_, _26257_, _42355_);
  and (_42987_, _26258_, _26256_);
  not (_26259_, \oc8051_golden_model_1.PC [4]);
  nor (_26260_, _01320_, _26259_);
  nand (_26261_, _25169_, _08879_);
  nand (_26262_, _08879_, _07678_);
  or (_26263_, _12202_, _12200_);
  and (_26265_, _26263_, _12203_);
  or (_26266_, _26265_, _11327_);
  or (_26267_, _12183_, _12248_);
  and (_26268_, _26267_, _12247_);
  and (_26269_, _26268_, _26266_);
  or (_26270_, _12183_, _09015_);
  or (_26271_, _12183_, _06267_);
  or (_26272_, _25304_, _12183_);
  nor (_26273_, _05602_, _26259_);
  and (_26274_, _05602_, _26259_);
  nor (_26276_, _26274_, _26273_);
  not (_26277_, _26276_);
  nand (_26278_, _26277_, _12254_);
  and (_26279_, _12400_, _12307_);
  or (_26280_, _12332_, _12330_);
  and (_26281_, _26280_, _12333_);
  and (_26282_, _26281_, _12398_);
  or (_26283_, _26282_, _26279_);
  and (_26284_, _26283_, _06423_);
  or (_26285_, _12183_, _06278_);
  or (_26287_, _26276_, _12404_);
  not (_26288_, _12404_);
  or (_26289_, _26281_, _12418_);
  or (_26290_, _12420_, _12307_);
  and (_26291_, _26290_, _06285_);
  and (_26292_, _26291_, _26289_);
  and (_26293_, _12430_, _12183_);
  and (_26294_, _26265_, _12432_);
  or (_26295_, _26294_, _26293_);
  or (_26296_, _26295_, _08736_);
  nand (_26298_, _08879_, _07152_);
  or (_26299_, _12183_, _07144_);
  and (_26300_, _26299_, _06756_);
  and (_26301_, _07454_, \oc8051_golden_model_1.PC [4]);
  or (_26302_, _26301_, _07143_);
  and (_26303_, _26302_, _26300_);
  nor (_26304_, _26277_, _24975_);
  or (_26305_, _26304_, _07152_);
  or (_26306_, _26305_, _26303_);
  and (_26307_, _26306_, _12453_);
  and (_26309_, _26307_, _26298_);
  and (_26310_, _26276_, _12448_);
  or (_26311_, _26310_, _08734_);
  or (_26312_, _26311_, _26309_);
  and (_26313_, _26312_, _12457_);
  and (_26314_, _26313_, _26296_);
  or (_26315_, _26314_, _26292_);
  and (_26316_, _26315_, _12409_);
  nor (_26317_, _26277_, _12411_);
  or (_26318_, _26317_, _06281_);
  or (_26320_, _26318_, _26316_);
  or (_26321_, _12183_, _06282_);
  and (_26322_, _26321_, _05949_);
  and (_26323_, _26322_, _26320_);
  nor (_26324_, _08879_, _05949_);
  or (_26325_, _26324_, _06354_);
  or (_26326_, _26325_, _26323_);
  or (_26327_, _12183_, _07169_);
  and (_26328_, _26327_, _26326_);
  or (_26329_, _26328_, _26288_);
  and (_26331_, _26329_, _26287_);
  or (_26332_, _26331_, _06345_);
  or (_26333_, _12183_, _06346_);
  and (_26334_, _26333_, _12468_);
  and (_26335_, _26334_, _26332_);
  nor (_26336_, _26277_, _12468_);
  or (_26337_, _26336_, _06277_);
  or (_26338_, _26337_, _26335_);
  and (_26339_, _26338_, _26285_);
  or (_26340_, _26339_, _12475_);
  nand (_26342_, _08879_, _12475_);
  and (_26343_, _26342_, _06778_);
  and (_26344_, _26343_, _26340_);
  nand (_26345_, _12183_, _06276_);
  nand (_26346_, _26345_, _12484_);
  or (_26347_, _26346_, _26344_);
  and (_26348_, _26281_, _25019_);
  and (_26349_, _12519_, _12307_);
  or (_26350_, _26349_, _12484_);
  or (_26351_, _26350_, _26348_);
  and (_26353_, _26351_, _06424_);
  and (_26354_, _26353_, _26347_);
  or (_26355_, _26354_, _26284_);
  and (_26356_, _26355_, _06420_);
  or (_26357_, _25279_, _12307_);
  or (_26358_, _26281_, _12540_);
  and (_26359_, _26358_, _06347_);
  and (_26360_, _26359_, _26357_);
  or (_26361_, _26281_, _12559_);
  or (_26362_, _12560_, _12307_);
  and (_26364_, _26362_, _06419_);
  and (_26365_, _26364_, _26361_);
  or (_26366_, _26365_, _12254_);
  or (_26367_, _26366_, _26360_);
  or (_26368_, _26367_, _26356_);
  and (_26369_, _26368_, _26278_);
  or (_26370_, _26369_, _06270_);
  or (_26371_, _12183_, _06271_);
  and (_26372_, _26371_, _05946_);
  and (_26373_, _26372_, _26370_);
  nor (_26375_, _08879_, _05946_);
  or (_26376_, _26375_, _25305_);
  or (_26377_, _26376_, _26373_);
  and (_26378_, _26377_, _26272_);
  or (_26379_, _26378_, _12589_);
  or (_26380_, _26276_, _12585_);
  and (_26381_, _26380_, _14014_);
  and (_26382_, _26381_, _26379_);
  and (_26383_, _12183_, _06371_);
  or (_26384_, _26383_, _25318_);
  or (_26386_, _26384_, _26382_);
  nand (_26387_, _08879_, _25318_);
  and (_26388_, _26387_, _14013_);
  and (_26389_, _26388_, _26386_);
  and (_26390_, _12183_, _06370_);
  or (_26391_, _26390_, _26389_);
  and (_26392_, _26391_, _12595_);
  nor (_26393_, _26277_, _12595_);
  or (_26394_, _26393_, _12600_);
  or (_26395_, _26394_, _26392_);
  or (_26397_, _12183_, _12599_);
  and (_26398_, _26397_, _05940_);
  and (_26399_, _26398_, _26395_);
  nor (_26400_, _26277_, _05940_);
  or (_26401_, _26400_, _06266_);
  or (_26402_, _26401_, _26399_);
  and (_26403_, _26402_, _26271_);
  or (_26404_, _26403_, _05974_);
  nand (_26405_, _08879_, _05974_);
  and (_26406_, _26405_, _06396_);
  and (_26408_, _26406_, _26404_);
  nand (_26409_, _12307_, _06395_);
  nand (_26410_, _26409_, _06261_);
  or (_26411_, _26410_, _26408_);
  or (_26412_, _12183_, _06261_);
  and (_26413_, _26412_, _06251_);
  and (_26414_, _26413_, _26411_);
  nand (_26415_, _12307_, _05972_);
  nand (_26416_, _26415_, _12252_);
  or (_26417_, _26416_, _26414_);
  or (_26419_, _26276_, _12252_);
  and (_26420_, _26419_, _06854_);
  and (_26421_, _26420_, _26417_);
  nor (_26422_, _12183_, _05997_);
  nor (_26423_, _26422_, _12624_);
  or (_26424_, _26423_, _26421_);
  nand (_26425_, _08879_, _05997_);
  and (_26426_, _26425_, _12631_);
  and (_26427_, _26426_, _26424_);
  and (_26428_, _26265_, _12630_);
  or (_26430_, _26428_, _09016_);
  or (_26431_, _26430_, _26427_);
  and (_26432_, _26431_, _26270_);
  or (_26433_, _26432_, _06215_);
  or (_26434_, _12307_, _06216_);
  and (_26435_, _26434_, _10892_);
  and (_26436_, _26435_, _26433_);
  and (_26437_, _12183_, _10891_);
  or (_26438_, _26437_, _12644_);
  or (_26439_, _26438_, _26436_);
  or (_26440_, _12659_, _12657_);
  nand (_26441_, _26440_, _12660_);
  nand (_26442_, _26441_, _12644_);
  and (_26443_, _26442_, _06860_);
  and (_26444_, _26443_, _26439_);
  and (_26445_, _12183_, _06329_);
  or (_26446_, _26445_, _06004_);
  or (_26447_, _26446_, _26444_);
  nand (_26448_, _08879_, _06004_);
  and (_26449_, _26448_, _12685_);
  and (_26452_, _26449_, _26447_);
  or (_26453_, _26452_, _26269_);
  and (_26454_, _26453_, _12695_);
  nor (_26455_, _26277_, _12695_);
  or (_26456_, _26455_, _12700_);
  or (_26457_, _26456_, _26454_);
  or (_26458_, _12699_, _12183_);
  and (_26459_, _26458_, _09025_);
  and (_26460_, _26459_, _26457_);
  and (_26461_, _12307_, _06398_);
  or (_26463_, _26461_, _06524_);
  or (_26464_, _26463_, _26460_);
  or (_26465_, _12183_, _09030_);
  and (_26466_, _26465_, _26464_);
  or (_26467_, _26466_, _06001_);
  nand (_26468_, _08879_, _06001_);
  and (_26469_, _26468_, _12712_);
  and (_26470_, _26469_, _26467_);
  or (_26471_, _26265_, _12248_);
  or (_26472_, _12183_, _11327_);
  and (_26474_, _26472_, _12711_);
  and (_26475_, _26474_, _26471_);
  or (_26476_, _26475_, _26470_);
  and (_26477_, _26476_, _12244_);
  nor (_26478_, _26277_, _12244_);
  or (_26479_, _26478_, _10970_);
  or (_26480_, _26479_, _26477_);
  or (_26481_, _12183_, _10969_);
  and (_26482_, _26481_, _07219_);
  and (_26483_, _26482_, _26480_);
  and (_26484_, _12307_, _06426_);
  or (_26485_, _26484_, _06532_);
  or (_26486_, _26485_, _26483_);
  or (_26487_, _12183_, _07217_);
  and (_26488_, _26487_, _26486_);
  or (_26489_, _26488_, _06013_);
  nand (_26490_, _08879_, _06013_);
  and (_26491_, _26490_, _12733_);
  and (_26492_, _26491_, _26489_);
  or (_26493_, _26265_, \oc8051_golden_model_1.PSW [7]);
  or (_26495_, _12183_, _10774_);
  and (_26496_, _26495_, _12732_);
  and (_26497_, _26496_, _26493_);
  or (_26498_, _26497_, _26492_);
  and (_26499_, _26498_, _12749_);
  nor (_26500_, _26277_, _12749_);
  or (_26501_, _26500_, _11008_);
  or (_26502_, _26501_, _26499_);
  or (_26503_, _12183_, _11007_);
  and (_26504_, _26503_, _07229_);
  and (_26506_, _26504_, _26502_);
  and (_26507_, _12307_, _06437_);
  or (_26508_, _26507_, _06535_);
  or (_26509_, _26508_, _26506_);
  or (_26510_, _12183_, _07231_);
  and (_26511_, _26510_, _26509_);
  or (_26512_, _26511_, _06008_);
  nand (_26513_, _08879_, _06008_);
  and (_26514_, _26513_, _12762_);
  and (_26515_, _26514_, _26512_);
  or (_26516_, _26265_, _10774_);
  or (_26517_, _12183_, \oc8051_golden_model_1.PSW [7]);
  and (_26518_, _26517_, _12239_);
  and (_26519_, _26518_, _26516_);
  or (_26520_, _26519_, _26515_);
  and (_26521_, _26520_, _12767_);
  nor (_26522_, _26277_, _12767_);
  or (_26523_, _26522_, _12770_);
  or (_26524_, _26523_, _26521_);
  or (_26525_, _12183_, _12769_);
  and (_26526_, _26525_, _12775_);
  and (_26527_, _26526_, _26524_);
  and (_26528_, _26276_, _11111_);
  or (_26529_, _26528_, _06543_);
  or (_26530_, _26529_, _26527_);
  or (_26531_, _09437_, _12782_);
  and (_26532_, _26531_, _26530_);
  or (_26533_, _26532_, _06011_);
  nand (_26534_, _08879_, _06011_);
  and (_26535_, _26534_, _12786_);
  and (_26536_, _26535_, _26533_);
  and (_26537_, _12307_, _25133_);
  and (_26538_, _26281_, _12970_);
  or (_26539_, _26538_, _26537_);
  and (_26540_, _26539_, _06436_);
  or (_26541_, _26540_, _26536_);
  and (_26542_, _26541_, _12129_);
  nor (_26543_, _26277_, _12129_);
  or (_26544_, _26543_, _12979_);
  or (_26545_, _26544_, _26542_);
  or (_26546_, _12978_, _12183_);
  and (_26547_, _26546_, _12981_);
  and (_26548_, _26547_, _26545_);
  and (_26549_, _26276_, _10472_);
  or (_26550_, _26549_, _06290_);
  or (_26551_, _26550_, _26548_);
  or (_26552_, _09437_, _06291_);
  and (_26553_, _26552_, _25143_);
  and (_26554_, _26553_, _26551_);
  nor (_26555_, _08879_, _25143_);
  or (_26556_, _26555_, _06434_);
  or (_26557_, _26556_, _26554_);
  or (_26558_, _12307_, _25133_);
  or (_26559_, _26281_, _12970_);
  and (_26560_, _26559_, _26558_);
  or (_26561_, _26560_, _06435_);
  and (_26562_, _26561_, _12998_);
  and (_26563_, _26562_, _26557_);
  nor (_26564_, _26277_, _12998_);
  or (_26565_, _26564_, _06559_);
  or (_26567_, _26565_, _26563_);
  or (_26568_, _12183_, _07240_);
  and (_26569_, _26568_, _13005_);
  and (_26570_, _26569_, _26567_);
  nor (_26571_, _26277_, _13005_);
  or (_26572_, _26571_, _07678_);
  or (_26573_, _26572_, _26570_);
  and (_26574_, _26573_, _26262_);
  or (_26575_, _26574_, _05932_);
  or (_26576_, _26560_, _05933_);
  and (_26578_, _26576_, _13019_);
  and (_26579_, _26578_, _26575_);
  nor (_26580_, _26277_, _13019_);
  or (_26581_, _26580_, _06566_);
  or (_26582_, _26581_, _26579_);
  or (_26583_, _12183_, _06570_);
  and (_26584_, _26583_, _13027_);
  and (_26585_, _26584_, _26582_);
  nor (_26586_, _26277_, _13027_);
  or (_26587_, _26586_, _25169_);
  or (_26588_, _26587_, _26585_);
  and (_26589_, _26588_, _26261_);
  or (_26590_, _26589_, _13035_);
  nand (_26591_, _26277_, _13035_);
  and (_26592_, _26591_, _01320_);
  and (_26593_, _26592_, _26590_);
  or (_26594_, _26593_, _26260_);
  and (_42988_, _26594_, _42355_);
  and (_26595_, _12178_, _06566_);
  and (_26596_, _12178_, _06559_);
  or (_26598_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  or (_26599_, _12178_, _05619_);
  and (_26600_, _26599_, _26598_);
  or (_26601_, _26600_, _12129_);
  or (_26602_, _09436_, _12782_);
  or (_26603_, _26600_, _12767_);
  or (_26604_, _26600_, _12749_);
  or (_26605_, _26600_, _12244_);
  or (_26606_, _26600_, _12695_);
  or (_26607_, _12178_, _09015_);
  nand (_26609_, _12179_, _06266_);
  or (_26610_, _25304_, _12178_);
  or (_26611_, _26600_, _12255_);
  and (_26612_, _08913_, _07152_);
  nand (_26613_, _12179_, _07143_);
  and (_26614_, _26613_, _06756_);
  and (_26615_, _07454_, \oc8051_golden_model_1.PC [5]);
  or (_26616_, _26615_, _07143_);
  and (_26617_, _26616_, _26614_);
  not (_26618_, _24975_);
  and (_26620_, _26600_, _26618_);
  or (_26621_, _26620_, _12448_);
  or (_26622_, _26621_, _26617_);
  and (_26623_, _26622_, _07858_);
  or (_26624_, _26623_, _26612_);
  or (_26625_, _26600_, _12453_);
  and (_26626_, _26625_, _26624_);
  or (_26627_, _26626_, _08734_);
  and (_26628_, _12430_, _12178_);
  or (_26629_, _12181_, _12180_);
  nand (_26631_, _26629_, _12204_);
  or (_26632_, _26629_, _12204_);
  and (_26633_, _26632_, _26631_);
  and (_26634_, _26633_, _12432_);
  or (_26635_, _26634_, _08736_);
  or (_26636_, _26635_, _26628_);
  and (_26637_, _26636_, _26627_);
  or (_26638_, _26637_, _07159_);
  or (_26639_, _26600_, _08639_);
  and (_26640_, _26639_, _06286_);
  and (_26642_, _26640_, _26638_);
  and (_26643_, _12418_, _12303_);
  or (_26644_, _12305_, _12304_);
  nand (_26645_, _26644_, _12334_);
  or (_26646_, _26644_, _12334_);
  and (_26647_, _26646_, _26645_);
  and (_26648_, _26647_, _12420_);
  or (_26649_, _26648_, _26643_);
  and (_26650_, _26649_, _06285_);
  or (_26651_, _26650_, _12410_);
  or (_26652_, _26651_, _26642_);
  or (_26653_, _26600_, _12409_);
  and (_26654_, _26653_, _06282_);
  and (_26655_, _26654_, _26652_);
  and (_26656_, _12178_, _06281_);
  or (_26657_, _26656_, _07460_);
  or (_26658_, _26657_, _26655_);
  or (_26659_, _08913_, _05949_);
  and (_26660_, _26659_, _07169_);
  and (_26661_, _26660_, _26658_);
  nand (_26662_, _12178_, _06354_);
  nand (_26663_, _26662_, _12404_);
  or (_26664_, _26663_, _26661_);
  or (_26665_, _26600_, _12404_);
  and (_26666_, _26665_, _06346_);
  and (_26667_, _26666_, _26664_);
  nand (_26668_, _12178_, _06345_);
  nand (_26669_, _26668_, _12468_);
  or (_26670_, _26669_, _26667_);
  or (_26671_, _26600_, _12468_);
  and (_26674_, _26671_, _06278_);
  and (_26675_, _26674_, _26670_);
  and (_26676_, _12178_, _06277_);
  or (_26677_, _26676_, _12475_);
  or (_26678_, _26677_, _26675_);
  or (_26679_, _08913_, _05955_);
  and (_26680_, _26679_, _06778_);
  and (_26681_, _26680_, _26678_);
  nand (_26682_, _12178_, _06276_);
  nand (_26683_, _26682_, _12484_);
  or (_26685_, _26683_, _26681_);
  and (_26686_, _12519_, _12303_);
  and (_26687_, _26647_, _25019_);
  or (_26688_, _26687_, _26686_);
  or (_26689_, _26688_, _12484_);
  and (_26690_, _26689_, _26685_);
  or (_26691_, _26690_, _06423_);
  and (_26692_, _12400_, _12303_);
  and (_26693_, _26647_, _12398_);
  or (_26694_, _26693_, _26692_);
  or (_26696_, _26694_, _06424_);
  and (_26697_, _26696_, _26691_);
  or (_26698_, _26697_, _06347_);
  and (_26699_, _26647_, _25279_);
  and (_26700_, _12540_, _12303_);
  or (_26701_, _26700_, _14105_);
  or (_26702_, _26701_, _26699_);
  and (_26703_, _26702_, _12528_);
  and (_26704_, _26703_, _26698_);
  or (_26705_, _26647_, _12559_);
  or (_26707_, _12560_, _12303_);
  and (_26708_, _26707_, _06419_);
  and (_26709_, _26708_, _26705_);
  or (_26710_, _26709_, _12254_);
  or (_26711_, _26710_, _26704_);
  and (_26712_, _26711_, _26611_);
  or (_26713_, _26712_, _06270_);
  nand (_26714_, _12179_, _06270_);
  and (_26715_, _26714_, _05946_);
  and (_26716_, _26715_, _26713_);
  and (_26717_, _08913_, _07458_);
  or (_26718_, _26717_, _25305_);
  or (_26719_, _26718_, _26716_);
  and (_26720_, _26719_, _26610_);
  or (_26721_, _26720_, _12589_);
  or (_26722_, _26600_, _12585_);
  and (_26723_, _26722_, _14014_);
  and (_26724_, _26723_, _26721_);
  and (_26725_, _12178_, _06371_);
  or (_26726_, _26725_, _25318_);
  or (_26728_, _26726_, _26724_);
  or (_26729_, _08913_, _05953_);
  and (_26730_, _26729_, _14013_);
  and (_26731_, _26730_, _26728_);
  nand (_26732_, _12178_, _06370_);
  nand (_26733_, _26732_, _12595_);
  or (_26734_, _26733_, _26731_);
  or (_26735_, _26600_, _12595_);
  and (_26736_, _26735_, _26734_);
  or (_26737_, _26736_, _12600_);
  or (_26739_, _12178_, _12599_);
  and (_26740_, _26739_, _05940_);
  and (_26741_, _26740_, _26737_);
  and (_26742_, _26600_, _05976_);
  or (_26743_, _26742_, _06266_);
  or (_26744_, _26743_, _26741_);
  and (_26745_, _26744_, _26609_);
  or (_26746_, _26745_, _05974_);
  or (_26747_, _08913_, _15174_);
  and (_26748_, _26747_, _06396_);
  and (_26750_, _26748_, _26746_);
  nand (_26751_, _12303_, _06395_);
  nand (_26752_, _26751_, _06261_);
  or (_26753_, _26752_, _26750_);
  or (_26754_, _12178_, _06261_);
  and (_26755_, _26754_, _06251_);
  and (_26756_, _26755_, _26753_);
  nand (_26757_, _12303_, _05972_);
  nand (_26758_, _26757_, _12252_);
  or (_26759_, _26758_, _26756_);
  or (_26761_, _26600_, _12252_);
  and (_26762_, _26761_, _06854_);
  and (_26763_, _26762_, _26759_);
  and (_26764_, _12178_, _06330_);
  or (_26765_, _26764_, _05997_);
  or (_26766_, _26765_, _26763_);
  or (_26767_, _08913_, _05998_);
  and (_26768_, _26767_, _12631_);
  and (_26769_, _26768_, _26766_);
  and (_26770_, _26633_, _12630_);
  or (_26772_, _26770_, _09016_);
  or (_26773_, _26772_, _26769_);
  and (_26774_, _26773_, _26607_);
  or (_26775_, _26774_, _06215_);
  or (_26776_, _12303_, _06216_);
  and (_26777_, _26776_, _10892_);
  and (_26778_, _26777_, _26775_);
  and (_26779_, _12178_, _10891_);
  or (_26780_, _26779_, _12644_);
  or (_26781_, _26780_, _26778_);
  nor (_26782_, _12662_, _12655_);
  or (_26783_, _26782_, _12663_);
  nand (_26784_, _26783_, _12644_);
  and (_26785_, _26784_, _06860_);
  and (_26786_, _26785_, _26781_);
  and (_26787_, _12178_, _06329_);
  or (_26788_, _26787_, _06004_);
  or (_26789_, _26788_, _26786_);
  or (_26790_, _08913_, _13852_);
  and (_26791_, _26790_, _12685_);
  and (_26793_, _26791_, _26789_);
  or (_26794_, _26633_, _11327_);
  nand (_26795_, _12179_, _11327_);
  and (_26796_, _26795_, _12247_);
  and (_26797_, _26796_, _26794_);
  or (_26798_, _26797_, _12697_);
  or (_26799_, _26798_, _26793_);
  and (_26800_, _26799_, _26606_);
  or (_26801_, _26800_, _12700_);
  or (_26802_, _12699_, _12178_);
  and (_26804_, _26802_, _09025_);
  and (_26805_, _26804_, _26801_);
  and (_26806_, _12303_, _06398_);
  or (_26807_, _26806_, _06524_);
  or (_26808_, _26807_, _26805_);
  nand (_26809_, _12179_, _06524_);
  and (_26810_, _26809_, _26808_);
  or (_26811_, _26810_, _06001_);
  not (_26812_, _06001_);
  or (_26813_, _08913_, _26812_);
  and (_26815_, _26813_, _12712_);
  and (_26816_, _26815_, _26811_);
  or (_26817_, _26633_, _12248_);
  or (_26818_, _12178_, _11327_);
  and (_26819_, _26818_, _12711_);
  and (_26820_, _26819_, _26817_);
  or (_26821_, _26820_, _12720_);
  or (_26822_, _26821_, _26816_);
  and (_26823_, _26822_, _26605_);
  or (_26824_, _26823_, _10970_);
  or (_26826_, _12178_, _10969_);
  and (_26827_, _26826_, _07219_);
  and (_26828_, _26827_, _26824_);
  and (_26829_, _12303_, _06426_);
  or (_26830_, _26829_, _06532_);
  or (_26831_, _26830_, _26828_);
  nand (_26832_, _12179_, _06532_);
  and (_26833_, _26832_, _26831_);
  or (_26834_, _26833_, _06013_);
  or (_26835_, _08913_, _15250_);
  and (_26837_, _26835_, _12733_);
  and (_26838_, _26837_, _26834_);
  or (_26839_, _26633_, \oc8051_golden_model_1.PSW [7]);
  or (_26840_, _12178_, _10774_);
  and (_26841_, _26840_, _12732_);
  and (_26842_, _26841_, _26839_);
  or (_26843_, _26842_, _12751_);
  or (_26844_, _26843_, _26838_);
  and (_26845_, _26844_, _26604_);
  or (_26846_, _26845_, _11008_);
  or (_26847_, _12178_, _11007_);
  and (_26848_, _26847_, _07229_);
  and (_26849_, _26848_, _26846_);
  and (_26850_, _12303_, _06437_);
  or (_26851_, _26850_, _06535_);
  or (_26852_, _26851_, _26849_);
  nand (_26853_, _12179_, _06535_);
  and (_26854_, _26853_, _26852_);
  or (_26855_, _26854_, _06008_);
  or (_26856_, _08913_, _06009_);
  and (_26858_, _26856_, _12762_);
  and (_26859_, _26858_, _26855_);
  or (_26860_, _26633_, _10774_);
  or (_26861_, _12178_, \oc8051_golden_model_1.PSW [7]);
  and (_26862_, _26861_, _12239_);
  and (_26863_, _26862_, _26860_);
  or (_26864_, _26863_, _12771_);
  or (_26865_, _26864_, _26859_);
  and (_26866_, _26865_, _26603_);
  or (_26867_, _26866_, _12770_);
  or (_26869_, _12178_, _12769_);
  and (_26870_, _26869_, _12775_);
  and (_26871_, _26870_, _26867_);
  and (_26872_, _26600_, _11111_);
  or (_26873_, _26872_, _06543_);
  or (_26874_, _26873_, _26871_);
  and (_26875_, _26874_, _26602_);
  or (_26876_, _26875_, _06011_);
  or (_26877_, _08913_, _09057_);
  and (_26878_, _26877_, _12786_);
  and (_26880_, _26878_, _26876_);
  or (_26881_, _26647_, _25133_);
  or (_26882_, _12303_, _12970_);
  and (_26883_, _26882_, _06436_);
  and (_26884_, _26883_, _26881_);
  or (_26885_, _26884_, _12790_);
  or (_26886_, _26885_, _26880_);
  and (_26887_, _26886_, _26601_);
  or (_26888_, _26887_, _12979_);
  or (_26889_, _12978_, _12178_);
  and (_26891_, _26889_, _12981_);
  and (_26892_, _26891_, _26888_);
  and (_26893_, _26600_, _10472_);
  or (_26894_, _26893_, _06290_);
  or (_26895_, _26894_, _26892_);
  or (_26896_, _09436_, _06291_);
  and (_26897_, _26896_, _26895_);
  or (_26898_, _26897_, _05994_);
  or (_26899_, _08913_, _25143_);
  and (_26900_, _26899_, _06435_);
  and (_26902_, _26900_, _26898_);
  or (_26903_, _12303_, _25133_);
  or (_26904_, _26647_, _12970_);
  and (_26905_, _26904_, _26903_);
  and (_26906_, _26905_, _06434_);
  or (_26907_, _26906_, _12999_);
  or (_26908_, _26907_, _26902_);
  or (_26909_, _26600_, _12998_);
  and (_26910_, _26909_, _07240_);
  and (_26911_, _26910_, _26908_);
  or (_26912_, _26911_, _26596_);
  and (_26913_, _26912_, _13005_);
  not (_26914_, _13005_);
  and (_26915_, _26600_, _26914_);
  or (_26916_, _26915_, _07678_);
  or (_26917_, _26916_, _26913_);
  or (_26918_, _08913_, _07252_);
  and (_26919_, _26918_, _05933_);
  and (_26920_, _26919_, _26917_);
  and (_26921_, _26905_, _05932_);
  or (_26923_, _26921_, _13020_);
  or (_26924_, _26923_, _26920_);
  or (_26925_, _26600_, _13019_);
  and (_26926_, _26925_, _06570_);
  and (_26927_, _26926_, _26924_);
  or (_26928_, _26927_, _26595_);
  and (_26929_, _26928_, _13027_);
  not (_26930_, _13027_);
  and (_26931_, _26600_, _26930_);
  or (_26932_, _26931_, _25169_);
  or (_26934_, _26932_, _26929_);
  or (_26935_, _25167_, _08913_);
  and (_26936_, _26935_, _13039_);
  and (_26937_, _26936_, _26934_);
  and (_26938_, _26600_, _13035_);
  or (_26939_, _26938_, _01324_);
  or (_26940_, _26939_, _26937_);
  or (_26941_, _01320_, \oc8051_golden_model_1.PC [5]);
  and (_26942_, _26941_, _42355_);
  and (_42989_, _26942_, _26940_);
  nand (_26944_, _08844_, _07678_);
  and (_26945_, _08739_, _12116_);
  nor (_26946_, _26945_, \oc8051_golden_model_1.PC [6]);
  nor (_26947_, _26946_, _12117_);
  not (_26948_, _26947_);
  nand (_26949_, _26948_, _10472_);
  nand (_26950_, _26948_, _12254_);
  nand (_26951_, _12172_, _06277_);
  or (_26952_, _26947_, _12404_);
  or (_26953_, _12336_, _12300_);
  and (_26955_, _26953_, _12337_);
  or (_26956_, _26955_, _12418_);
  or (_26957_, _12420_, _12296_);
  and (_26958_, _26957_, _06285_);
  and (_26959_, _26958_, _26956_);
  and (_26960_, _12430_, _12171_);
  or (_26961_, _12206_, _12175_);
  and (_26962_, _26961_, _12207_);
  and (_26963_, _26962_, _12432_);
  or (_26964_, _26963_, _26960_);
  or (_26966_, _26964_, _08736_);
  nand (_26967_, _08844_, _07152_);
  nand (_26968_, _12172_, _07143_);
  and (_26969_, _26968_, _06756_);
  and (_26970_, _07454_, \oc8051_golden_model_1.PC [6]);
  or (_26971_, _26970_, _07143_);
  and (_26972_, _26971_, _26969_);
  nor (_26973_, _26948_, _24975_);
  or (_26974_, _26973_, _07152_);
  or (_26975_, _26974_, _26972_);
  and (_26977_, _26975_, _12453_);
  and (_26978_, _26977_, _26967_);
  and (_26979_, _26947_, _12448_);
  or (_26980_, _26979_, _08734_);
  or (_26981_, _26980_, _26978_);
  and (_26982_, _26981_, _12457_);
  and (_26983_, _26982_, _26966_);
  or (_26984_, _26983_, _26959_);
  and (_26985_, _26984_, _12409_);
  nor (_26986_, _26948_, _12411_);
  or (_26988_, _26986_, _06281_);
  or (_26989_, _26988_, _26985_);
  nand (_26990_, _12172_, _06281_);
  and (_26991_, _26990_, _05949_);
  and (_26992_, _26991_, _26989_);
  nor (_26993_, _08844_, _05949_);
  or (_26994_, _26993_, _06354_);
  or (_26995_, _26994_, _26992_);
  nand (_26996_, _12172_, _06354_);
  and (_26997_, _26996_, _26995_);
  or (_26998_, _26997_, _26288_);
  and (_26999_, _26998_, _26952_);
  or (_27000_, _26999_, _06345_);
  nand (_27001_, _12172_, _06345_);
  and (_27002_, _27001_, _12468_);
  and (_27003_, _27002_, _27000_);
  nor (_27004_, _26948_, _12468_);
  or (_27005_, _27004_, _06277_);
  or (_27006_, _27005_, _27003_);
  and (_27007_, _27006_, _26951_);
  or (_27009_, _27007_, _12475_);
  nand (_27010_, _08844_, _12475_);
  and (_27011_, _27010_, _06778_);
  nand (_27012_, _27011_, _27009_);
  nand (_27013_, _12171_, _06276_);
  and (_27014_, _27013_, _12484_);
  and (_27015_, _27014_, _27012_);
  not (_27016_, _26955_);
  or (_27017_, _27016_, _12519_);
  nand (_27018_, _12519_, _12296_);
  and (_27020_, _27018_, _12485_);
  and (_27021_, _27020_, _27017_);
  or (_27022_, _27021_, _27015_);
  nand (_27023_, _27022_, _06424_);
  or (_27024_, _12398_, _12297_);
  or (_27025_, _27016_, _12400_);
  and (_27026_, _27025_, _06423_);
  and (_27027_, _27026_, _27024_);
  nor (_27028_, _27027_, _06347_);
  and (_27029_, _27028_, _27023_);
  nor (_27031_, _27016_, _12540_);
  and (_27032_, _12540_, _12296_);
  or (_27033_, _27032_, _27031_);
  and (_27034_, _27033_, _06347_);
  or (_27035_, _27034_, _27029_);
  and (_27036_, _27035_, _12528_);
  or (_27037_, _26955_, _12559_);
  nand (_27038_, _12559_, _12297_);
  and (_27039_, _27038_, _06419_);
  and (_27040_, _27039_, _27037_);
  or (_27042_, _27040_, _12254_);
  or (_27043_, _27042_, _27036_);
  and (_27044_, _27043_, _26950_);
  or (_27045_, _27044_, _06270_);
  nand (_27046_, _12172_, _06270_);
  and (_27047_, _27046_, _05946_);
  and (_27048_, _27047_, _27045_);
  nor (_27049_, _08844_, _05946_);
  or (_27050_, _27049_, _25305_);
  or (_27051_, _27050_, _27048_);
  or (_27053_, _25304_, _12171_);
  and (_27054_, _27053_, _27051_);
  or (_27055_, _27054_, _12589_);
  or (_27056_, _26947_, _12585_);
  and (_27057_, _27056_, _14014_);
  and (_27058_, _27057_, _27055_);
  and (_27059_, _12171_, _06371_);
  or (_27060_, _27059_, _25318_);
  or (_27061_, _27060_, _27058_);
  nand (_27062_, _08844_, _25318_);
  and (_27063_, _27062_, _14013_);
  and (_27064_, _27063_, _27061_);
  nand (_27065_, _12171_, _06370_);
  nand (_27066_, _27065_, _12595_);
  or (_27067_, _27066_, _27064_);
  or (_27068_, _26947_, _12595_);
  and (_27069_, _27068_, _12599_);
  and (_27070_, _27069_, _27067_);
  nor (_27071_, _12172_, _12599_);
  or (_27072_, _27071_, _05976_);
  or (_27074_, _27072_, _27070_);
  or (_27075_, _26947_, _05940_);
  and (_27076_, _27075_, _27074_);
  or (_27077_, _27076_, _06266_);
  nand (_27078_, _12172_, _06266_);
  and (_27079_, _27078_, _15174_);
  and (_27080_, _27079_, _27077_);
  nor (_27081_, _08844_, _15174_);
  or (_27082_, _27081_, _06395_);
  or (_27083_, _27082_, _27080_);
  nand (_27085_, _12297_, _06395_);
  and (_27086_, _27085_, _06261_);
  and (_27087_, _27086_, _27083_);
  nor (_27088_, _12172_, _06261_);
  or (_27089_, _27088_, _05972_);
  or (_27090_, _27089_, _27087_);
  nand (_27091_, _12297_, _05972_);
  and (_27092_, _27091_, _12252_);
  and (_27093_, _27092_, _27090_);
  nor (_27094_, _26948_, _12252_);
  or (_27096_, _27094_, _06330_);
  or (_27097_, _27096_, _27093_);
  nand (_27098_, _12172_, _06330_);
  and (_27099_, _27098_, _05998_);
  and (_27100_, _27099_, _27097_);
  nor (_27101_, _08844_, _05998_);
  or (_27102_, _27101_, _12630_);
  or (_27103_, _27102_, _27100_);
  or (_27104_, _26962_, _12631_);
  and (_27105_, _27104_, _09015_);
  and (_27107_, _27105_, _27103_);
  nor (_27108_, _12172_, _09015_);
  or (_27109_, _27108_, _06215_);
  or (_27110_, _27109_, _27107_);
  nand (_27111_, _12297_, _06215_);
  and (_27112_, _27111_, _10892_);
  and (_27113_, _27112_, _27110_);
  and (_27114_, _12171_, _10891_);
  or (_27115_, _27114_, _12644_);
  or (_27116_, _27115_, _27113_);
  or (_27118_, _12664_, _12652_);
  and (_27119_, _27118_, _12665_);
  or (_27120_, _27119_, _25380_);
  and (_27121_, _27120_, _06860_);
  and (_27122_, _27121_, _27116_);
  and (_27123_, _12171_, _06329_);
  or (_27124_, _27123_, _06004_);
  or (_27125_, _27124_, _27122_);
  nand (_27126_, _08844_, _06004_);
  and (_27127_, _27126_, _12685_);
  and (_27129_, _27127_, _27125_);
  or (_27130_, _26962_, _11327_);
  nand (_27131_, _12172_, _11327_);
  and (_27132_, _27131_, _12247_);
  and (_27133_, _27132_, _27130_);
  or (_27134_, _27133_, _12697_);
  or (_27135_, _27134_, _27129_);
  or (_27136_, _26947_, _12695_);
  and (_27137_, _27136_, _12699_);
  and (_27138_, _27137_, _27135_);
  nor (_27140_, _12699_, _12172_);
  or (_27141_, _27140_, _06398_);
  or (_27142_, _27141_, _27138_);
  nand (_27143_, _12297_, _06398_);
  and (_27144_, _27143_, _27142_);
  or (_27145_, _27144_, _06524_);
  nand (_27146_, _12172_, _06524_);
  and (_27147_, _27146_, _26812_);
  and (_27148_, _27147_, _27145_);
  nor (_27149_, _08844_, _26812_);
  or (_27151_, _27149_, _27148_);
  and (_27152_, _27151_, _12712_);
  or (_27153_, _26962_, _12248_);
  or (_27154_, _12171_, _11327_);
  and (_27155_, _27154_, _12711_);
  and (_27156_, _27155_, _27153_);
  or (_27157_, _27156_, _12720_);
  or (_27158_, _27157_, _27152_);
  or (_27159_, _26947_, _12244_);
  and (_27160_, _27159_, _10969_);
  and (_27162_, _27160_, _27158_);
  nor (_27163_, _12172_, _10969_);
  or (_27164_, _27163_, _06426_);
  or (_27165_, _27164_, _27162_);
  nand (_27166_, _12297_, _06426_);
  and (_27167_, _27166_, _27165_);
  or (_27168_, _27167_, _06532_);
  nand (_27169_, _12172_, _06532_);
  and (_27170_, _27169_, _15250_);
  and (_27171_, _27170_, _27168_);
  nor (_27173_, _08844_, _15250_);
  or (_27174_, _27173_, _27171_);
  and (_27175_, _27174_, _12733_);
  or (_27176_, _26962_, \oc8051_golden_model_1.PSW [7]);
  or (_27177_, _12171_, _10774_);
  and (_27178_, _27177_, _12732_);
  and (_27179_, _27178_, _27176_);
  or (_27180_, _27179_, _12751_);
  or (_27181_, _27180_, _27175_);
  or (_27182_, _26947_, _12749_);
  and (_27184_, _27182_, _11007_);
  and (_27185_, _27184_, _27181_);
  nor (_27186_, _12172_, _11007_);
  or (_27187_, _27186_, _06437_);
  or (_27188_, _27187_, _27185_);
  nand (_27189_, _12297_, _06437_);
  and (_27190_, _27189_, _27188_);
  or (_27191_, _27190_, _06535_);
  nand (_27192_, _12172_, _06535_);
  and (_27193_, _27192_, _06009_);
  and (_27195_, _27193_, _27191_);
  nor (_27196_, _08844_, _06009_);
  or (_27197_, _27196_, _27195_);
  and (_27198_, _27197_, _12762_);
  or (_27199_, _26962_, _10774_);
  or (_27200_, _12171_, \oc8051_golden_model_1.PSW [7]);
  and (_27201_, _27200_, _12239_);
  and (_27202_, _27201_, _27199_);
  or (_27203_, _27202_, _12771_);
  or (_27204_, _27203_, _27198_);
  or (_27206_, _26947_, _12767_);
  and (_27207_, _27206_, _12769_);
  and (_27208_, _27207_, _27204_);
  nor (_27209_, _12172_, _12769_);
  or (_27210_, _27209_, _11111_);
  or (_27211_, _27210_, _27208_);
  nand (_27212_, _26948_, _11111_);
  and (_27213_, _27212_, _12782_);
  and (_27214_, _27213_, _27211_);
  and (_27215_, _09435_, _06543_);
  or (_27217_, _27215_, _06011_);
  or (_27218_, _27217_, _27214_);
  nand (_27219_, _08844_, _06011_);
  and (_27220_, _27219_, _12786_);
  and (_27221_, _27220_, _27218_);
  nand (_27222_, _27016_, _12970_);
  or (_27223_, _12296_, _12970_);
  and (_27224_, _27223_, _06436_);
  and (_27225_, _27224_, _27222_);
  or (_27226_, _27225_, _12790_);
  or (_27228_, _27226_, _27221_);
  or (_27229_, _26947_, _12129_);
  and (_27230_, _27229_, _12978_);
  and (_27231_, _27230_, _27228_);
  nor (_27232_, _12978_, _12172_);
  or (_27233_, _27232_, _10472_);
  or (_27234_, _27233_, _27231_);
  and (_27235_, _27234_, _26949_);
  or (_27236_, _27235_, _06290_);
  or (_27237_, _09435_, _06291_);
  and (_27238_, _27237_, _25143_);
  and (_27239_, _27238_, _27236_);
  nor (_27240_, _08844_, _25143_);
  or (_27241_, _27240_, _06434_);
  or (_27242_, _27241_, _27239_);
  or (_27243_, _26955_, _12970_);
  nand (_27244_, _12297_, _12970_);
  and (_27245_, _27244_, _27243_);
  or (_27246_, _27245_, _06435_);
  and (_27247_, _27246_, _27242_);
  or (_27250_, _27247_, _12999_);
  or (_27251_, _26947_, _12998_);
  and (_27252_, _27251_, _27250_);
  or (_27253_, _27252_, _06559_);
  nand (_27254_, _12172_, _06559_);
  and (_27255_, _27254_, _13005_);
  and (_27256_, _27255_, _27253_);
  nor (_27257_, _26948_, _13005_);
  or (_27258_, _27257_, _07678_);
  or (_27259_, _27258_, _27256_);
  and (_27261_, _27259_, _26944_);
  or (_27262_, _27261_, _05932_);
  or (_27263_, _27245_, _05933_);
  and (_27264_, _27263_, _13019_);
  and (_27265_, _27264_, _27262_);
  nor (_27266_, _26948_, _13019_);
  or (_27267_, _27266_, _06566_);
  or (_27268_, _27267_, _27265_);
  nand (_27269_, _12172_, _06566_);
  and (_27270_, _27269_, _13027_);
  and (_27272_, _27270_, _27268_);
  nor (_27273_, _26948_, _13027_);
  or (_27274_, _27273_, _25169_);
  or (_27275_, _27274_, _27272_);
  nand (_27276_, _25169_, _08844_);
  and (_27277_, _27276_, _13039_);
  and (_27278_, _27277_, _27275_);
  and (_27279_, _26947_, _13035_);
  or (_27280_, _27279_, _01324_);
  or (_27281_, _27280_, _27278_);
  or (_27283_, _01320_, \oc8051_golden_model_1.PC [6]);
  and (_27284_, _27283_, _42355_);
  and (_42990_, _27284_, _27281_);
  and (_27285_, _08744_, _06566_);
  and (_27286_, _08744_, _06559_);
  nor (_27287_, _12117_, \oc8051_golden_model_1.PC [7]);
  nor (_27288_, _27287_, _12118_);
  or (_27289_, _27288_, _12129_);
  or (_27290_, _27288_, _12767_);
  or (_27291_, _27288_, _12749_);
  or (_27293_, _27288_, _12244_);
  or (_27294_, _27288_, _12695_);
  or (_27295_, _09015_, _08744_);
  or (_27296_, _27288_, _12595_);
  or (_27297_, _25304_, _08744_);
  or (_27298_, _27288_, _12255_);
  or (_27299_, _12167_, _12168_);
  nand (_27300_, _27299_, _12208_);
  or (_27301_, _27299_, _12208_);
  and (_27302_, _27301_, _27300_);
  and (_27304_, _27302_, _25203_);
  and (_27305_, _12430_, _08744_);
  or (_27306_, _27305_, _27304_);
  and (_27307_, _27306_, _08734_);
  nor (_27308_, _08582_, _07858_);
  nand (_27309_, _08773_, _07143_);
  and (_27310_, _27309_, _06756_);
  and (_27311_, _07454_, \oc8051_golden_model_1.PC [7]);
  or (_27312_, _27311_, _07143_);
  and (_27313_, _27312_, _27310_);
  and (_27315_, _27288_, _26618_);
  or (_27316_, _27315_, _12448_);
  or (_27317_, _27316_, _27313_);
  and (_27318_, _27317_, _07858_);
  or (_27319_, _27318_, _27308_);
  or (_27320_, _27288_, _12453_);
  and (_27321_, _27320_, _08736_);
  and (_27322_, _27321_, _27319_);
  or (_27323_, _27322_, _07159_);
  or (_27324_, _27323_, _27307_);
  or (_27326_, _27288_, _08639_);
  and (_27327_, _27326_, _06286_);
  and (_27328_, _27327_, _27324_);
  or (_27329_, _12292_, _12293_);
  nand (_27330_, _27329_, _12338_);
  or (_27331_, _27329_, _12338_);
  and (_27332_, _27331_, _27330_);
  and (_27333_, _27332_, _12420_);
  and (_27334_, _12418_, _09405_);
  or (_27335_, _27334_, _27333_);
  and (_27337_, _27335_, _06285_);
  or (_27338_, _27337_, _12410_);
  or (_27339_, _27338_, _27328_);
  or (_27340_, _27288_, _12409_);
  and (_27341_, _27340_, _06282_);
  and (_27342_, _27341_, _27339_);
  and (_27343_, _08744_, _06281_);
  or (_27344_, _27343_, _07460_);
  or (_27345_, _27344_, _27342_);
  nand (_27346_, _08582_, _07460_);
  and (_27348_, _27346_, _07169_);
  and (_27349_, _27348_, _27345_);
  nand (_27350_, _08744_, _06354_);
  nand (_27351_, _27350_, _12404_);
  or (_27352_, _27351_, _27349_);
  or (_27353_, _27288_, _12404_);
  and (_27354_, _27353_, _06346_);
  and (_27355_, _27354_, _27352_);
  nand (_27356_, _08744_, _06345_);
  nand (_27357_, _27356_, _12468_);
  or (_27359_, _27357_, _27355_);
  or (_27360_, _27288_, _12468_);
  and (_27361_, _27360_, _06278_);
  and (_27362_, _27361_, _27359_);
  and (_27363_, _08744_, _06277_);
  or (_27364_, _27363_, _12475_);
  or (_27365_, _27364_, _27362_);
  nand (_27366_, _08582_, _12475_);
  and (_27367_, _27366_, _06778_);
  and (_27368_, _27367_, _27365_);
  nand (_27370_, _08744_, _06276_);
  nand (_27371_, _27370_, _12484_);
  or (_27372_, _27371_, _27368_);
  and (_27373_, _27332_, _25019_);
  and (_27374_, _12519_, _09405_);
  or (_27375_, _27374_, _12484_);
  or (_27376_, _27375_, _27373_);
  and (_27377_, _27376_, _27372_);
  or (_27378_, _27377_, _06423_);
  or (_27379_, _27332_, _12400_);
  or (_27381_, _12398_, _09405_);
  and (_27382_, _27381_, _27379_);
  or (_27383_, _27382_, _06424_);
  and (_27384_, _27383_, _06420_);
  and (_27385_, _27384_, _27378_);
  or (_27386_, _27332_, _12559_);
  or (_27387_, _12560_, _09405_);
  and (_27388_, _27387_, _06419_);
  and (_27389_, _27388_, _27386_);
  or (_27390_, _27389_, _12254_);
  or (_27392_, _25279_, _09405_);
  or (_27393_, _27332_, _12540_);
  and (_27394_, _27393_, _06347_);
  and (_27395_, _27394_, _27392_);
  or (_27396_, _27395_, _27390_);
  or (_27397_, _27396_, _27385_);
  and (_27398_, _27397_, _27298_);
  or (_27399_, _27398_, _06270_);
  nand (_27400_, _08773_, _06270_);
  and (_27401_, _27400_, _05946_);
  and (_27403_, _27401_, _27399_);
  nor (_27404_, _08582_, _05946_);
  or (_27405_, _27404_, _25305_);
  or (_27406_, _27405_, _27403_);
  and (_27407_, _27406_, _27297_);
  or (_27408_, _27407_, _12589_);
  or (_27409_, _27288_, _12585_);
  and (_27410_, _27409_, _14014_);
  and (_27411_, _27410_, _27408_);
  and (_27412_, _08744_, _06371_);
  or (_27414_, _27412_, _25318_);
  or (_27415_, _27414_, _27411_);
  nand (_27416_, _08582_, _25318_);
  and (_27417_, _27416_, _14013_);
  and (_27418_, _27417_, _27415_);
  nand (_27419_, _08744_, _06370_);
  nand (_27420_, _27419_, _12595_);
  or (_27421_, _27420_, _27418_);
  and (_27422_, _27421_, _27296_);
  or (_27423_, _27422_, _12600_);
  or (_27425_, _12599_, _08744_);
  and (_27426_, _27425_, _05940_);
  and (_27427_, _27426_, _27423_);
  and (_27428_, _27288_, _05976_);
  or (_27429_, _27428_, _06266_);
  or (_27430_, _27429_, _27427_);
  nand (_27431_, _08773_, _06266_);
  and (_27432_, _27431_, _27430_);
  or (_27433_, _27432_, _05974_);
  nand (_27434_, _08582_, _05974_);
  and (_27436_, _27434_, _06396_);
  and (_27437_, _27436_, _27433_);
  nand (_27438_, _09405_, _06395_);
  nand (_27439_, _27438_, _06261_);
  or (_27440_, _27439_, _27437_);
  or (_27441_, _08744_, _06261_);
  and (_27442_, _27441_, _06251_);
  and (_27443_, _27442_, _27440_);
  nand (_27444_, _09405_, _05972_);
  nand (_27445_, _27444_, _12252_);
  or (_27447_, _27445_, _27443_);
  or (_27448_, _27288_, _12252_);
  and (_27449_, _27448_, _06854_);
  and (_27450_, _27449_, _27447_);
  and (_27451_, _08744_, _06330_);
  or (_27452_, _27451_, _05997_);
  or (_27453_, _27452_, _27450_);
  nand (_27454_, _08582_, _05997_);
  and (_27455_, _27454_, _12631_);
  and (_27456_, _27455_, _27453_);
  and (_27458_, _27302_, _12630_);
  or (_27459_, _27458_, _09016_);
  or (_27460_, _27459_, _27456_);
  and (_27461_, _27460_, _27295_);
  or (_27462_, _27461_, _06215_);
  or (_27463_, _09405_, _06216_);
  and (_27464_, _27463_, _10892_);
  and (_27465_, _27464_, _27462_);
  and (_27466_, _10891_, _08744_);
  or (_27467_, _27466_, _12644_);
  or (_27469_, _27467_, _27465_);
  not (_27470_, _12666_);
  or (_27471_, _12649_, _12648_);
  nor (_27472_, _27471_, _27470_);
  and (_27473_, _27471_, _27470_);
  or (_27474_, _27473_, _27472_);
  or (_27475_, _27474_, _25380_);
  and (_27476_, _27475_, _06860_);
  and (_27477_, _27476_, _27469_);
  and (_27478_, _08744_, _06329_);
  or (_27480_, _27478_, _06004_);
  or (_27481_, _27480_, _27477_);
  nand (_27482_, _08582_, _06004_);
  and (_27483_, _27482_, _12685_);
  and (_27484_, _27483_, _27481_);
  or (_27485_, _27302_, _11327_);
  nand (_27486_, _11327_, _08773_);
  and (_27487_, _27486_, _12247_);
  and (_27488_, _27487_, _27485_);
  or (_27489_, _27488_, _12697_);
  or (_27491_, _27489_, _27484_);
  and (_27492_, _27491_, _27294_);
  or (_27493_, _27492_, _12700_);
  or (_27494_, _12699_, _08744_);
  and (_27495_, _27494_, _09025_);
  and (_27496_, _27495_, _27493_);
  and (_27497_, _09405_, _06398_);
  or (_27498_, _27497_, _06524_);
  or (_27499_, _27498_, _27496_);
  nand (_27500_, _08773_, _06524_);
  and (_27502_, _27500_, _27499_);
  or (_27503_, _27502_, _06001_);
  nand (_27504_, _08582_, _06001_);
  and (_27505_, _27504_, _12712_);
  and (_27506_, _27505_, _27503_);
  or (_27507_, _27302_, _12248_);
  or (_27508_, _11327_, _08744_);
  and (_27509_, _27508_, _12711_);
  and (_27510_, _27509_, _27507_);
  or (_27511_, _27510_, _12720_);
  or (_27513_, _27511_, _27506_);
  and (_27514_, _27513_, _27293_);
  or (_27515_, _27514_, _10970_);
  or (_27516_, _10969_, _08744_);
  and (_27517_, _27516_, _07219_);
  and (_27518_, _27517_, _27515_);
  and (_27519_, _09405_, _06426_);
  or (_27520_, _27519_, _06532_);
  or (_27521_, _27520_, _27518_);
  nand (_27522_, _08773_, _06532_);
  and (_27524_, _27522_, _27521_);
  or (_27525_, _27524_, _06013_);
  nand (_27526_, _08582_, _06013_);
  and (_27527_, _27526_, _12733_);
  and (_27528_, _27527_, _27525_);
  or (_27529_, _27302_, \oc8051_golden_model_1.PSW [7]);
  or (_27530_, _08744_, _10774_);
  and (_27531_, _27530_, _12732_);
  and (_27532_, _27531_, _27529_);
  or (_27533_, _27532_, _12751_);
  or (_27535_, _27533_, _27528_);
  and (_27536_, _27535_, _27291_);
  or (_27537_, _27536_, _11008_);
  or (_27538_, _11007_, _08744_);
  and (_27539_, _27538_, _07229_);
  and (_27540_, _27539_, _27537_);
  and (_27541_, _09405_, _06437_);
  or (_27542_, _27541_, _06535_);
  or (_27543_, _27542_, _27540_);
  nand (_27544_, _08773_, _06535_);
  and (_27546_, _27544_, _27543_);
  or (_27547_, _27546_, _06008_);
  nand (_27548_, _08582_, _06008_);
  and (_27549_, _27548_, _12762_);
  and (_27550_, _27549_, _27547_);
  or (_27551_, _27302_, _10774_);
  or (_27552_, _08744_, \oc8051_golden_model_1.PSW [7]);
  and (_27553_, _27552_, _12239_);
  and (_27554_, _27553_, _27551_);
  or (_27555_, _27554_, _12771_);
  or (_27557_, _27555_, _27550_);
  and (_27558_, _27557_, _27290_);
  or (_27559_, _27558_, _12770_);
  or (_27560_, _12769_, _08744_);
  and (_27561_, _27560_, _12775_);
  and (_27562_, _27561_, _27559_);
  and (_27563_, _27288_, _11111_);
  or (_27564_, _27563_, _06543_);
  or (_27565_, _27564_, _27562_);
  or (_27566_, _08731_, _12782_);
  and (_27568_, _27566_, _27565_);
  or (_27569_, _27568_, _06011_);
  nand (_27570_, _08582_, _06011_);
  and (_27571_, _27570_, _12786_);
  and (_27572_, _27571_, _27569_);
  or (_27573_, _27332_, _25133_);
  or (_27574_, _09405_, _12970_);
  and (_27575_, _27574_, _06436_);
  and (_27576_, _27575_, _27573_);
  or (_27577_, _27576_, _12790_);
  or (_27579_, _27577_, _27572_);
  and (_27580_, _27579_, _27289_);
  or (_27581_, _27580_, _12979_);
  or (_27582_, _12978_, _08744_);
  and (_27583_, _27582_, _12981_);
  and (_27584_, _27583_, _27581_);
  and (_27585_, _27288_, _10472_);
  or (_27586_, _27585_, _06290_);
  or (_27587_, _27586_, _27584_);
  or (_27588_, _08731_, _06291_);
  and (_27590_, _27588_, _27587_);
  or (_27591_, _27590_, _05994_);
  nand (_27592_, _08582_, _05994_);
  and (_27593_, _27592_, _06435_);
  and (_27594_, _27593_, _27591_);
  or (_27595_, _09405_, _25133_);
  or (_27596_, _27332_, _12970_);
  and (_27597_, _27596_, _27595_);
  and (_27598_, _27597_, _06434_);
  or (_27599_, _27598_, _12999_);
  or (_27601_, _27599_, _27594_);
  or (_27602_, _27288_, _12998_);
  and (_27603_, _27602_, _07240_);
  and (_27604_, _27603_, _27601_);
  or (_27605_, _27604_, _27286_);
  and (_27606_, _27605_, _13005_);
  and (_27607_, _27288_, _26914_);
  or (_27608_, _27607_, _07678_);
  or (_27609_, _27608_, _27606_);
  nand (_27610_, _08582_, _07678_);
  and (_27612_, _27610_, _05933_);
  and (_27613_, _27612_, _27609_);
  and (_27614_, _27597_, _05932_);
  or (_27615_, _27614_, _13020_);
  or (_27616_, _27615_, _27613_);
  or (_27617_, _27288_, _13019_);
  and (_27618_, _27617_, _06570_);
  and (_27619_, _27618_, _27616_);
  or (_27620_, _27619_, _27285_);
  and (_27621_, _27620_, _13027_);
  and (_27623_, _27288_, _26930_);
  or (_27624_, _27623_, _25169_);
  or (_27625_, _27624_, _27621_);
  nand (_27626_, _25169_, _08582_);
  and (_27627_, _27626_, _13039_);
  and (_27628_, _27627_, _27625_);
  and (_27629_, _27288_, _13035_);
  or (_27630_, _27629_, _01324_);
  or (_27631_, _27630_, _27628_);
  or (_27632_, _01320_, \oc8051_golden_model_1.PC [7]);
  and (_27634_, _27632_, _42355_);
  and (_42991_, _27634_, _27631_);
  and (_27635_, _06432_, _06248_);
  or (_27636_, _12342_, _07219_);
  or (_27637_, _12212_, _09015_);
  or (_27638_, _12398_, _12342_);
  or (_27639_, _12345_, _12340_);
  and (_27640_, _27639_, _12346_);
  or (_27641_, _27640_, _12400_);
  and (_27642_, _27641_, _06423_);
  and (_27644_, _27642_, _27638_);
  and (_27645_, _12212_, _06277_);
  nor (_27646_, _06354_, _07460_);
  and (_27647_, _12212_, _06281_);
  or (_27648_, _12420_, _12342_);
  or (_27649_, _27640_, _12418_);
  and (_27650_, _27649_, _27648_);
  or (_27651_, _27650_, _06286_);
  and (_27652_, _12430_, _12212_);
  or (_27653_, _12215_, _12210_);
  and (_27655_, _27653_, _12216_);
  and (_27656_, _27655_, _12432_);
  or (_27657_, _27656_, _27652_);
  or (_27658_, _27657_, _08736_);
  nor (_27659_, _12118_, \oc8051_golden_model_1.PC [8]);
  nor (_27660_, _27659_, _12119_);
  or (_27661_, _27660_, _24975_);
  or (_27662_, _12212_, _07144_);
  nor (_27663_, _07143_, \oc8051_golden_model_1.PC [8]);
  nand (_27664_, _27663_, _07454_);
  and (_27666_, _27664_, _27662_);
  or (_27667_, _27666_, _06755_);
  and (_27668_, _27667_, _27661_);
  or (_27669_, _27668_, _25213_);
  or (_27670_, _27660_, _12453_);
  and (_27671_, _27670_, _27669_);
  or (_27672_, _27671_, _08734_);
  and (_27673_, _27672_, _08639_);
  and (_27674_, _27673_, _27658_);
  and (_27675_, _27660_, _07159_);
  or (_27677_, _27675_, _06285_);
  or (_27678_, _27677_, _27674_);
  and (_27679_, _27678_, _27651_);
  or (_27680_, _27679_, _12410_);
  or (_27681_, _27660_, _12409_);
  and (_27682_, _27681_, _06282_);
  and (_27683_, _27682_, _27680_);
  or (_27684_, _27683_, _27647_);
  and (_27685_, _27684_, _27646_);
  nand (_27686_, _12212_, _06354_);
  nand (_27688_, _27686_, _12404_);
  or (_27689_, _27688_, _27685_);
  or (_27690_, _27660_, _12404_);
  and (_27691_, _27690_, _06346_);
  and (_27692_, _27691_, _27689_);
  nand (_27693_, _12212_, _06345_);
  nand (_27694_, _27693_, _12468_);
  or (_27695_, _27694_, _27692_);
  or (_27696_, _27660_, _12468_);
  and (_27697_, _27696_, _06278_);
  and (_27699_, _27697_, _27695_);
  or (_27700_, _27699_, _27645_);
  and (_27701_, _27700_, _12476_);
  nand (_27702_, _12212_, _06276_);
  nand (_27703_, _27702_, _12484_);
  or (_27704_, _27703_, _27701_);
  and (_27705_, _12519_, _12342_);
  and (_27706_, _27640_, _25019_);
  or (_27707_, _27706_, _27705_);
  or (_27708_, _27707_, _12484_);
  and (_27710_, _27708_, _06424_);
  and (_27711_, _27710_, _27704_);
  or (_27712_, _27711_, _27644_);
  and (_27713_, _27712_, _06420_);
  and (_27714_, _12540_, _12342_);
  and (_27715_, _27640_, _25279_);
  or (_27716_, _27715_, _27714_);
  and (_27717_, _27716_, _06347_);
  or (_27718_, _27640_, _12559_);
  or (_27719_, _12560_, _12342_);
  and (_27721_, _27719_, _06419_);
  and (_27722_, _27721_, _27718_);
  or (_27723_, _27722_, _12254_);
  or (_27724_, _27723_, _27717_);
  or (_27725_, _27724_, _27713_);
  or (_27726_, _27660_, _12255_);
  and (_27727_, _27726_, _06271_);
  and (_27728_, _27727_, _27725_);
  and (_27729_, _12212_, _06270_);
  or (_27730_, _27729_, _07458_);
  or (_27732_, _27730_, _27728_);
  and (_27733_, _27732_, _25304_);
  and (_27734_, _25305_, _12212_);
  or (_27735_, _27734_, _12589_);
  or (_27736_, _27735_, _27733_);
  or (_27737_, _27660_, _12585_);
  and (_27738_, _27737_, _14014_);
  and (_27739_, _27738_, _27736_);
  and (_27740_, _12212_, _06371_);
  or (_27741_, _27740_, _25318_);
  or (_27743_, _27741_, _27739_);
  and (_27744_, _27743_, _14013_);
  nand (_27745_, _12212_, _06370_);
  nand (_27746_, _27745_, _12595_);
  or (_27747_, _27746_, _27744_);
  or (_27748_, _27660_, _12595_);
  and (_27749_, _27748_, _12599_);
  and (_27750_, _27749_, _27747_);
  and (_27751_, _12212_, _12600_);
  or (_27752_, _27751_, _05976_);
  or (_27754_, _27752_, _27750_);
  or (_27755_, _27660_, _05940_);
  and (_27756_, _27755_, _27754_);
  or (_27757_, _27756_, _06266_);
  or (_27758_, _12212_, _06267_);
  nor (_27759_, _06395_, _05974_);
  and (_27760_, _27759_, _27758_);
  and (_27761_, _27760_, _27757_);
  nand (_27762_, _12342_, _06395_);
  nand (_27763_, _27762_, _06261_);
  or (_27765_, _27763_, _27761_);
  or (_27766_, _12212_, _06261_);
  and (_27767_, _27766_, _06251_);
  and (_27768_, _27767_, _27765_);
  nand (_27769_, _12342_, _05972_);
  nand (_27770_, _27769_, _12252_);
  or (_27771_, _27770_, _27768_);
  or (_27772_, _27660_, _12252_);
  and (_27773_, _27772_, _06854_);
  and (_27774_, _27773_, _27771_);
  and (_27776_, _12212_, _06330_);
  or (_27777_, _27776_, _27774_);
  nor (_27778_, _12630_, _05997_);
  and (_27779_, _27778_, _27777_);
  and (_27780_, _27655_, _12630_);
  or (_27781_, _27780_, _09016_);
  or (_27782_, _27781_, _27779_);
  and (_27783_, _27782_, _27637_);
  or (_27784_, _27783_, _06215_);
  or (_27785_, _12342_, _06216_);
  and (_27787_, _27785_, _10892_);
  and (_27788_, _27787_, _27784_);
  and (_27789_, _12212_, _10891_);
  or (_27790_, _27789_, _12644_);
  or (_27791_, _27790_, _27788_);
  nor (_27792_, _12668_, \oc8051_golden_model_1.DPH [0]);
  nor (_27793_, _27792_, _12669_);
  or (_27794_, _27793_, _25380_);
  and (_27795_, _27794_, _06860_);
  and (_27796_, _27795_, _27791_);
  and (_27798_, _12212_, _06329_);
  or (_27799_, _27798_, _06004_);
  or (_27800_, _27799_, _27796_);
  and (_27801_, _27800_, _12685_);
  or (_27802_, _27655_, _11327_);
  or (_27803_, _12212_, _12248_);
  and (_27804_, _27803_, _12247_);
  and (_27805_, _27804_, _27802_);
  or (_27806_, _27805_, _12697_);
  or (_27807_, _27806_, _27801_);
  or (_27809_, _27660_, _12695_);
  and (_27810_, _27809_, _12699_);
  and (_27811_, _27810_, _27807_);
  and (_27812_, _12700_, _12212_);
  or (_27813_, _27812_, _06398_);
  or (_27814_, _27813_, _27811_);
  or (_27815_, _12342_, _09025_);
  and (_27816_, _27815_, _09030_);
  and (_27817_, _27816_, _27814_);
  and (_27818_, _12212_, _06524_);
  or (_27820_, _27818_, _06001_);
  or (_27821_, _27820_, _27817_);
  and (_27822_, _27821_, _12712_);
  or (_27823_, _27655_, _12248_);
  or (_27824_, _12212_, _11327_);
  and (_27825_, _27824_, _12711_);
  and (_27826_, _27825_, _27823_);
  or (_27827_, _27826_, _12720_);
  or (_27828_, _27827_, _27822_);
  or (_27829_, _27660_, _12244_);
  and (_27831_, _27829_, _10969_);
  and (_27832_, _27831_, _27828_);
  and (_27833_, _12212_, _10970_);
  or (_27834_, _27833_, _06426_);
  or (_27835_, _27834_, _27832_);
  and (_27836_, _27835_, _27636_);
  or (_27837_, _27836_, _06532_);
  or (_27838_, _12212_, _07217_);
  nor (_27839_, _12732_, _06013_);
  and (_27840_, _27839_, _27838_);
  and (_27842_, _27840_, _27837_);
  or (_27843_, _27655_, \oc8051_golden_model_1.PSW [7]);
  or (_27844_, _12212_, _10774_);
  and (_27845_, _27844_, _12732_);
  and (_27846_, _27845_, _27843_);
  or (_27847_, _27846_, _12751_);
  or (_27848_, _27847_, _27842_);
  or (_27849_, _27660_, _12749_);
  and (_27850_, _27849_, _11007_);
  and (_27851_, _27850_, _27848_);
  and (_27853_, _12212_, _11008_);
  or (_27854_, _27853_, _27851_);
  and (_27855_, _27854_, _07229_);
  and (_27856_, _12342_, _06437_);
  or (_27857_, _27856_, _06535_);
  or (_27858_, _27857_, _27855_);
  nor (_27859_, _12239_, _06008_);
  or (_27860_, _12212_, _07231_);
  and (_27861_, _27860_, _27859_);
  and (_27862_, _27861_, _27858_);
  or (_27864_, _27655_, _10774_);
  or (_27865_, _12212_, \oc8051_golden_model_1.PSW [7]);
  and (_27866_, _27865_, _12239_);
  and (_27867_, _27866_, _27864_);
  or (_27868_, _27867_, _12771_);
  or (_27869_, _27868_, _27862_);
  or (_27870_, _27660_, _12767_);
  and (_27871_, _27870_, _12769_);
  and (_27872_, _27871_, _27869_);
  and (_27873_, _12212_, _12770_);
  or (_27874_, _27873_, _11111_);
  or (_27875_, _27874_, _27872_);
  or (_27876_, _27660_, _12775_);
  and (_27877_, _27876_, _12782_);
  and (_27878_, _27877_, _27875_);
  and (_27879_, _07135_, _06543_);
  or (_27880_, _27879_, _06011_);
  or (_27881_, _27880_, _27878_);
  and (_27882_, _27881_, _12786_);
  or (_27883_, _27640_, _25133_);
  or (_27886_, _12342_, _12970_);
  and (_27887_, _27886_, _06436_);
  and (_27888_, _27887_, _27883_);
  or (_27889_, _27888_, _12790_);
  or (_27890_, _27889_, _27882_);
  or (_27891_, _27660_, _12129_);
  and (_27892_, _27891_, _12978_);
  and (_27893_, _27892_, _27890_);
  and (_27894_, _12979_, _12212_);
  or (_27895_, _27894_, _10472_);
  or (_27897_, _27895_, _27893_);
  or (_27898_, _27660_, _12981_);
  and (_27899_, _27898_, _06291_);
  and (_27900_, _27899_, _27897_);
  and (_27901_, _07135_, _06290_);
  or (_27902_, _27901_, _05994_);
  or (_27903_, _27902_, _27900_);
  and (_27904_, _27903_, _06435_);
  or (_27905_, _12342_, _25133_);
  or (_27906_, _27640_, _12970_);
  and (_27908_, _27906_, _27905_);
  and (_27909_, _27908_, _06434_);
  or (_27910_, _27909_, _12999_);
  or (_27911_, _27910_, _27904_);
  or (_27912_, _27660_, _12998_);
  and (_27913_, _27912_, _07240_);
  and (_27914_, _27913_, _27911_);
  nand (_27915_, _12212_, _06559_);
  nand (_27916_, _27915_, _13005_);
  or (_27917_, _27916_, _27914_);
  or (_27919_, _27660_, _13005_);
  and (_27920_, _27919_, _06433_);
  and (_27921_, _27920_, _27917_);
  or (_27922_, _27921_, _27635_);
  nor (_27923_, _05991_, _05932_);
  and (_27924_, _27923_, _27922_);
  and (_27925_, _27908_, _05932_);
  or (_27926_, _27925_, _13020_);
  or (_27927_, _27926_, _27924_);
  or (_27928_, _27660_, _13019_);
  and (_27930_, _27928_, _06570_);
  and (_27931_, _27930_, _27927_);
  nand (_27932_, _12212_, _06566_);
  nand (_27933_, _27932_, _13027_);
  or (_27934_, _27933_, _27931_);
  or (_27935_, _27660_, _13027_);
  and (_27936_, _27935_, _13030_);
  and (_27937_, _27936_, _27934_);
  and (_27938_, _06393_, _06248_);
  or (_27939_, _27938_, _27937_);
  and (_27941_, _27939_, _13036_);
  and (_27942_, _27660_, _13035_);
  or (_27943_, _27942_, _01324_);
  or (_27944_, _27943_, _27941_);
  or (_27945_, _01320_, \oc8051_golden_model_1.PC [8]);
  and (_27946_, _27945_, _42355_);
  and (_42992_, _27946_, _27944_);
  nor (_27947_, _06995_, _13030_);
  nor (_27948_, _06995_, _06433_);
  nor (_27949_, _12119_, \oc8051_golden_model_1.PC [9]);
  nor (_27951_, _27949_, _12120_);
  or (_27952_, _27951_, _12129_);
  or (_27953_, _27951_, _12767_);
  and (_27954_, _12287_, _06437_);
  or (_27955_, _27951_, _12749_);
  and (_27956_, _12287_, _06426_);
  or (_27957_, _27951_, _12244_);
  and (_27958_, _12287_, _06398_);
  or (_27959_, _27951_, _12695_);
  or (_27960_, _12162_, _09015_);
  and (_27962_, _12162_, _06330_);
  and (_27963_, _12162_, _06370_);
  or (_27964_, _27951_, _12585_);
  or (_27965_, _27951_, _12255_);
  or (_27966_, _12398_, _12287_);
  not (_27967_, _12343_);
  and (_27968_, _12346_, _27967_);
  and (_27969_, _27968_, _12290_);
  nor (_27970_, _27968_, _12290_);
  or (_27971_, _27970_, _27969_);
  or (_27973_, _27971_, _12400_);
  and (_27974_, _27973_, _06423_);
  and (_27975_, _27974_, _27966_);
  and (_27976_, _12430_, _12162_);
  not (_27977_, _12213_);
  and (_27978_, _12216_, _27977_);
  and (_27979_, _27978_, _12165_);
  nor (_27980_, _27978_, _12165_);
  or (_27981_, _27980_, _27979_);
  and (_27982_, _27981_, _12432_);
  or (_27984_, _27982_, _08736_);
  or (_27985_, _27984_, _27976_);
  and (_27986_, _27951_, _06755_);
  or (_27987_, _27951_, _12453_);
  or (_27988_, _07455_, \oc8051_golden_model_1.PC [9]);
  or (_27989_, _27951_, _07454_);
  and (_27990_, _27989_, _27988_);
  or (_27991_, _27990_, _07143_);
  or (_27992_, _12162_, _07144_);
  and (_27993_, _27992_, _06756_);
  and (_27995_, _27993_, _27991_);
  or (_27996_, _27995_, _25213_);
  and (_27997_, _27996_, _27987_);
  or (_27998_, _27997_, _08734_);
  or (_27999_, _27998_, _27986_);
  and (_28000_, _27999_, _27985_);
  or (_28001_, _28000_, _07159_);
  or (_28002_, _27951_, _08639_);
  and (_28003_, _28002_, _06286_);
  and (_28004_, _28003_, _28001_);
  or (_28006_, _27971_, _12418_);
  or (_28007_, _12420_, _12287_);
  and (_28008_, _28007_, _06285_);
  and (_28009_, _28008_, _28006_);
  or (_28010_, _28009_, _12410_);
  or (_28011_, _28010_, _28004_);
  or (_28012_, _27951_, _12409_);
  and (_28013_, _28012_, _06282_);
  and (_28014_, _28013_, _28011_);
  and (_28015_, _12162_, _06281_);
  or (_28017_, _28015_, _07460_);
  or (_28018_, _28017_, _28014_);
  and (_28019_, _28018_, _07169_);
  nand (_28020_, _12162_, _06354_);
  nand (_28021_, _28020_, _12404_);
  or (_28022_, _28021_, _28019_);
  or (_28023_, _27951_, _12404_);
  and (_28024_, _28023_, _06346_);
  and (_28025_, _28024_, _28022_);
  nand (_28026_, _12162_, _06345_);
  nand (_28028_, _28026_, _12468_);
  or (_28029_, _28028_, _28025_);
  or (_28030_, _27951_, _12468_);
  and (_28031_, _28030_, _06278_);
  and (_28032_, _28031_, _28029_);
  and (_28033_, _12162_, _06277_);
  or (_28034_, _28033_, _12475_);
  or (_28035_, _28034_, _28032_);
  and (_28036_, _28035_, _06778_);
  nand (_28037_, _12162_, _06276_);
  nand (_28039_, _28037_, _12484_);
  or (_28040_, _28039_, _28036_);
  and (_28041_, _12519_, _12287_);
  and (_28042_, _27971_, _25019_);
  or (_28043_, _28042_, _28041_);
  or (_28044_, _28043_, _12484_);
  and (_28045_, _28044_, _06424_);
  and (_28046_, _28045_, _28040_);
  or (_28047_, _28046_, _27975_);
  and (_28048_, _28047_, _06420_);
  or (_28050_, _25279_, _12287_);
  or (_28051_, _27971_, _12540_);
  and (_28052_, _28051_, _06347_);
  and (_28053_, _28052_, _28050_);
  or (_28054_, _27971_, _12559_);
  or (_28055_, _12560_, _12287_);
  and (_28056_, _28055_, _06419_);
  and (_28057_, _28056_, _28054_);
  or (_28058_, _28057_, _12254_);
  or (_28059_, _28058_, _28053_);
  or (_28061_, _28059_, _28048_);
  and (_28062_, _28061_, _27965_);
  or (_28063_, _28062_, _06270_);
  or (_28064_, _12162_, _06271_);
  and (_28065_, _28064_, _12573_);
  and (_28066_, _28065_, _25303_);
  and (_28067_, _28066_, _28063_);
  and (_28068_, _25305_, _12162_);
  or (_28069_, _28068_, _12589_);
  or (_28070_, _28069_, _28067_);
  and (_28072_, _28070_, _27964_);
  or (_28073_, _28072_, _06371_);
  nor (_28074_, _06370_, _25318_);
  or (_28075_, _12162_, _14014_);
  and (_28076_, _28075_, _28074_);
  and (_28077_, _28076_, _28073_);
  or (_28078_, _28077_, _27963_);
  and (_28079_, _28078_, _12595_);
  and (_28080_, _27951_, _12601_);
  or (_28081_, _28080_, _12600_);
  or (_28083_, _28081_, _28079_);
  or (_28084_, _12162_, _12599_);
  and (_28085_, _28084_, _05940_);
  and (_28086_, _28085_, _28083_);
  and (_28087_, _27951_, _05976_);
  or (_28088_, _28087_, _06266_);
  or (_28089_, _28088_, _28086_);
  or (_28090_, _12162_, _06267_);
  and (_28091_, _28090_, _27759_);
  and (_28092_, _28091_, _28089_);
  nand (_28094_, _12287_, _06395_);
  nand (_28095_, _28094_, _06261_);
  or (_28096_, _28095_, _28092_);
  or (_28097_, _12162_, _06261_);
  and (_28098_, _28097_, _06251_);
  and (_28099_, _28098_, _28096_);
  nand (_28100_, _12287_, _05972_);
  nand (_28101_, _28100_, _12252_);
  or (_28102_, _28101_, _28099_);
  or (_28103_, _27951_, _12252_);
  and (_28105_, _28103_, _06854_);
  and (_28106_, _28105_, _28102_);
  or (_28107_, _28106_, _27962_);
  and (_28108_, _28107_, _27778_);
  and (_28109_, _27981_, _12630_);
  or (_28110_, _28109_, _09016_);
  or (_28111_, _28110_, _28108_);
  and (_28112_, _28111_, _27960_);
  or (_28113_, _28112_, _06215_);
  or (_28114_, _12287_, _06216_);
  and (_28116_, _28114_, _10892_);
  and (_28117_, _28116_, _28113_);
  and (_28118_, _12162_, _10891_);
  or (_28119_, _28118_, _12644_);
  or (_28120_, _28119_, _28117_);
  nor (_28121_, _12669_, \oc8051_golden_model_1.DPH [1]);
  nor (_28122_, _28121_, _12670_);
  or (_28123_, _28122_, _25380_);
  and (_28124_, _28123_, _06860_);
  and (_28125_, _28124_, _28120_);
  and (_28127_, _12162_, _06329_);
  or (_28128_, _28127_, _06004_);
  or (_28129_, _28128_, _28125_);
  and (_28130_, _28129_, _12685_);
  or (_28131_, _27981_, _11327_);
  or (_28132_, _12162_, _12248_);
  and (_28133_, _28132_, _12247_);
  and (_28134_, _28133_, _28131_);
  or (_28135_, _28134_, _12697_);
  or (_28136_, _28135_, _28130_);
  and (_28138_, _28136_, _27959_);
  or (_28139_, _28138_, _12700_);
  or (_28140_, _12699_, _12162_);
  and (_28141_, _28140_, _09025_);
  and (_28142_, _28141_, _28139_);
  or (_28143_, _28142_, _27958_);
  and (_28144_, _28143_, _09030_);
  and (_28145_, _12162_, _06524_);
  or (_28146_, _28145_, _06001_);
  or (_28147_, _28146_, _28144_);
  and (_28149_, _28147_, _12712_);
  or (_28150_, _27981_, _12248_);
  or (_28151_, _12162_, _11327_);
  and (_28152_, _28151_, _12711_);
  and (_28153_, _28152_, _28150_);
  or (_28154_, _28153_, _12720_);
  or (_28155_, _28154_, _28149_);
  and (_28156_, _28155_, _27957_);
  or (_28157_, _28156_, _10970_);
  or (_28158_, _12162_, _10969_);
  and (_28160_, _28158_, _07219_);
  and (_28161_, _28160_, _28157_);
  or (_28162_, _28161_, _27956_);
  and (_28163_, _28162_, _07217_);
  and (_28164_, _12162_, _06532_);
  or (_28165_, _28164_, _06013_);
  or (_28166_, _28165_, _28163_);
  and (_28167_, _28166_, _12733_);
  or (_28168_, _27981_, \oc8051_golden_model_1.PSW [7]);
  or (_28169_, _12162_, _10774_);
  and (_28171_, _28169_, _12732_);
  and (_28172_, _28171_, _28168_);
  or (_28173_, _28172_, _12751_);
  or (_28174_, _28173_, _28167_);
  and (_28175_, _28174_, _27955_);
  or (_28176_, _28175_, _11008_);
  or (_28177_, _12162_, _11007_);
  and (_28178_, _28177_, _07229_);
  and (_28179_, _28178_, _28176_);
  or (_28180_, _28179_, _27954_);
  and (_28181_, _28180_, _07231_);
  and (_28182_, _12162_, _06535_);
  or (_28183_, _28182_, _06008_);
  or (_28184_, _28183_, _28181_);
  and (_28185_, _28184_, _12762_);
  or (_28186_, _27981_, _10774_);
  or (_28187_, _12162_, \oc8051_golden_model_1.PSW [7]);
  and (_28188_, _28187_, _12239_);
  and (_28189_, _28188_, _28186_);
  or (_28190_, _28189_, _12771_);
  or (_28193_, _28190_, _28185_);
  and (_28194_, _28193_, _27953_);
  or (_28195_, _28194_, _12770_);
  or (_28196_, _12162_, _12769_);
  and (_28197_, _28196_, _12775_);
  and (_28198_, _28197_, _28195_);
  and (_28199_, _27951_, _11111_);
  or (_28200_, _28199_, _06543_);
  or (_28201_, _28200_, _28198_);
  or (_28202_, _09422_, _12782_);
  nor (_28204_, _06436_, _06011_);
  and (_28205_, _28204_, _28202_);
  and (_28206_, _28205_, _28201_);
  or (_28207_, _27971_, _25133_);
  or (_28208_, _12287_, _12970_);
  and (_28209_, _28208_, _06436_);
  and (_28210_, _28209_, _28207_);
  or (_28211_, _28210_, _12790_);
  or (_28212_, _28211_, _28206_);
  and (_28213_, _28212_, _27952_);
  or (_28215_, _28213_, _12979_);
  or (_28216_, _12978_, _12162_);
  and (_28217_, _28216_, _12981_);
  and (_28218_, _28217_, _28215_);
  and (_28219_, _27951_, _10472_);
  or (_28220_, _28219_, _06290_);
  or (_28221_, _28220_, _28218_);
  or (_28222_, _09422_, _06291_);
  nor (_28223_, _06434_, _05994_);
  and (_28224_, _28223_, _28222_);
  and (_28226_, _28224_, _28221_);
  or (_28227_, _27971_, _12970_);
  or (_28228_, _12287_, _25133_);
  and (_28229_, _28228_, _28227_);
  and (_28230_, _28229_, _06434_);
  or (_28231_, _28230_, _12999_);
  or (_28232_, _28231_, _28226_);
  or (_28233_, _27951_, _12998_);
  and (_28234_, _28233_, _07240_);
  and (_28235_, _28234_, _28232_);
  nand (_28237_, _12162_, _06559_);
  nand (_28238_, _28237_, _13005_);
  or (_28239_, _28238_, _28235_);
  or (_28240_, _27951_, _13005_);
  and (_28241_, _28240_, _06433_);
  and (_28242_, _28241_, _28239_);
  or (_28243_, _28242_, _27948_);
  and (_28244_, _28243_, _27923_);
  and (_28245_, _28229_, _05932_);
  or (_28246_, _28245_, _13020_);
  or (_28248_, _28246_, _28244_);
  or (_28249_, _27951_, _13019_);
  and (_28250_, _28249_, _06570_);
  and (_28251_, _28250_, _28248_);
  nand (_28252_, _12162_, _06566_);
  nand (_28253_, _28252_, _13027_);
  or (_28254_, _28253_, _28251_);
  or (_28255_, _27951_, _13027_);
  and (_28256_, _28255_, _13030_);
  and (_28257_, _28256_, _28254_);
  or (_28259_, _28257_, _27947_);
  and (_28260_, _28259_, _13036_);
  and (_28261_, _27951_, _13035_);
  or (_28262_, _28261_, _01324_);
  or (_28263_, _28262_, _28260_);
  or (_28264_, _01320_, \oc8051_golden_model_1.PC [9]);
  and (_28265_, _28264_, _42355_);
  and (_42993_, _28265_, _28263_);
  nor (_28266_, _12120_, \oc8051_golden_model_1.PC [10]);
  nor (_28267_, _28266_, _12121_);
  not (_28269_, _28267_);
  nand (_28270_, _28269_, _10472_);
  nand (_28271_, _28269_, _11111_);
  or (_28272_, _12281_, _07229_);
  or (_28273_, _12281_, _07219_);
  or (_28274_, _12281_, _09025_);
  nor (_28275_, _28269_, _12252_);
  and (_28276_, _14881_, _06370_);
  and (_28277_, _12400_, _12281_);
  or (_28278_, _12349_, _12347_);
  nand (_28280_, _28278_, _12284_);
  or (_28281_, _28278_, _12284_);
  and (_28282_, _28281_, _28280_);
  and (_28283_, _28282_, _12398_);
  or (_28284_, _28283_, _28277_);
  and (_28285_, _28284_, _06423_);
  nor (_28286_, _28269_, _12468_);
  or (_28287_, _28267_, _12404_);
  nor (_28288_, _28269_, _12411_);
  or (_28289_, _28282_, _12418_);
  or (_28291_, _12420_, _12281_);
  and (_28292_, _28291_, _06285_);
  and (_28293_, _28292_, _28289_);
  and (_28294_, _12430_, _12156_);
  or (_28295_, _12219_, _12217_);
  and (_28296_, _28295_, _12159_);
  nor (_28297_, _28295_, _12159_);
  nor (_28298_, _28297_, _28296_);
  and (_28299_, _28298_, _12432_);
  or (_28300_, _28299_, _28294_);
  or (_28302_, _28300_, _08736_);
  and (_28303_, _12156_, _07143_);
  and (_28304_, _07144_, \oc8051_golden_model_1.PC [10]);
  and (_28305_, _28304_, _07454_);
  or (_28306_, _28305_, _28303_);
  and (_28307_, _28306_, _06756_);
  or (_28308_, _28307_, _07152_);
  and (_28309_, _28308_, _12453_);
  nor (_28310_, _26618_, _12448_);
  nor (_28311_, _28310_, _28269_);
  or (_28313_, _28311_, _08734_);
  or (_28314_, _28313_, _28309_);
  and (_28315_, _28314_, _12457_);
  and (_28316_, _28315_, _28302_);
  or (_28317_, _28316_, _28293_);
  and (_28318_, _28317_, _12409_);
  or (_28319_, _28318_, _28288_);
  and (_28320_, _28319_, _06361_);
  nor (_28321_, _14881_, _06361_);
  nand (_28322_, _12404_, _05949_);
  or (_28324_, _28322_, _28321_);
  or (_28325_, _28324_, _28320_);
  and (_28326_, _28325_, _28287_);
  or (_28327_, _28326_, _06345_);
  nand (_28328_, _14881_, _06345_);
  and (_28329_, _28328_, _12468_);
  and (_28330_, _28329_, _28327_);
  or (_28331_, _28330_, _28286_);
  and (_28332_, _28331_, _06278_);
  and (_28333_, _12156_, _06277_);
  or (_28335_, _28333_, _12475_);
  or (_28336_, _28335_, _28332_);
  and (_28337_, _28336_, _06778_);
  nand (_28338_, _12156_, _06276_);
  nand (_28339_, _28338_, _12484_);
  or (_28340_, _28339_, _28337_);
  and (_28341_, _28282_, _25019_);
  and (_28342_, _12519_, _12281_);
  or (_28343_, _28342_, _12484_);
  or (_28344_, _28343_, _28341_);
  and (_28346_, _28344_, _06424_);
  and (_28347_, _28346_, _28340_);
  or (_28348_, _28347_, _28285_);
  and (_28349_, _28348_, _06420_);
  or (_28350_, _28282_, _12559_);
  or (_28351_, _12560_, _12281_);
  and (_28352_, _28351_, _06419_);
  and (_28353_, _28352_, _28350_);
  or (_28354_, _28353_, _12254_);
  or (_28355_, _28282_, _12540_);
  or (_28357_, _25279_, _12281_);
  and (_28358_, _28357_, _06347_);
  and (_28359_, _28358_, _28355_);
  or (_28360_, _28359_, _28354_);
  or (_28361_, _28360_, _28349_);
  nand (_28362_, _28269_, _12254_);
  and (_28363_, _28362_, _06271_);
  and (_28364_, _28363_, _28361_);
  or (_28365_, _28364_, _07458_);
  and (_28366_, _28365_, _25304_);
  nand (_28368_, _25304_, _06271_);
  and (_28369_, _28368_, _12156_);
  or (_28370_, _28369_, _12589_);
  or (_28371_, _28370_, _28366_);
  or (_28372_, _28267_, _12585_);
  and (_28373_, _28372_, _14014_);
  nand (_28374_, _28373_, _28371_);
  nand (_28375_, _12156_, _06371_);
  and (_28376_, _28375_, _28074_);
  and (_28377_, _28376_, _28374_);
  or (_28379_, _28377_, _28276_);
  and (_28380_, _28379_, _12595_);
  nor (_28381_, _28267_, _12595_);
  or (_28382_, _28381_, _12600_);
  or (_28383_, _28382_, _28380_);
  or (_28384_, _14881_, _12599_);
  and (_28385_, _28384_, _05940_);
  and (_28386_, _28385_, _28383_);
  nor (_28387_, _28267_, _05940_);
  or (_28388_, _28387_, _06266_);
  nor (_28390_, _28388_, _28386_);
  nand (_28391_, _12156_, _06266_);
  nand (_28392_, _28391_, _27759_);
  or (_28393_, _28392_, _28390_);
  or (_28394_, _12281_, _06396_);
  and (_28395_, _28394_, _06261_);
  and (_28396_, _28395_, _28393_);
  nor (_28397_, _14881_, _06261_);
  or (_28398_, _28397_, _05972_);
  or (_28399_, _28398_, _28396_);
  or (_28401_, _12281_, _06251_);
  and (_28402_, _28401_, _12252_);
  and (_28403_, _28402_, _28399_);
  or (_28404_, _28403_, _28275_);
  and (_28405_, _28404_, _06854_);
  nand (_28406_, _12156_, _06330_);
  nand (_28407_, _28406_, _27778_);
  or (_28408_, _28407_, _28405_);
  or (_28409_, _28298_, _12631_);
  and (_28410_, _28409_, _09015_);
  and (_28412_, _28410_, _28408_);
  nor (_28413_, _14881_, _09015_);
  or (_28414_, _28413_, _06215_);
  or (_28415_, _28414_, _28412_);
  or (_28416_, _12281_, _06216_);
  and (_28417_, _28416_, _10892_);
  and (_28418_, _28417_, _28415_);
  and (_28419_, _12156_, _10891_);
  or (_28420_, _28419_, _12644_);
  or (_28421_, _28420_, _28418_);
  nor (_28423_, _12670_, \oc8051_golden_model_1.DPH [2]);
  nor (_28424_, _28423_, _12671_);
  or (_28425_, _28424_, _25380_);
  and (_28426_, _28425_, _06860_);
  and (_28427_, _28426_, _28421_);
  and (_28428_, _12156_, _06329_);
  or (_28429_, _28428_, _28427_);
  nand (_28430_, _07387_, _05930_);
  and (_28431_, _28430_, _28429_);
  or (_28432_, _28298_, _11327_);
  or (_28434_, _12156_, _12248_);
  and (_28435_, _28434_, _12247_);
  and (_28436_, _28435_, _28432_);
  or (_28437_, _28436_, _12697_);
  or (_28438_, _28437_, _28431_);
  or (_28439_, _28267_, _12695_);
  and (_28440_, _28439_, _12699_);
  and (_28441_, _28440_, _28438_);
  nor (_28442_, _12699_, _14881_);
  or (_28443_, _28442_, _06398_);
  or (_28445_, _28443_, _28441_);
  and (_28446_, _28445_, _28274_);
  or (_28447_, _28446_, _06524_);
  nand (_28448_, _14881_, _06524_);
  nor (_28449_, _12711_, _06001_);
  and (_28450_, _28449_, _28448_);
  and (_28451_, _28450_, _28447_);
  or (_28452_, _28298_, _12248_);
  or (_28453_, _12156_, _11327_);
  and (_28454_, _28453_, _12711_);
  and (_28456_, _28454_, _28452_);
  or (_28457_, _28456_, _12720_);
  or (_28458_, _28457_, _28451_);
  or (_28459_, _28267_, _12244_);
  and (_28460_, _28459_, _10969_);
  and (_28461_, _28460_, _28458_);
  nor (_28462_, _14881_, _10969_);
  or (_28463_, _28462_, _06426_);
  or (_28464_, _28463_, _28461_);
  and (_28465_, _28464_, _28273_);
  or (_28467_, _28465_, _06532_);
  nand (_28468_, _14881_, _06532_);
  and (_28469_, _28468_, _27839_);
  and (_28470_, _28469_, _28467_);
  or (_28471_, _28298_, \oc8051_golden_model_1.PSW [7]);
  or (_28472_, _12156_, _10774_);
  and (_28473_, _28472_, _12732_);
  and (_28474_, _28473_, _28471_);
  or (_28475_, _28474_, _12751_);
  or (_28476_, _28475_, _28470_);
  or (_28478_, _28267_, _12749_);
  and (_28479_, _28478_, _11007_);
  and (_28480_, _28479_, _28476_);
  nor (_28481_, _14881_, _11007_);
  or (_28482_, _28481_, _06437_);
  or (_28483_, _28482_, _28480_);
  and (_28484_, _28483_, _28272_);
  or (_28485_, _28484_, _06535_);
  nand (_28486_, _14881_, _06535_);
  and (_28487_, _28486_, _27859_);
  and (_28489_, _28487_, _28485_);
  or (_28490_, _28298_, _10774_);
  or (_28491_, _12156_, \oc8051_golden_model_1.PSW [7]);
  and (_28492_, _28491_, _12239_);
  and (_28493_, _28492_, _28490_);
  or (_28494_, _28493_, _12771_);
  or (_28495_, _28494_, _28489_);
  or (_28496_, _28267_, _12767_);
  and (_28497_, _28496_, _12769_);
  and (_28498_, _28497_, _28495_);
  nor (_28500_, _14881_, _12769_);
  or (_28501_, _28500_, _11111_);
  or (_28502_, _28501_, _28498_);
  and (_28503_, _28502_, _28271_);
  or (_28504_, _28503_, _06543_);
  or (_28505_, _08662_, _12782_);
  and (_28506_, _28505_, _28204_);
  and (_28507_, _28506_, _28504_);
  or (_28508_, _28282_, _25133_);
  or (_28509_, _12281_, _12970_);
  and (_28511_, _28509_, _06436_);
  and (_28512_, _28511_, _28508_);
  or (_28513_, _28512_, _12790_);
  or (_28514_, _28513_, _28507_);
  or (_28515_, _28267_, _12129_);
  and (_28516_, _28515_, _12978_);
  and (_28517_, _28516_, _28514_);
  nor (_28518_, _12978_, _14881_);
  or (_28519_, _28518_, _10472_);
  or (_28520_, _28519_, _28517_);
  and (_28522_, _28520_, _28270_);
  or (_28523_, _28522_, _06290_);
  or (_28524_, _08662_, _06291_);
  and (_28525_, _28524_, _28223_);
  and (_28526_, _28525_, _28523_);
  or (_28527_, _12281_, _25133_);
  or (_28528_, _28282_, _12970_);
  and (_28529_, _28528_, _28527_);
  and (_28530_, _28529_, _06434_);
  or (_28531_, _28530_, _12999_);
  or (_28532_, _28531_, _28526_);
  or (_28533_, _28267_, _12998_);
  and (_28534_, _28533_, _28532_);
  or (_28535_, _28534_, _06559_);
  nand (_28536_, _14881_, _06559_);
  and (_28537_, _28536_, _13005_);
  and (_28538_, _28537_, _28535_);
  nor (_28539_, _28269_, _13005_);
  or (_28540_, _28539_, _06432_);
  or (_28541_, _28540_, _28538_);
  nand (_28544_, _06646_, _06432_);
  and (_28545_, _28544_, _27923_);
  and (_28546_, _28545_, _28541_);
  and (_28547_, _28529_, _05932_);
  or (_28548_, _28547_, _13020_);
  or (_28549_, _28548_, _28546_);
  or (_28550_, _28267_, _13019_);
  and (_28551_, _28550_, _28549_);
  or (_28552_, _28551_, _06566_);
  nand (_28553_, _14881_, _06566_);
  and (_28555_, _28553_, _13027_);
  and (_28556_, _28555_, _28552_);
  nor (_28557_, _28269_, _13027_);
  or (_28558_, _28557_, _06393_);
  or (_28559_, _28558_, _28556_);
  nand (_28560_, _06646_, _06393_);
  and (_28561_, _28560_, _13036_);
  and (_28562_, _28561_, _28559_);
  and (_28563_, _28267_, _13035_);
  or (_28564_, _28563_, _01324_);
  or (_28566_, _28564_, _28562_);
  or (_28567_, _01320_, \oc8051_golden_model_1.PC [10]);
  and (_28568_, _28567_, _42355_);
  and (_42994_, _28568_, _28566_);
  or (_28569_, _09421_, _06291_);
  nor (_28570_, _12121_, \oc8051_golden_model_1.PC [11]);
  nor (_28571_, _28570_, _12122_);
  or (_28572_, _28571_, _12129_);
  or (_28573_, _28571_, _12767_);
  or (_28574_, _28571_, _12749_);
  or (_28576_, _28571_, _12695_);
  or (_28577_, _12151_, _09015_);
  and (_28578_, _12276_, _05972_);
  and (_28579_, _12400_, _12276_);
  not (_28580_, _12282_);
  and (_28581_, _28280_, _28580_);
  and (_28582_, _28581_, _12279_);
  nor (_28583_, _28581_, _12279_);
  or (_28584_, _28583_, _28582_);
  and (_28585_, _28584_, _12398_);
  or (_28587_, _28585_, _06424_);
  or (_28588_, _28587_, _28579_);
  and (_28589_, _12151_, _06345_);
  or (_28590_, _12406_, _12151_);
  or (_28591_, _12420_, _12276_);
  or (_28592_, _28584_, _12418_);
  and (_28593_, _28592_, _06285_);
  and (_28594_, _28593_, _28591_);
  and (_28595_, _12430_, _12151_);
  nor (_28596_, _28296_, _12157_);
  and (_28598_, _28596_, _12154_);
  nor (_28599_, _28596_, _12154_);
  or (_28600_, _28599_, _28598_);
  and (_28601_, _28600_, _25203_);
  or (_28602_, _28601_, _08736_);
  or (_28603_, _28602_, _28595_);
  or (_28604_, _12151_, _07858_);
  or (_28605_, _28571_, _12453_);
  and (_28606_, _28605_, _25213_);
  or (_28607_, _28571_, _28310_);
  or (_28609_, _12151_, _07144_);
  nor (_28610_, _07143_, \oc8051_golden_model_1.PC [11]);
  nand (_28611_, _28610_, _07454_);
  and (_28612_, _28611_, _28609_);
  or (_28613_, _28612_, _06755_);
  and (_28614_, _28613_, _28607_);
  or (_28615_, _28614_, _28606_);
  and (_28616_, _28615_, _28604_);
  or (_28617_, _28616_, _08734_);
  and (_28618_, _28617_, _12457_);
  and (_28620_, _28618_, _28603_);
  or (_28621_, _28620_, _28594_);
  and (_28622_, _28621_, _12409_);
  not (_28623_, _12411_);
  and (_28624_, _28571_, _28623_);
  or (_28625_, _28624_, _12407_);
  or (_28626_, _28625_, _28622_);
  and (_28627_, _28626_, _28590_);
  or (_28628_, _28627_, _26288_);
  or (_28629_, _28571_, _12404_);
  and (_28631_, _28629_, _06346_);
  and (_28632_, _28631_, _28628_);
  or (_28633_, _28632_, _28589_);
  and (_28634_, _28633_, _12468_);
  and (_28635_, _28571_, _12473_);
  or (_28636_, _28635_, _12478_);
  or (_28637_, _28636_, _28634_);
  or (_28638_, _12477_, _12151_);
  and (_28639_, _28638_, _28637_);
  or (_28640_, _28639_, _12485_);
  and (_28642_, _12519_, _12276_);
  and (_28643_, _28584_, _25019_);
  or (_28644_, _28643_, _28642_);
  or (_28645_, _28644_, _12484_);
  and (_28646_, _28645_, _28640_);
  or (_28647_, _28646_, _06423_);
  and (_28648_, _28647_, _28588_);
  and (_28649_, _28648_, _06420_);
  and (_28650_, _28584_, _25279_);
  and (_28651_, _12540_, _12276_);
  or (_28653_, _28651_, _28650_);
  and (_28654_, _28653_, _06347_);
  or (_28655_, _28584_, _12559_);
  or (_28656_, _12560_, _12276_);
  and (_28657_, _28656_, _06419_);
  and (_28658_, _28657_, _28655_);
  or (_28659_, _28658_, _28654_);
  or (_28660_, _28659_, _28649_);
  and (_28661_, _28660_, _12255_);
  nand (_28662_, _28571_, _12254_);
  nand (_28664_, _28662_, _12579_);
  or (_28665_, _28664_, _28661_);
  or (_28666_, _12579_, _12151_);
  and (_28667_, _28666_, _12585_);
  and (_28668_, _28667_, _28665_);
  and (_28669_, _28571_, _12589_);
  or (_28670_, _28669_, _12592_);
  or (_28671_, _28670_, _28668_);
  or (_28672_, _12591_, _12151_);
  and (_28673_, _28672_, _12595_);
  and (_28675_, _28673_, _28671_);
  and (_28676_, _28571_, _12601_);
  or (_28677_, _28676_, _12600_);
  or (_28678_, _28677_, _28675_);
  or (_28679_, _12151_, _12599_);
  and (_28680_, _28679_, _05940_);
  and (_28681_, _28680_, _28678_);
  nand (_28682_, _28571_, _05976_);
  nand (_28683_, _28682_, _12609_);
  or (_28684_, _28683_, _28681_);
  or (_28686_, _12609_, _12151_);
  and (_28687_, _28686_, _06396_);
  and (_28688_, _28687_, _28684_);
  nand (_28689_, _12276_, _06395_);
  nand (_28690_, _28689_, _06261_);
  or (_28691_, _28690_, _28688_);
  or (_28692_, _12151_, _06261_);
  and (_28693_, _28692_, _06251_);
  and (_28694_, _28693_, _28691_);
  or (_28695_, _28694_, _28578_);
  and (_28697_, _28695_, _12252_);
  and (_28698_, _28571_, _12626_);
  or (_28699_, _28698_, _12625_);
  or (_28700_, _28699_, _28697_);
  or (_28701_, _12624_, _12151_);
  and (_28702_, _28701_, _12631_);
  and (_28703_, _28702_, _28700_);
  and (_28704_, _28600_, _12630_);
  or (_28705_, _28704_, _09016_);
  or (_28706_, _28705_, _28703_);
  and (_28708_, _28706_, _28577_);
  or (_28709_, _28708_, _06215_);
  or (_28710_, _12276_, _06216_);
  and (_28711_, _28710_, _10892_);
  and (_28712_, _28711_, _28709_);
  and (_28713_, _12151_, _10891_);
  or (_28714_, _28713_, _28712_);
  and (_28715_, _28714_, _25380_);
  or (_28716_, _12671_, \oc8051_golden_model_1.DPH [3]);
  nor (_28717_, _12672_, _25380_);
  and (_28719_, _28717_, _28716_);
  or (_28720_, _28719_, _12681_);
  or (_28721_, _28720_, _28715_);
  or (_28722_, _12680_, _12151_);
  and (_28723_, _28722_, _12685_);
  and (_28724_, _28723_, _28721_);
  or (_28725_, _28600_, _11327_);
  or (_28726_, _12151_, _12248_);
  and (_28727_, _28726_, _12247_);
  and (_28728_, _28727_, _28725_);
  or (_28730_, _28728_, _12697_);
  or (_28731_, _28730_, _28724_);
  and (_28732_, _28731_, _28576_);
  or (_28733_, _28732_, _12700_);
  or (_28734_, _12699_, _12151_);
  and (_28735_, _28734_, _09025_);
  and (_28736_, _28735_, _28733_);
  nand (_28737_, _12276_, _06398_);
  nand (_28738_, _28737_, _12708_);
  or (_28739_, _28738_, _28736_);
  or (_28741_, _12708_, _12151_);
  and (_28742_, _28741_, _12712_);
  and (_28743_, _28742_, _28739_);
  or (_28744_, _28600_, _12248_);
  or (_28745_, _12151_, _11327_);
  and (_28746_, _28745_, _12711_);
  and (_28747_, _28746_, _28744_);
  or (_28748_, _28747_, _28743_);
  and (_28749_, _28748_, _12244_);
  and (_28750_, _28571_, _12720_);
  or (_28752_, _28750_, _10970_);
  or (_28753_, _28752_, _28749_);
  or (_28754_, _12151_, _10969_);
  and (_28755_, _28754_, _07219_);
  and (_28756_, _28755_, _28753_);
  nand (_28757_, _12276_, _06426_);
  nand (_28758_, _28757_, _12729_);
  or (_28759_, _28758_, _28756_);
  or (_28760_, _12729_, _12151_);
  and (_28761_, _28760_, _12733_);
  and (_28763_, _28761_, _28759_);
  or (_28764_, _28600_, \oc8051_golden_model_1.PSW [7]);
  or (_28765_, _12151_, _10774_);
  and (_28766_, _28765_, _12732_);
  and (_28767_, _28766_, _28764_);
  or (_28768_, _28767_, _12751_);
  or (_28769_, _28768_, _28763_);
  and (_28770_, _28769_, _28574_);
  or (_28771_, _28770_, _11008_);
  or (_28772_, _12151_, _11007_);
  and (_28774_, _28772_, _07229_);
  and (_28775_, _28774_, _28771_);
  nand (_28776_, _12276_, _06437_);
  nand (_28777_, _28776_, _12759_);
  or (_28778_, _28777_, _28775_);
  or (_28779_, _12759_, _12151_);
  and (_28780_, _28779_, _12762_);
  and (_28781_, _28780_, _28778_);
  or (_28782_, _28600_, _10774_);
  or (_28783_, _12151_, \oc8051_golden_model_1.PSW [7]);
  and (_28785_, _28783_, _12239_);
  and (_28786_, _28785_, _28782_);
  or (_28787_, _28786_, _12771_);
  or (_28788_, _28787_, _28781_);
  and (_28789_, _28788_, _28573_);
  or (_28790_, _28789_, _12770_);
  or (_28791_, _12151_, _12769_);
  and (_28792_, _28791_, _12775_);
  and (_28793_, _28792_, _28790_);
  and (_28794_, _28571_, _11111_);
  or (_28796_, _28794_, _06543_);
  or (_28797_, _28796_, _28793_);
  or (_28798_, _09421_, _12782_);
  and (_28799_, _28798_, _28797_);
  or (_28800_, _28799_, _06011_);
  or (_28801_, _12151_, _09057_);
  and (_28802_, _28801_, _12786_);
  and (_28803_, _28802_, _28800_);
  or (_28804_, _28584_, _25133_);
  or (_28805_, _12276_, _12970_);
  and (_28807_, _28805_, _06436_);
  and (_28808_, _28807_, _28804_);
  or (_28809_, _28808_, _12790_);
  or (_28810_, _28809_, _28803_);
  and (_28811_, _28810_, _28572_);
  or (_28812_, _28811_, _12979_);
  or (_28813_, _12978_, _12151_);
  and (_28814_, _28813_, _12981_);
  and (_28815_, _28814_, _28812_);
  and (_28816_, _28571_, _10472_);
  or (_28818_, _28816_, _06290_);
  or (_28819_, _28818_, _28815_);
  and (_28820_, _28819_, _28569_);
  or (_28821_, _28820_, _05994_);
  or (_28822_, _12151_, _25143_);
  and (_28823_, _28822_, _06435_);
  and (_28824_, _28823_, _28821_);
  or (_28825_, _28584_, _12970_);
  or (_28826_, _12276_, _25133_);
  and (_28827_, _28826_, _28825_);
  and (_28829_, _28827_, _06434_);
  or (_28830_, _28829_, _12999_);
  or (_28831_, _28830_, _28824_);
  or (_28832_, _28571_, _12998_);
  and (_28833_, _28832_, _07240_);
  and (_28834_, _28833_, _28831_);
  nand (_28835_, _12151_, _06559_);
  nand (_28836_, _28835_, _13005_);
  or (_28837_, _28836_, _28834_);
  or (_28838_, _28571_, _13005_);
  and (_28840_, _28838_, _06433_);
  and (_28841_, _28840_, _28837_);
  nor (_28842_, _06433_, _06212_);
  or (_28843_, _28842_, _05991_);
  or (_28844_, _28843_, _28841_);
  or (_28845_, _12151_, _14666_);
  and (_28846_, _28845_, _05933_);
  and (_28847_, _28846_, _28844_);
  and (_28848_, _28827_, _05932_);
  or (_28849_, _28848_, _13020_);
  or (_28851_, _28849_, _28847_);
  or (_28852_, _28571_, _13019_);
  and (_28853_, _28852_, _06570_);
  and (_28854_, _28853_, _28851_);
  nand (_28855_, _12151_, _06566_);
  nand (_28856_, _28855_, _13027_);
  or (_28857_, _28856_, _28854_);
  or (_28858_, _28571_, _13027_);
  and (_28859_, _28858_, _13030_);
  and (_28860_, _28859_, _28857_);
  nor (_28862_, _13030_, _06212_);
  or (_28863_, _28862_, _05989_);
  or (_28864_, _28863_, _28860_);
  or (_28865_, _12151_, _05990_);
  and (_28866_, _28865_, _13039_);
  and (_28867_, _28866_, _28864_);
  and (_28868_, _28571_, _13035_);
  or (_28869_, _28868_, _01324_);
  or (_28870_, _28869_, _28867_);
  or (_28871_, _01320_, \oc8051_golden_model_1.PC [11]);
  and (_28873_, _28871_, _42355_);
  and (_42995_, _28873_, _28870_);
  and (_28874_, _01324_, \oc8051_golden_model_1.PC [12]);
  nand (_28875_, _06961_, _06393_);
  and (_28876_, _28875_, _05990_);
  nor (_28877_, _12122_, \oc8051_golden_model_1.PC [12]);
  nor (_28878_, _28877_, _12123_);
  or (_28879_, _28878_, _12981_);
  nor (_28880_, _12759_, _15304_);
  nor (_28881_, _12729_, _15304_);
  nor (_28883_, _12708_, _15304_);
  nand (_28884_, _15304_, _06345_);
  or (_28885_, _12355_, _12353_);
  and (_28886_, _28885_, _12356_);
  or (_28887_, _28886_, _12418_);
  or (_28888_, _12420_, _12273_);
  and (_28889_, _28888_, _06285_);
  and (_28890_, _28889_, _28887_);
  and (_28891_, _12430_, _12148_);
  or (_28892_, _12225_, _12223_);
  and (_28894_, _28892_, _12226_);
  and (_28895_, _28894_, _12432_);
  or (_28896_, _28895_, _28891_);
  or (_28897_, _28896_, _08736_);
  or (_28898_, _28878_, _12453_);
  or (_28899_, _12448_, _12148_);
  and (_28900_, _28899_, _28898_);
  or (_28901_, _28900_, _24979_);
  not (_28902_, _28310_);
  and (_28903_, _28878_, _28902_);
  nand (_28904_, _15304_, _07143_);
  and (_28905_, _28904_, _06756_);
  and (_28906_, _07454_, \oc8051_golden_model_1.PC [12]);
  or (_28907_, _28906_, _07143_);
  and (_28908_, _28907_, _28905_);
  or (_28909_, _28908_, _07152_);
  or (_28910_, _28909_, _28903_);
  and (_28911_, _28910_, _28901_);
  or (_28912_, _28911_, _08734_);
  and (_28913_, _28912_, _12457_);
  and (_28916_, _28913_, _28897_);
  or (_28917_, _28916_, _28890_);
  and (_28918_, _28917_, _12409_);
  and (_28919_, _28878_, _28623_);
  or (_28920_, _28919_, _12407_);
  or (_28921_, _28920_, _28918_);
  or (_28922_, _12406_, _12148_);
  and (_28923_, _28922_, _12404_);
  and (_28924_, _28923_, _28921_);
  and (_28925_, _28878_, _26288_);
  or (_28927_, _28925_, _06345_);
  or (_28928_, _28927_, _28924_);
  and (_28929_, _28928_, _28884_);
  or (_28930_, _28929_, _12473_);
  or (_28931_, _28878_, _12468_);
  and (_28932_, _28931_, _12477_);
  and (_28933_, _28932_, _28930_);
  or (_28934_, _12477_, _15304_);
  nand (_28935_, _28934_, _12484_);
  or (_28936_, _28935_, _28933_);
  and (_28938_, _12519_, _12273_);
  and (_28939_, _28886_, _25019_);
  or (_28940_, _28939_, _28938_);
  or (_28941_, _28940_, _12484_);
  and (_28942_, _28941_, _06424_);
  and (_28943_, _28942_, _28936_);
  or (_28944_, _12398_, _12273_);
  or (_28945_, _28886_, _12400_);
  and (_28946_, _28945_, _06423_);
  and (_28947_, _28946_, _28944_);
  or (_28949_, _28947_, _28943_);
  and (_28950_, _28949_, _06420_);
  or (_28951_, _28886_, _12559_);
  or (_28952_, _12560_, _12273_);
  and (_28953_, _28952_, _06419_);
  and (_28954_, _28953_, _28951_);
  or (_28955_, _28954_, _12254_);
  or (_28956_, _28886_, _12540_);
  or (_28957_, _25279_, _12273_);
  and (_28958_, _28957_, _06347_);
  and (_28960_, _28958_, _28956_);
  or (_28961_, _28960_, _28955_);
  or (_28962_, _28961_, _28950_);
  or (_28963_, _28878_, _12255_);
  and (_28964_, _28963_, _12579_);
  and (_28965_, _28964_, _28962_);
  nor (_28966_, _12579_, _15304_);
  or (_28967_, _28966_, _12589_);
  or (_28968_, _28967_, _28965_);
  or (_28969_, _28878_, _12585_);
  and (_28971_, _28969_, _12591_);
  and (_28972_, _28971_, _28968_);
  or (_28973_, _12591_, _15304_);
  nand (_28974_, _28973_, _12595_);
  or (_28975_, _28974_, _28972_);
  or (_28976_, _28878_, _12595_);
  and (_28977_, _28976_, _12599_);
  and (_28978_, _28977_, _28975_);
  nor (_28979_, _15304_, _12599_);
  or (_28980_, _28979_, _05976_);
  or (_28982_, _28980_, _28978_);
  or (_28983_, _28878_, _05940_);
  and (_28984_, _28983_, _12609_);
  and (_28985_, _28984_, _28982_);
  nor (_28986_, _12609_, _15304_);
  or (_28987_, _28986_, _06395_);
  or (_28988_, _28987_, _28985_);
  or (_28989_, _12273_, _06396_);
  and (_28990_, _28989_, _06261_);
  and (_28991_, _28990_, _28988_);
  nor (_28993_, _15304_, _06261_);
  or (_28994_, _28993_, _05972_);
  or (_28995_, _28994_, _28991_);
  or (_28996_, _12273_, _06251_);
  and (_28997_, _28996_, _12252_);
  and (_28998_, _28997_, _28995_);
  and (_28999_, _28878_, _12626_);
  or (_29000_, _28999_, _12625_);
  or (_29001_, _29000_, _28998_);
  or (_29002_, _12624_, _12148_);
  and (_29004_, _29002_, _12631_);
  and (_29005_, _29004_, _29001_);
  and (_29006_, _28894_, _12630_);
  or (_29007_, _29006_, _29005_);
  and (_29008_, _29007_, _09015_);
  nor (_29009_, _15304_, _09015_);
  or (_29010_, _29009_, _06215_);
  or (_29011_, _29010_, _29008_);
  or (_29012_, _12273_, _06216_);
  and (_29013_, _29012_, _10892_);
  and (_29015_, _29013_, _29011_);
  and (_29016_, _12148_, _10891_);
  or (_29017_, _29016_, _12644_);
  or (_29018_, _29017_, _29015_);
  nor (_29019_, _12672_, \oc8051_golden_model_1.DPH [4]);
  nor (_29020_, _29019_, _12673_);
  or (_29021_, _29020_, _25380_);
  and (_29022_, _29021_, _29018_);
  or (_29023_, _29022_, _12681_);
  or (_29024_, _12680_, _12148_);
  and (_29026_, _29024_, _12685_);
  and (_29027_, _29026_, _29023_);
  or (_29028_, _28894_, _11327_);
  or (_29029_, _12148_, _12248_);
  and (_29030_, _29029_, _12247_);
  and (_29031_, _29030_, _29028_);
  or (_29032_, _29031_, _12697_);
  or (_29033_, _29032_, _29027_);
  or (_29034_, _28878_, _12695_);
  and (_29035_, _29034_, _12699_);
  and (_29037_, _29035_, _29033_);
  nor (_29038_, _12699_, _15304_);
  or (_29039_, _29038_, _06398_);
  or (_29040_, _29039_, _29037_);
  or (_29041_, _12273_, _09025_);
  and (_29042_, _29041_, _12708_);
  and (_29043_, _29042_, _29040_);
  or (_29044_, _29043_, _28883_);
  and (_29045_, _29044_, _12712_);
  or (_29046_, _28894_, _12248_);
  or (_29048_, _12148_, _11327_);
  and (_29049_, _29048_, _12711_);
  and (_29050_, _29049_, _29046_);
  or (_29051_, _29050_, _12720_);
  or (_29052_, _29051_, _29045_);
  or (_29053_, _28878_, _12244_);
  and (_29054_, _29053_, _10969_);
  and (_29055_, _29054_, _29052_);
  nor (_29056_, _15304_, _10969_);
  or (_29057_, _29056_, _06426_);
  or (_29059_, _29057_, _29055_);
  or (_29060_, _12273_, _07219_);
  and (_29061_, _29060_, _12729_);
  and (_29062_, _29061_, _29059_);
  or (_29063_, _29062_, _28881_);
  and (_29064_, _29063_, _12733_);
  or (_29065_, _28894_, \oc8051_golden_model_1.PSW [7]);
  or (_29066_, _12148_, _10774_);
  and (_29067_, _29066_, _12732_);
  and (_29068_, _29067_, _29065_);
  or (_29070_, _29068_, _12751_);
  or (_29071_, _29070_, _29064_);
  or (_29072_, _28878_, _12749_);
  and (_29073_, _29072_, _11007_);
  and (_29074_, _29073_, _29071_);
  nor (_29075_, _15304_, _11007_);
  or (_29076_, _29075_, _06437_);
  or (_29077_, _29076_, _29074_);
  or (_29078_, _12273_, _07229_);
  and (_29079_, _29078_, _12759_);
  and (_29081_, _29079_, _29077_);
  or (_29082_, _29081_, _28880_);
  and (_29083_, _29082_, _12762_);
  or (_29084_, _28894_, _10774_);
  or (_29085_, _12148_, \oc8051_golden_model_1.PSW [7]);
  and (_29086_, _29085_, _12239_);
  and (_29087_, _29086_, _29084_);
  or (_29088_, _29087_, _12771_);
  or (_29089_, _29088_, _29083_);
  or (_29090_, _28878_, _12767_);
  and (_29092_, _29090_, _12769_);
  and (_29093_, _29092_, _29089_);
  nor (_29094_, _15304_, _12769_);
  or (_29095_, _29094_, _11111_);
  or (_29096_, _29095_, _29093_);
  or (_29097_, _28878_, _12775_);
  and (_29098_, _29097_, _12782_);
  and (_29099_, _29098_, _29096_);
  and (_29100_, _09420_, _06543_);
  or (_29101_, _29100_, _06011_);
  or (_29103_, _29101_, _29099_);
  nand (_29104_, _15304_, _06011_);
  and (_29105_, _29104_, _12786_);
  and (_29106_, _29105_, _29103_);
  or (_29107_, _28886_, _25133_);
  or (_29108_, _12273_, _12970_);
  and (_29109_, _29108_, _06436_);
  and (_29110_, _29109_, _29107_);
  or (_29111_, _29110_, _12790_);
  or (_29112_, _29111_, _29106_);
  or (_29114_, _28878_, _12129_);
  and (_29115_, _29114_, _12978_);
  and (_29116_, _29115_, _29112_);
  nor (_29117_, _12978_, _15304_);
  or (_29118_, _29117_, _10472_);
  or (_29119_, _29118_, _29116_);
  and (_29120_, _29119_, _28879_);
  or (_29121_, _29120_, _06290_);
  or (_29122_, _09420_, _06291_);
  and (_29123_, _29122_, _25143_);
  and (_29125_, _29123_, _29121_);
  and (_29126_, _12148_, _05994_);
  or (_29127_, _29126_, _06434_);
  or (_29128_, _29127_, _29125_);
  or (_29129_, _28886_, _12970_);
  or (_29130_, _12273_, _25133_);
  and (_29131_, _29130_, _29129_);
  or (_29132_, _29131_, _06435_);
  and (_29133_, _29132_, _29128_);
  or (_29134_, _29133_, _12999_);
  or (_29136_, _28878_, _12998_);
  and (_29137_, _29136_, _29134_);
  or (_29138_, _29137_, _06559_);
  nand (_29139_, _15304_, _06559_);
  and (_29140_, _29139_, _13005_);
  and (_29141_, _29140_, _29138_);
  and (_29142_, _28878_, _26914_);
  or (_29143_, _29142_, _06432_);
  or (_29144_, _29143_, _29141_);
  nand (_29145_, _06961_, _06432_);
  and (_29147_, _29145_, _14666_);
  and (_29148_, _29147_, _29144_);
  and (_29149_, _12148_, _05991_);
  or (_29150_, _29149_, _05932_);
  or (_29151_, _29150_, _29148_);
  or (_29152_, _29131_, _05933_);
  and (_29153_, _29152_, _13019_);
  and (_29154_, _29153_, _29151_);
  and (_29155_, _28878_, _13020_);
  or (_29156_, _29155_, _06566_);
  or (_29158_, _29156_, _29154_);
  nand (_29159_, _15304_, _06566_);
  and (_29160_, _29159_, _13027_);
  and (_29161_, _29160_, _29158_);
  and (_29162_, _28878_, _26930_);
  or (_29163_, _29162_, _06393_);
  or (_29164_, _29163_, _29161_);
  and (_29165_, _29164_, _28876_);
  and (_29166_, _12148_, _05989_);
  or (_29167_, _29166_, _13035_);
  or (_29169_, _29167_, _29165_);
  or (_29170_, _28878_, _13039_);
  and (_29171_, _29170_, _01320_);
  and (_29172_, _29171_, _29169_);
  or (_29173_, _29172_, _28874_);
  and (_42996_, _29173_, _42355_);
  and (_29174_, _01324_, \oc8051_golden_model_1.PC [13]);
  nor (_29175_, _12123_, \oc8051_golden_model_1.PC [13]);
  nor (_29176_, _29175_, _12124_);
  or (_29177_, _29176_, _13027_);
  or (_29179_, _09419_, _06291_);
  or (_29180_, _29176_, _12129_);
  or (_29181_, _29176_, _12767_);
  or (_29182_, _29176_, _12749_);
  or (_29183_, _12146_, _12145_);
  not (_29184_, _29183_);
  nor (_29185_, _29184_, _12227_);
  and (_29186_, _29184_, _12227_);
  or (_29187_, _29186_, _29185_);
  or (_29188_, _29187_, _12248_);
  or (_29190_, _12144_, _11327_);
  and (_29191_, _29190_, _12711_);
  and (_29192_, _29191_, _29188_);
  or (_29193_, _29176_, _12695_);
  or (_29194_, _12144_, _09015_);
  and (_29195_, _12269_, _05972_);
  and (_29196_, _12400_, _12269_);
  or (_29197_, _12271_, _12270_);
  not (_29198_, _29197_);
  nor (_29199_, _29198_, _12357_);
  and (_29201_, _29198_, _12357_);
  or (_29202_, _29201_, _29199_);
  and (_29203_, _29202_, _12398_);
  or (_29204_, _29203_, _29196_);
  or (_29205_, _29204_, _06424_);
  and (_29206_, _12144_, _06345_);
  or (_29207_, _12406_, _12144_);
  or (_29208_, _29202_, _12418_);
  or (_29209_, _12420_, _12269_);
  and (_29210_, _29209_, _06285_);
  and (_29212_, _29210_, _29208_);
  and (_29213_, _12430_, _12144_);
  and (_29214_, _29187_, _25203_);
  or (_29215_, _29214_, _08736_);
  or (_29216_, _29215_, _29213_);
  or (_29217_, _29176_, _28310_);
  or (_29218_, _12144_, _07858_);
  or (_29219_, _12144_, _07144_);
  nor (_29220_, _07143_, \oc8051_golden_model_1.PC [13]);
  nand (_29221_, _29220_, _07454_);
  and (_29223_, _29221_, _29219_);
  nand (_29224_, _24979_, _06756_);
  or (_29225_, _29224_, _29223_);
  and (_29226_, _29225_, _29218_);
  and (_29227_, _29226_, _29217_);
  or (_29228_, _29227_, _08734_);
  and (_29229_, _29228_, _12457_);
  and (_29230_, _29229_, _29216_);
  or (_29231_, _29230_, _29212_);
  and (_29232_, _29231_, _12409_);
  and (_29234_, _29176_, _28623_);
  or (_29235_, _29234_, _12407_);
  or (_29236_, _29235_, _29232_);
  and (_29237_, _29236_, _29207_);
  or (_29238_, _29237_, _26288_);
  or (_29239_, _29176_, _12404_);
  and (_29240_, _29239_, _06346_);
  and (_29241_, _29240_, _29238_);
  or (_29242_, _29241_, _29206_);
  and (_29243_, _29242_, _12468_);
  and (_29245_, _29176_, _12473_);
  or (_29246_, _29245_, _12478_);
  or (_29247_, _29246_, _29243_);
  or (_29248_, _12477_, _12144_);
  and (_29249_, _29248_, _12484_);
  and (_29250_, _29249_, _29247_);
  or (_29251_, _25019_, _12269_);
  or (_29252_, _29202_, _12519_);
  and (_29253_, _29252_, _12485_);
  and (_29254_, _29253_, _29251_);
  or (_29256_, _29254_, _06423_);
  or (_29257_, _29256_, _29250_);
  and (_29258_, _29257_, _29205_);
  or (_29259_, _29258_, _06347_);
  and (_29260_, _29202_, _25279_);
  and (_29261_, _12540_, _12269_);
  or (_29262_, _29261_, _14105_);
  or (_29263_, _29262_, _29260_);
  and (_29264_, _29263_, _12528_);
  and (_29265_, _29264_, _29259_);
  or (_29267_, _29202_, _12559_);
  or (_29268_, _12560_, _12269_);
  and (_29269_, _29268_, _06419_);
  and (_29270_, _29269_, _29267_);
  or (_29271_, _29270_, _29265_);
  and (_29272_, _29271_, _12255_);
  nand (_29273_, _29176_, _12254_);
  nand (_29274_, _29273_, _12579_);
  or (_29275_, _29274_, _29272_);
  or (_29276_, _12579_, _12144_);
  and (_29278_, _29276_, _12585_);
  and (_29279_, _29278_, _29275_);
  and (_29280_, _29176_, _12589_);
  or (_29281_, _29280_, _12592_);
  or (_29282_, _29281_, _29279_);
  or (_29283_, _12591_, _12144_);
  and (_29284_, _29283_, _12595_);
  and (_29285_, _29284_, _29282_);
  and (_29286_, _29176_, _12601_);
  or (_29287_, _29286_, _12600_);
  or (_29289_, _29287_, _29285_);
  or (_29290_, _12144_, _12599_);
  and (_29291_, _29290_, _05940_);
  and (_29292_, _29291_, _29289_);
  nand (_29293_, _29176_, _05976_);
  nand (_29294_, _29293_, _12609_);
  or (_29295_, _29294_, _29292_);
  or (_29296_, _12609_, _12144_);
  and (_29297_, _29296_, _06396_);
  and (_29298_, _29297_, _29295_);
  nand (_29300_, _12269_, _06395_);
  nand (_29301_, _29300_, _06261_);
  or (_29302_, _29301_, _29298_);
  or (_29303_, _12144_, _06261_);
  and (_29304_, _29303_, _06251_);
  and (_29305_, _29304_, _29302_);
  or (_29306_, _29305_, _29195_);
  and (_29307_, _29306_, _12252_);
  and (_29308_, _29176_, _12626_);
  or (_29309_, _29308_, _12625_);
  or (_29311_, _29309_, _29307_);
  or (_29312_, _12624_, _12144_);
  and (_29313_, _29312_, _12631_);
  and (_29314_, _29313_, _29311_);
  and (_29315_, _29187_, _12630_);
  or (_29316_, _29315_, _09016_);
  or (_29317_, _29316_, _29314_);
  and (_29318_, _29317_, _29194_);
  or (_29319_, _29318_, _06215_);
  or (_29320_, _12269_, _06216_);
  and (_29322_, _29320_, _10892_);
  and (_29323_, _29322_, _29319_);
  and (_29324_, _12144_, _10891_);
  or (_29325_, _29324_, _29323_);
  and (_29326_, _29325_, _25380_);
  or (_29327_, _12673_, \oc8051_golden_model_1.DPH [5]);
  nor (_29328_, _12674_, _25380_);
  and (_29329_, _29328_, _29327_);
  or (_29330_, _29329_, _12681_);
  or (_29331_, _29330_, _29326_);
  or (_29333_, _12680_, _12144_);
  and (_29334_, _29333_, _12685_);
  and (_29335_, _29334_, _29331_);
  or (_29336_, _29187_, _11327_);
  or (_29337_, _12144_, _12248_);
  and (_29338_, _29337_, _12247_);
  and (_29339_, _29338_, _29336_);
  or (_29340_, _29339_, _12697_);
  or (_29341_, _29340_, _29335_);
  and (_29342_, _29341_, _29193_);
  or (_29344_, _29342_, _12700_);
  or (_29345_, _12699_, _12144_);
  and (_29346_, _29345_, _09025_);
  and (_29347_, _29346_, _29344_);
  nand (_29348_, _12269_, _06398_);
  nand (_29349_, _29348_, _12708_);
  or (_29350_, _29349_, _29347_);
  or (_29351_, _12708_, _12144_);
  and (_29352_, _29351_, _12712_);
  and (_29353_, _29352_, _29350_);
  or (_29355_, _29353_, _29192_);
  and (_29356_, _29355_, _12244_);
  and (_29357_, _29176_, _12720_);
  or (_29358_, _29357_, _10970_);
  or (_29359_, _29358_, _29356_);
  or (_29360_, _12144_, _10969_);
  and (_29361_, _29360_, _07219_);
  and (_29362_, _29361_, _29359_);
  nand (_29363_, _12269_, _06426_);
  nand (_29364_, _29363_, _12729_);
  or (_29366_, _29364_, _29362_);
  or (_29367_, _12729_, _12144_);
  and (_29368_, _29367_, _12733_);
  and (_29369_, _29368_, _29366_);
  or (_29370_, _29187_, \oc8051_golden_model_1.PSW [7]);
  or (_29371_, _12144_, _10774_);
  and (_29372_, _29371_, _12732_);
  and (_29373_, _29372_, _29370_);
  or (_29374_, _29373_, _12751_);
  or (_29375_, _29374_, _29369_);
  and (_29377_, _29375_, _29182_);
  or (_29378_, _29377_, _11008_);
  or (_29379_, _12144_, _11007_);
  and (_29380_, _29379_, _07229_);
  and (_29381_, _29380_, _29378_);
  nand (_29382_, _12269_, _06437_);
  nand (_29383_, _29382_, _12759_);
  or (_29384_, _29383_, _29381_);
  or (_29385_, _12759_, _12144_);
  and (_29386_, _29385_, _12762_);
  and (_29388_, _29386_, _29384_);
  or (_29389_, _29187_, _10774_);
  or (_29390_, _12144_, \oc8051_golden_model_1.PSW [7]);
  and (_29391_, _29390_, _12239_);
  and (_29392_, _29391_, _29389_);
  or (_29393_, _29392_, _12771_);
  or (_29394_, _29393_, _29388_);
  and (_29395_, _29394_, _29181_);
  or (_29396_, _29395_, _12770_);
  or (_29397_, _12144_, _12769_);
  and (_29399_, _29397_, _12775_);
  and (_29400_, _29399_, _29396_);
  and (_29401_, _29176_, _11111_);
  or (_29402_, _29401_, _06543_);
  or (_29403_, _29402_, _29400_);
  or (_29404_, _09419_, _12782_);
  and (_29405_, _29404_, _29403_);
  or (_29406_, _29405_, _06011_);
  or (_29407_, _12144_, _09057_);
  and (_29408_, _29407_, _12786_);
  and (_29410_, _29408_, _29406_);
  or (_29411_, _29202_, _25133_);
  or (_29412_, _12269_, _12970_);
  and (_29413_, _29412_, _06436_);
  and (_29414_, _29413_, _29411_);
  or (_29415_, _29414_, _12790_);
  or (_29416_, _29415_, _29410_);
  and (_29417_, _29416_, _29180_);
  or (_29418_, _29417_, _12979_);
  or (_29419_, _12978_, _12144_);
  and (_29421_, _29419_, _12981_);
  and (_29422_, _29421_, _29418_);
  and (_29423_, _29176_, _10472_);
  or (_29424_, _29423_, _06290_);
  or (_29425_, _29424_, _29422_);
  and (_29426_, _29425_, _29179_);
  or (_29427_, _29426_, _05994_);
  or (_29428_, _12144_, _25143_);
  and (_29429_, _29428_, _06435_);
  and (_29430_, _29429_, _29427_);
  or (_29431_, _12269_, _25133_);
  or (_29432_, _29202_, _12970_);
  and (_29433_, _29432_, _29431_);
  and (_29434_, _29433_, _06434_);
  or (_29435_, _29434_, _12999_);
  or (_29436_, _29435_, _29430_);
  or (_29437_, _29176_, _12998_);
  and (_29438_, _29437_, _07240_);
  and (_29439_, _29438_, _29436_);
  nand (_29440_, _12144_, _06559_);
  nand (_29443_, _29440_, _13005_);
  or (_29444_, _29443_, _29439_);
  or (_29445_, _29176_, _13005_);
  and (_29446_, _29445_, _06433_);
  and (_29447_, _29446_, _29444_);
  nor (_29448_, _06604_, _06433_);
  or (_29449_, _29448_, _05991_);
  or (_29450_, _29449_, _29447_);
  or (_29451_, _12144_, _14666_);
  and (_29452_, _29451_, _05933_);
  and (_29454_, _29452_, _29450_);
  and (_29455_, _29433_, _05932_);
  or (_29456_, _29455_, _13020_);
  or (_29457_, _29456_, _29454_);
  or (_29458_, _29176_, _13019_);
  and (_29459_, _29458_, _06570_);
  and (_29460_, _29459_, _29457_);
  nand (_29461_, _12144_, _06566_);
  nand (_29462_, _29461_, _13027_);
  or (_29463_, _29462_, _29460_);
  and (_29465_, _29463_, _29177_);
  or (_29466_, _29465_, _06393_);
  nand (_29467_, _06604_, _06393_);
  and (_29468_, _29467_, _05990_);
  and (_29469_, _29468_, _29466_);
  and (_29470_, _12144_, _05989_);
  or (_29471_, _29470_, _13035_);
  or (_29472_, _29471_, _29469_);
  or (_29473_, _29176_, _13039_);
  and (_29474_, _29473_, _01320_);
  and (_29476_, _29474_, _29472_);
  or (_29477_, _29476_, _29174_);
  and (_42998_, _29477_, _42355_);
  or (_29478_, _12124_, \oc8051_golden_model_1.PC [14]);
  and (_29479_, _29478_, _12125_);
  or (_29480_, _29479_, _12981_);
  not (_29481_, _12139_);
  nor (_29482_, _12759_, _29481_);
  nor (_29483_, _12729_, _29481_);
  nor (_29484_, _12708_, _29481_);
  nor (_29486_, _12680_, _29481_);
  and (_29487_, _12400_, _12264_);
  or (_29488_, _12359_, _12267_);
  and (_29489_, _29488_, _12360_);
  and (_29490_, _29489_, _12398_);
  or (_29491_, _29490_, _06424_);
  or (_29492_, _29491_, _29487_);
  and (_29493_, _12519_, _12264_);
  and (_29494_, _29489_, _25019_);
  or (_29495_, _29494_, _29493_);
  or (_29497_, _29495_, _12484_);
  or (_29498_, _12139_, _06346_);
  or (_29499_, _29489_, _12418_);
  or (_29500_, _12420_, _12264_);
  and (_29501_, _29500_, _06285_);
  and (_29502_, _29501_, _29499_);
  and (_29503_, _12430_, _12139_);
  or (_29504_, _12229_, _12142_);
  and (_29505_, _29504_, _12230_);
  and (_29506_, _29505_, _12432_);
  or (_29508_, _29506_, _29503_);
  or (_29509_, _29508_, _08736_);
  or (_29510_, _29479_, _12453_);
  or (_29511_, _12448_, _12139_);
  and (_29512_, _29511_, _29510_);
  or (_29513_, _29512_, _24979_);
  and (_29514_, _29479_, _28902_);
  nand (_29515_, _29481_, _07143_);
  and (_29516_, _29515_, _06756_);
  and (_29517_, _07454_, \oc8051_golden_model_1.PC [14]);
  or (_29519_, _29517_, _07143_);
  and (_29520_, _29519_, _29516_);
  or (_29521_, _29520_, _07152_);
  or (_29522_, _29521_, _29514_);
  and (_29523_, _29522_, _29513_);
  or (_29524_, _29523_, _08734_);
  and (_29525_, _29524_, _12457_);
  and (_29526_, _29525_, _29509_);
  or (_29527_, _29526_, _29502_);
  and (_29528_, _29527_, _12409_);
  and (_29530_, _29479_, _28623_);
  or (_29531_, _29530_, _12407_);
  or (_29532_, _29531_, _29528_);
  or (_29533_, _12406_, _12139_);
  and (_29534_, _29533_, _12404_);
  and (_29535_, _29534_, _29532_);
  and (_29536_, _29479_, _26288_);
  or (_29537_, _29536_, _06345_);
  or (_29538_, _29537_, _29535_);
  and (_29539_, _29538_, _29498_);
  or (_29541_, _29539_, _12473_);
  or (_29542_, _29479_, _12468_);
  and (_29543_, _29542_, _12477_);
  and (_29544_, _29543_, _29541_);
  or (_29545_, _12477_, _29481_);
  nand (_29546_, _29545_, _12484_);
  or (_29547_, _29546_, _29544_);
  and (_29548_, _29547_, _29497_);
  or (_29549_, _29548_, _06423_);
  and (_29550_, _29549_, _06420_);
  and (_29552_, _29550_, _29492_);
  or (_29553_, _29489_, _12559_);
  or (_29554_, _12560_, _12264_);
  and (_29555_, _29554_, _06419_);
  and (_29556_, _29555_, _29553_);
  or (_29557_, _29556_, _12254_);
  or (_29558_, _25279_, _12264_);
  or (_29559_, _29489_, _12540_);
  and (_29560_, _29559_, _06347_);
  and (_29561_, _29560_, _29558_);
  or (_29563_, _29561_, _29557_);
  or (_29564_, _29563_, _29552_);
  or (_29565_, _29479_, _12255_);
  and (_29566_, _29565_, _12579_);
  and (_29567_, _29566_, _29564_);
  nor (_29568_, _12579_, _29481_);
  or (_29569_, _29568_, _12589_);
  or (_29570_, _29569_, _29567_);
  or (_29571_, _29479_, _12585_);
  and (_29572_, _29571_, _12591_);
  and (_29574_, _29572_, _29570_);
  or (_29575_, _12591_, _29481_);
  nand (_29576_, _29575_, _12595_);
  or (_29577_, _29576_, _29574_);
  or (_29578_, _29479_, _12595_);
  and (_29579_, _29578_, _12599_);
  and (_29580_, _29579_, _29577_);
  nor (_29581_, _29481_, _12599_);
  or (_29582_, _29581_, _05976_);
  or (_29583_, _29582_, _29580_);
  or (_29585_, _29479_, _05940_);
  and (_29586_, _29585_, _12609_);
  and (_29587_, _29586_, _29583_);
  nor (_29588_, _12609_, _29481_);
  or (_29589_, _29588_, _06395_);
  or (_29590_, _29589_, _29587_);
  or (_29591_, _12264_, _06396_);
  and (_29592_, _29591_, _06261_);
  and (_29593_, _29592_, _29590_);
  nor (_29594_, _29481_, _06261_);
  or (_29596_, _29594_, _05972_);
  or (_29597_, _29596_, _29593_);
  or (_29598_, _12264_, _06251_);
  and (_29599_, _29598_, _12252_);
  and (_29600_, _29599_, _29597_);
  and (_29601_, _29479_, _12626_);
  or (_29602_, _29601_, _12625_);
  or (_29603_, _29602_, _29600_);
  or (_29604_, _12624_, _12139_);
  and (_29605_, _29604_, _12631_);
  and (_29607_, _29605_, _29603_);
  and (_29608_, _29505_, _12630_);
  or (_29609_, _29608_, _09016_);
  or (_29610_, _29609_, _29607_);
  or (_29611_, _12139_, _09015_);
  and (_29612_, _29611_, _29610_);
  or (_29613_, _29612_, _06215_);
  or (_29614_, _12264_, _06216_);
  and (_29615_, _29614_, _10892_);
  and (_29616_, _29615_, _29613_);
  and (_29618_, _12139_, _10891_);
  or (_29619_, _29618_, _12644_);
  or (_29620_, _29619_, _29616_);
  nor (_29621_, _12674_, \oc8051_golden_model_1.DPH [6]);
  nor (_29622_, _29621_, _12675_);
  or (_29623_, _29622_, _25380_);
  and (_29624_, _29623_, _12680_);
  and (_29625_, _29624_, _29620_);
  or (_29626_, _29625_, _29486_);
  and (_29627_, _29626_, _12685_);
  or (_29629_, _29505_, _11327_);
  or (_29630_, _12139_, _12248_);
  and (_29631_, _29630_, _12247_);
  and (_29632_, _29631_, _29629_);
  or (_29633_, _29632_, _12697_);
  or (_29634_, _29633_, _29627_);
  or (_29635_, _29479_, _12695_);
  and (_29636_, _29635_, _12699_);
  and (_29637_, _29636_, _29634_);
  nor (_29638_, _12699_, _29481_);
  or (_29640_, _29638_, _06398_);
  or (_29641_, _29640_, _29637_);
  or (_29642_, _12264_, _09025_);
  and (_29643_, _29642_, _12708_);
  and (_29644_, _29643_, _29641_);
  or (_29645_, _29644_, _29484_);
  and (_29646_, _29645_, _12712_);
  or (_29647_, _29505_, _12248_);
  or (_29648_, _12139_, _11327_);
  and (_29649_, _29648_, _12711_);
  and (_29651_, _29649_, _29647_);
  or (_29652_, _29651_, _12720_);
  or (_29653_, _29652_, _29646_);
  or (_29654_, _29479_, _12244_);
  and (_29655_, _29654_, _10969_);
  and (_29656_, _29655_, _29653_);
  nor (_29657_, _29481_, _10969_);
  or (_29658_, _29657_, _06426_);
  or (_29659_, _29658_, _29656_);
  or (_29660_, _12264_, _07219_);
  and (_29662_, _29660_, _12729_);
  and (_29663_, _29662_, _29659_);
  or (_29664_, _29663_, _29483_);
  and (_29665_, _29664_, _12733_);
  or (_29666_, _29505_, \oc8051_golden_model_1.PSW [7]);
  or (_29667_, _12139_, _10774_);
  and (_29668_, _29667_, _12732_);
  and (_29669_, _29668_, _29666_);
  or (_29670_, _29669_, _12751_);
  or (_29671_, _29670_, _29665_);
  or (_29673_, _29479_, _12749_);
  and (_29674_, _29673_, _11007_);
  and (_29675_, _29674_, _29671_);
  nor (_29676_, _29481_, _11007_);
  or (_29677_, _29676_, _06437_);
  or (_29678_, _29677_, _29675_);
  or (_29679_, _12264_, _07229_);
  and (_29680_, _29679_, _12759_);
  and (_29681_, _29680_, _29678_);
  or (_29682_, _29681_, _29482_);
  and (_29684_, _29682_, _12762_);
  or (_29685_, _29505_, _10774_);
  or (_29686_, _12139_, \oc8051_golden_model_1.PSW [7]);
  and (_29687_, _29686_, _12239_);
  and (_29688_, _29687_, _29685_);
  or (_29689_, _29688_, _12771_);
  or (_29690_, _29689_, _29684_);
  or (_29691_, _29479_, _12767_);
  and (_29692_, _29691_, _12769_);
  and (_29693_, _29692_, _29690_);
  nor (_29695_, _29481_, _12769_);
  or (_29696_, _29695_, _11111_);
  or (_29697_, _29696_, _29693_);
  or (_29698_, _29479_, _12775_);
  and (_29699_, _29698_, _12782_);
  and (_29700_, _29699_, _29697_);
  and (_29701_, _09418_, _06543_);
  or (_29702_, _29701_, _06011_);
  or (_29703_, _29702_, _29700_);
  or (_29704_, _12139_, _09057_);
  and (_29705_, _29704_, _12786_);
  and (_29706_, _29705_, _29703_);
  or (_29707_, _12264_, _12970_);
  or (_29708_, _29489_, _25133_);
  and (_29709_, _29708_, _06436_);
  and (_29710_, _29709_, _29707_);
  or (_29711_, _29710_, _12790_);
  or (_29712_, _29711_, _29706_);
  or (_29713_, _29479_, _12129_);
  and (_29714_, _29713_, _12978_);
  and (_29717_, _29714_, _29712_);
  nor (_29718_, _12978_, _29481_);
  or (_29719_, _29718_, _10472_);
  or (_29720_, _29719_, _29717_);
  and (_29721_, _29720_, _29480_);
  or (_29722_, _29721_, _06290_);
  or (_29723_, _09418_, _06291_);
  and (_29724_, _29723_, _25143_);
  and (_29725_, _29724_, _29722_);
  and (_29726_, _12139_, _05994_);
  or (_29728_, _29726_, _06434_);
  or (_29729_, _29728_, _29725_);
  or (_29730_, _12264_, _25133_);
  or (_29731_, _29489_, _12970_);
  and (_29732_, _29731_, _29730_);
  or (_29733_, _29732_, _06435_);
  and (_29734_, _29733_, _29729_);
  or (_29735_, _29734_, _12999_);
  or (_29736_, _29479_, _12998_);
  and (_29737_, _29736_, _29735_);
  or (_29739_, _29737_, _06559_);
  or (_29740_, _12139_, _07240_);
  and (_29741_, _29740_, _13005_);
  and (_29742_, _29741_, _29739_);
  and (_29743_, _29479_, _26914_);
  or (_29744_, _29743_, _06432_);
  or (_29745_, _29744_, _29742_);
  nand (_29746_, _06432_, _06325_);
  and (_29747_, _29746_, _14666_);
  and (_29748_, _29747_, _29745_);
  and (_29750_, _12139_, _05991_);
  or (_29751_, _29750_, _05932_);
  or (_29752_, _29751_, _29748_);
  or (_29753_, _29732_, _05933_);
  and (_29754_, _29753_, _13019_);
  and (_29755_, _29754_, _29752_);
  and (_29756_, _29479_, _13020_);
  or (_29757_, _29756_, _06566_);
  or (_29758_, _29757_, _29755_);
  or (_29759_, _12139_, _06570_);
  and (_29761_, _29759_, _13027_);
  and (_29762_, _29761_, _29758_);
  and (_29763_, _29479_, _26930_);
  or (_29764_, _29763_, _06393_);
  or (_29765_, _29764_, _29762_);
  nand (_29766_, _06393_, _06325_);
  and (_29767_, _29766_, _13036_);
  and (_29768_, _29767_, _29765_);
  and (_29769_, _29479_, _13035_);
  and (_29770_, _12139_, _05989_);
  or (_29772_, _29770_, _01324_);
  or (_29773_, _29772_, _29769_);
  or (_29774_, _29773_, _29768_);
  or (_29775_, _01320_, \oc8051_golden_model_1.PC [14]);
  and (_29776_, _29775_, _42355_);
  and (_42999_, _29776_, _29774_);
  nand (_29777_, _11254_, _07876_);
  and (_29778_, _13046_, \oc8051_golden_model_1.P2 [0]);
  nor (_29779_, _29778_, _07217_);
  nand (_29780_, _29779_, _29777_);
  and (_29782_, _07876_, _07135_);
  or (_29783_, _29782_, _29778_);
  or (_29784_, _29783_, _06260_);
  nor (_29785_, _08374_, _13046_);
  or (_29786_, _29785_, _29778_);
  and (_29787_, _29786_, _06285_);
  and (_29788_, _07144_, \oc8051_golden_model_1.P2 [0]);
  and (_29789_, _07876_, \oc8051_golden_model_1.ACC [0]);
  or (_29790_, _29789_, _29778_);
  and (_29791_, _29790_, _07143_);
  or (_29793_, _29791_, _29788_);
  and (_29794_, _29793_, _06286_);
  or (_29795_, _29794_, _06281_);
  or (_29796_, _29795_, _29787_);
  and (_29797_, _14326_, _08614_);
  and (_29798_, _13051_, \oc8051_golden_model_1.P2 [0]);
  or (_29799_, _29798_, _06282_);
  or (_29800_, _29799_, _29797_);
  and (_29801_, _29800_, _07169_);
  and (_29802_, _29801_, _29796_);
  and (_29804_, _29783_, _06354_);
  or (_29805_, _29804_, _06345_);
  or (_29806_, _29805_, _29802_);
  or (_29807_, _29790_, _06346_);
  and (_29808_, _29807_, _06278_);
  and (_29809_, _29808_, _29806_);
  and (_29810_, _29778_, _06277_);
  or (_29811_, _29810_, _06270_);
  or (_29812_, _29811_, _29809_);
  or (_29813_, _29786_, _06271_);
  and (_29815_, _29813_, _06267_);
  and (_29816_, _29815_, _29812_);
  and (_29817_, _14358_, _08614_);
  or (_29818_, _29817_, _29798_);
  and (_29819_, _29818_, _06266_);
  or (_29820_, _29819_, _06259_);
  or (_29821_, _29820_, _29816_);
  and (_29822_, _29821_, _29784_);
  or (_29823_, _29822_, _09486_);
  and (_29824_, _09384_, _07876_);
  or (_29826_, _29778_, _06258_);
  or (_29827_, _29826_, _29824_);
  and (_29828_, _29827_, _06251_);
  and (_29829_, _29828_, _29823_);
  and (_29830_, _14413_, _07876_);
  or (_29831_, _29830_, _29778_);
  and (_29832_, _29831_, _05972_);
  or (_29833_, _29832_, _29829_);
  or (_29834_, _29833_, _10080_);
  and (_29835_, _14311_, _07876_);
  or (_29837_, _29778_, _09025_);
  or (_29838_, _29837_, _29835_);
  and (_29839_, _07876_, _08929_);
  or (_29840_, _29839_, _29778_);
  or (_29841_, _29840_, _06216_);
  and (_29842_, _29841_, _09030_);
  and (_29843_, _29842_, _29838_);
  and (_29844_, _29843_, _29834_);
  nor (_29845_, _12532_, _13046_);
  or (_29846_, _29845_, _29778_);
  and (_29848_, _29777_, _06524_);
  and (_29849_, _29848_, _29846_);
  or (_29850_, _29849_, _29844_);
  and (_29851_, _29850_, _07219_);
  nand (_29852_, _29840_, _06426_);
  nor (_29853_, _29852_, _29785_);
  or (_29854_, _29853_, _06532_);
  or (_29855_, _29854_, _29851_);
  and (_29856_, _29855_, _29780_);
  or (_29857_, _29856_, _06437_);
  and (_29859_, _14307_, _07876_);
  or (_29860_, _29778_, _07229_);
  or (_29861_, _29860_, _29859_);
  and (_29862_, _29861_, _07231_);
  and (_29863_, _29862_, _29857_);
  and (_29864_, _29846_, _06535_);
  or (_29865_, _29864_, _06559_);
  or (_29866_, _29865_, _29863_);
  or (_29867_, _29786_, _07240_);
  and (_29868_, _29867_, _29866_);
  or (_29870_, _29868_, _05932_);
  or (_29871_, _29778_, _05933_);
  and (_29872_, _29871_, _29870_);
  or (_29873_, _29872_, _06566_);
  or (_29874_, _29786_, _06570_);
  and (_29875_, _29874_, _01320_);
  and (_29876_, _29875_, _29873_);
  nor (_29877_, \oc8051_golden_model_1.P2 [0], rst);
  nor (_29878_, _29877_, _00000_);
  or (_43000_, _29878_, _29876_);
  nor (_29880_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_29881_, _29880_, _00000_);
  and (_29882_, _13046_, \oc8051_golden_model_1.P2 [1]);
  nor (_29883_, _11252_, _13046_);
  or (_29884_, _29883_, _29882_);
  or (_29885_, _29884_, _07231_);
  and (_29886_, _07876_, _09422_);
  or (_29887_, _29886_, _29882_);
  or (_29888_, _29887_, _07169_);
  or (_29889_, _07876_, \oc8051_golden_model_1.P2 [1]);
  and (_29891_, _14520_, _07876_);
  not (_29892_, _29891_);
  and (_29893_, _29892_, _29889_);
  or (_29894_, _29893_, _06286_);
  and (_29895_, _07876_, \oc8051_golden_model_1.ACC [1]);
  or (_29896_, _29895_, _29882_);
  and (_29897_, _29896_, _07143_);
  and (_29898_, _07144_, \oc8051_golden_model_1.P2 [1]);
  or (_29899_, _29898_, _06285_);
  or (_29900_, _29899_, _29897_);
  and (_29902_, _29900_, _06282_);
  and (_29903_, _29902_, _29894_);
  and (_29904_, _13051_, \oc8051_golden_model_1.P2 [1]);
  and (_29905_, _14508_, _08614_);
  or (_29906_, _29905_, _29904_);
  and (_29907_, _29906_, _06281_);
  or (_29908_, _29907_, _06354_);
  or (_29909_, _29908_, _29903_);
  and (_29910_, _29909_, _29888_);
  or (_29911_, _29910_, _06345_);
  or (_29913_, _29896_, _06346_);
  and (_29914_, _29913_, _06278_);
  and (_29915_, _29914_, _29911_);
  and (_29916_, _14511_, _08614_);
  or (_29917_, _29916_, _29904_);
  and (_29918_, _29917_, _06277_);
  or (_29919_, _29918_, _06270_);
  or (_29920_, _29919_, _29915_);
  and (_29921_, _29905_, _14507_);
  or (_29922_, _29904_, _06271_);
  or (_29924_, _29922_, _29921_);
  and (_29925_, _29924_, _06267_);
  and (_29926_, _29925_, _29920_);
  or (_29927_, _29904_, _14551_);
  and (_29928_, _29927_, _06266_);
  and (_29929_, _29928_, _29906_);
  or (_29930_, _29929_, _06259_);
  or (_29931_, _29930_, _29926_);
  or (_29932_, _29887_, _06260_);
  and (_29933_, _29932_, _29931_);
  or (_29935_, _29933_, _09486_);
  and (_29936_, _09339_, _07876_);
  or (_29937_, _29882_, _06258_);
  or (_29938_, _29937_, _29936_);
  and (_29939_, _29938_, _06251_);
  and (_29940_, _29939_, _29935_);
  and (_29941_, _14607_, _07876_);
  or (_29942_, _29941_, _29882_);
  and (_29943_, _29942_, _05972_);
  or (_29944_, _29943_, _29940_);
  and (_29946_, _29944_, _06399_);
  or (_29947_, _14505_, _13046_);
  and (_29948_, _29947_, _06398_);
  nand (_29949_, _07876_, _07031_);
  and (_29950_, _29949_, _06215_);
  or (_29951_, _29950_, _29948_);
  and (_29952_, _29951_, _29889_);
  or (_29953_, _29952_, _06524_);
  or (_29954_, _29953_, _29946_);
  nand (_29955_, _11251_, _07876_);
  and (_29957_, _29955_, _29884_);
  or (_29958_, _29957_, _09030_);
  and (_29959_, _29958_, _07219_);
  and (_29960_, _29959_, _29954_);
  or (_29961_, _14503_, _13046_);
  and (_29962_, _29889_, _06426_);
  and (_29963_, _29962_, _29961_);
  or (_29964_, _29963_, _06532_);
  or (_29965_, _29964_, _29960_);
  nor (_29966_, _29882_, _07217_);
  nand (_29968_, _29966_, _29955_);
  and (_29969_, _29968_, _07229_);
  and (_29970_, _29969_, _29965_);
  or (_29971_, _29949_, _08325_);
  and (_29972_, _29889_, _06437_);
  and (_29973_, _29972_, _29971_);
  or (_29974_, _29973_, _06535_);
  or (_29975_, _29974_, _29970_);
  and (_29976_, _29975_, _29885_);
  or (_29977_, _29976_, _06559_);
  or (_29979_, _29893_, _07240_);
  and (_29980_, _29979_, _05933_);
  and (_29981_, _29980_, _29977_);
  and (_29982_, _29917_, _05932_);
  or (_29983_, _29982_, _06566_);
  or (_29984_, _29983_, _29981_);
  or (_29985_, _29882_, _06570_);
  or (_29986_, _29985_, _29891_);
  and (_29987_, _29986_, _01320_);
  and (_29988_, _29987_, _29984_);
  or (_43002_, _29988_, _29881_);
  and (_29990_, _13046_, \oc8051_golden_model_1.P2 [2]);
  and (_29991_, _07876_, _08662_);
  or (_29992_, _29991_, _29990_);
  or (_29993_, _29992_, _06260_);
  or (_29994_, _29992_, _07169_);
  and (_29995_, _14703_, _07876_);
  or (_29996_, _29995_, _29990_);
  or (_29997_, _29996_, _06286_);
  and (_29998_, _07876_, \oc8051_golden_model_1.ACC [2]);
  or (_30000_, _29998_, _29990_);
  and (_30001_, _30000_, _07143_);
  and (_30002_, _07144_, \oc8051_golden_model_1.P2 [2]);
  or (_30003_, _30002_, _06285_);
  or (_30004_, _30003_, _30001_);
  and (_30005_, _30004_, _06282_);
  and (_30006_, _30005_, _29997_);
  and (_30007_, _13051_, \oc8051_golden_model_1.P2 [2]);
  and (_30008_, _14716_, _08614_);
  or (_30009_, _30008_, _30007_);
  and (_30011_, _30009_, _06281_);
  or (_30012_, _30011_, _06354_);
  or (_30013_, _30012_, _30006_);
  and (_30014_, _30013_, _29994_);
  or (_30015_, _30014_, _06345_);
  or (_30016_, _30000_, _06346_);
  and (_30017_, _30016_, _06278_);
  and (_30018_, _30017_, _30015_);
  and (_30019_, _14699_, _08614_);
  or (_30020_, _30019_, _30007_);
  and (_30022_, _30020_, _06277_);
  or (_30023_, _30022_, _06270_);
  or (_30024_, _30023_, _30018_);
  and (_30025_, _30008_, _14731_);
  or (_30026_, _30007_, _06271_);
  or (_30027_, _30026_, _30025_);
  and (_30028_, _30027_, _06267_);
  and (_30029_, _30028_, _30024_);
  and (_30030_, _14749_, _08614_);
  or (_30031_, _30030_, _30007_);
  and (_30033_, _30031_, _06266_);
  or (_30034_, _30033_, _06259_);
  or (_30035_, _30034_, _30029_);
  and (_30036_, _30035_, _29993_);
  or (_30037_, _30036_, _09486_);
  and (_30038_, _09293_, _07876_);
  or (_30039_, _29990_, _06258_);
  or (_30040_, _30039_, _30038_);
  and (_30041_, _30040_, _06251_);
  and (_30042_, _30041_, _30037_);
  and (_30044_, _14804_, _07876_);
  or (_30045_, _29990_, _30044_);
  and (_30046_, _30045_, _05972_);
  or (_30047_, _30046_, _30042_);
  or (_30048_, _30047_, _10080_);
  and (_30049_, _14697_, _07876_);
  or (_30050_, _29990_, _09025_);
  or (_30051_, _30050_, _30049_);
  and (_30052_, _07876_, _08980_);
  or (_30053_, _30052_, _29990_);
  or (_30055_, _30053_, _06216_);
  and (_30056_, _30055_, _09030_);
  and (_30057_, _30056_, _30051_);
  and (_30058_, _30057_, _30048_);
  and (_30059_, _11250_, _07876_);
  or (_30060_, _30059_, _29990_);
  and (_30061_, _30060_, _06524_);
  or (_30062_, _30061_, _30058_);
  and (_30063_, _30062_, _07219_);
  or (_30064_, _29990_, _08424_);
  and (_30066_, _30053_, _06426_);
  and (_30067_, _30066_, _30064_);
  or (_30068_, _30067_, _30063_);
  and (_30069_, _30068_, _07217_);
  and (_30070_, _30000_, _06532_);
  and (_30071_, _30070_, _30064_);
  or (_30072_, _30071_, _06437_);
  or (_30073_, _30072_, _30069_);
  and (_30074_, _14694_, _07876_);
  or (_30075_, _29990_, _07229_);
  or (_30077_, _30075_, _30074_);
  and (_30078_, _30077_, _07231_);
  and (_30079_, _30078_, _30073_);
  nor (_30080_, _11249_, _13046_);
  or (_30081_, _30080_, _29990_);
  and (_30082_, _30081_, _06535_);
  or (_30083_, _30082_, _06559_);
  or (_30084_, _30083_, _30079_);
  or (_30085_, _29996_, _07240_);
  and (_30086_, _30085_, _05933_);
  and (_30088_, _30086_, _30084_);
  and (_30089_, _30020_, _05932_);
  or (_30090_, _30089_, _06566_);
  or (_30091_, _30090_, _30088_);
  and (_30092_, _14873_, _07876_);
  or (_30093_, _29990_, _06570_);
  or (_30094_, _30093_, _30092_);
  and (_30095_, _30094_, _01320_);
  and (_30096_, _30095_, _30091_);
  nor (_30097_, \oc8051_golden_model_1.P2 [2], rst);
  nor (_30099_, _30097_, _00000_);
  or (_43003_, _30099_, _30096_);
  and (_30100_, _13046_, \oc8051_golden_model_1.P2 [3]);
  and (_30101_, _07876_, _09421_);
  or (_30102_, _30101_, _30100_);
  or (_30103_, _30102_, _06260_);
  and (_30104_, _14900_, _07876_);
  or (_30105_, _30104_, _30100_);
  or (_30106_, _30105_, _06286_);
  and (_30107_, _07876_, \oc8051_golden_model_1.ACC [3]);
  or (_30109_, _30107_, _30100_);
  and (_30110_, _30109_, _07143_);
  and (_30111_, _07144_, \oc8051_golden_model_1.P2 [3]);
  or (_30112_, _30111_, _06285_);
  or (_30113_, _30112_, _30110_);
  and (_30114_, _30113_, _06282_);
  and (_30115_, _30114_, _30106_);
  and (_30116_, _13051_, \oc8051_golden_model_1.P2 [3]);
  and (_30117_, _14897_, _08614_);
  or (_30118_, _30117_, _30116_);
  and (_30120_, _30118_, _06281_);
  or (_30121_, _30120_, _06354_);
  or (_30122_, _30121_, _30115_);
  or (_30123_, _30102_, _07169_);
  and (_30124_, _30123_, _30122_);
  or (_30125_, _30124_, _06345_);
  or (_30126_, _30109_, _06346_);
  and (_30127_, _30126_, _06278_);
  and (_30128_, _30127_, _30125_);
  and (_30129_, _14895_, _08614_);
  or (_30131_, _30129_, _30116_);
  and (_30132_, _30131_, _06277_);
  or (_30133_, _30132_, _06270_);
  or (_30134_, _30133_, _30128_);
  or (_30135_, _30116_, _14926_);
  and (_30136_, _30135_, _30118_);
  or (_30137_, _30136_, _06271_);
  and (_30138_, _30137_, _06267_);
  and (_30139_, _30138_, _30134_);
  and (_30140_, _14943_, _08614_);
  or (_30142_, _30140_, _30116_);
  and (_30143_, _30142_, _06266_);
  or (_30144_, _30143_, _06259_);
  or (_30145_, _30144_, _30139_);
  and (_30146_, _30145_, _30103_);
  or (_30147_, _30146_, _09486_);
  and (_30148_, _09247_, _07876_);
  or (_30149_, _30100_, _06258_);
  or (_30150_, _30149_, _30148_);
  and (_30151_, _30150_, _06251_);
  and (_30153_, _30151_, _30147_);
  and (_30154_, _14998_, _07876_);
  or (_30155_, _30100_, _30154_);
  and (_30156_, _30155_, _05972_);
  or (_30157_, _30156_, _30153_);
  or (_30158_, _30157_, _10080_);
  and (_30159_, _14893_, _07876_);
  or (_30160_, _30100_, _09025_);
  or (_30161_, _30160_, _30159_);
  and (_30162_, _07876_, _08809_);
  or (_30164_, _30162_, _30100_);
  or (_30165_, _30164_, _06216_);
  and (_30166_, _30165_, _09030_);
  and (_30167_, _30166_, _30161_);
  and (_30168_, _30167_, _30158_);
  and (_30169_, _12529_, _07876_);
  or (_30170_, _30169_, _30100_);
  and (_30171_, _30170_, _06524_);
  or (_30172_, _30171_, _30168_);
  and (_30173_, _30172_, _07219_);
  or (_30175_, _30100_, _08280_);
  and (_30176_, _30164_, _06426_);
  and (_30177_, _30176_, _30175_);
  or (_30178_, _30177_, _30173_);
  and (_30179_, _30178_, _07217_);
  and (_30180_, _30109_, _06532_);
  and (_30181_, _30180_, _30175_);
  or (_30182_, _30181_, _06437_);
  or (_30183_, _30182_, _30179_);
  and (_30184_, _14890_, _07876_);
  or (_30186_, _30100_, _07229_);
  or (_30187_, _30186_, _30184_);
  and (_30188_, _30187_, _07231_);
  and (_30189_, _30188_, _30183_);
  nor (_30190_, _11247_, _13046_);
  or (_30191_, _30190_, _30100_);
  and (_30192_, _30191_, _06535_);
  or (_30193_, _30192_, _06559_);
  or (_30194_, _30193_, _30189_);
  or (_30195_, _30105_, _07240_);
  and (_30197_, _30195_, _05933_);
  and (_30198_, _30197_, _30194_);
  and (_30199_, _30131_, _05932_);
  or (_30200_, _30199_, _06566_);
  or (_30201_, _30200_, _30198_);
  and (_30202_, _15068_, _07876_);
  or (_30203_, _30100_, _06570_);
  or (_30204_, _30203_, _30202_);
  and (_30205_, _30204_, _01320_);
  and (_30206_, _30205_, _30201_);
  nor (_30208_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_30209_, _30208_, _00000_);
  or (_43004_, _30209_, _30206_);
  nor (_30210_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_30211_, _30210_, _00000_);
  and (_30212_, _13046_, \oc8051_golden_model_1.P2 [4]);
  and (_30213_, _09420_, _07876_);
  or (_30214_, _30213_, _30212_);
  or (_30215_, _30214_, _06260_);
  and (_30216_, _13051_, \oc8051_golden_model_1.P2 [4]);
  and (_30218_, _15145_, _08614_);
  or (_30219_, _30218_, _30216_);
  and (_30220_, _30219_, _06277_);
  and (_30221_, _15133_, _07876_);
  or (_30222_, _30221_, _30212_);
  or (_30223_, _30222_, _06286_);
  and (_30224_, _07876_, \oc8051_golden_model_1.ACC [4]);
  or (_30225_, _30224_, _30212_);
  and (_30226_, _30225_, _07143_);
  and (_30227_, _07144_, \oc8051_golden_model_1.P2 [4]);
  or (_30229_, _30227_, _06285_);
  or (_30230_, _30229_, _30226_);
  and (_30231_, _30230_, _06282_);
  and (_30232_, _30231_, _30223_);
  and (_30233_, _15116_, _08614_);
  or (_30234_, _30233_, _30216_);
  and (_30235_, _30234_, _06281_);
  or (_30236_, _30235_, _06354_);
  or (_30237_, _30236_, _30232_);
  or (_30238_, _30214_, _07169_);
  and (_30240_, _30238_, _30237_);
  or (_30241_, _30240_, _06345_);
  or (_30242_, _30225_, _06346_);
  and (_30243_, _30242_, _06278_);
  and (_30244_, _30243_, _30241_);
  or (_30245_, _30244_, _30220_);
  and (_30246_, _30245_, _06271_);
  or (_30247_, _30216_, _15152_);
  and (_30248_, _30247_, _06270_);
  and (_30249_, _30248_, _30234_);
  or (_30251_, _30249_, _30246_);
  and (_30252_, _30251_, _06267_);
  and (_30253_, _15170_, _08614_);
  or (_30254_, _30253_, _30216_);
  and (_30255_, _30254_, _06266_);
  or (_30256_, _30255_, _06259_);
  or (_30257_, _30256_, _30252_);
  and (_30258_, _30257_, _30215_);
  or (_30259_, _30258_, _09486_);
  and (_30260_, _09437_, _07876_);
  or (_30262_, _30212_, _06258_);
  or (_30263_, _30262_, _30260_);
  and (_30264_, _30263_, _06251_);
  and (_30265_, _30264_, _30259_);
  and (_30266_, _15226_, _07876_);
  or (_30267_, _30266_, _30212_);
  and (_30268_, _30267_, _05972_);
  or (_30269_, _30268_, _10080_);
  or (_30270_, _30269_, _30265_);
  and (_30271_, _15114_, _07876_);
  or (_30273_, _30212_, _09025_);
  or (_30274_, _30273_, _30271_);
  and (_30275_, _08919_, _07876_);
  or (_30276_, _30275_, _30212_);
  or (_30277_, _30276_, _06216_);
  and (_30278_, _30277_, _09030_);
  and (_30279_, _30278_, _30274_);
  and (_30280_, _30279_, _30270_);
  and (_30281_, _11245_, _07876_);
  or (_30282_, _30281_, _30212_);
  and (_30284_, _30282_, _06524_);
  or (_30285_, _30284_, _30280_);
  and (_30286_, _30285_, _07219_);
  or (_30287_, _30212_, _08528_);
  and (_30288_, _30276_, _06426_);
  and (_30289_, _30288_, _30287_);
  or (_30290_, _30289_, _30286_);
  and (_30291_, _30290_, _07217_);
  and (_30292_, _30225_, _06532_);
  and (_30293_, _30292_, _30287_);
  or (_30295_, _30293_, _06437_);
  or (_30296_, _30295_, _30291_);
  and (_30297_, _15111_, _07876_);
  or (_30298_, _30212_, _07229_);
  or (_30299_, _30298_, _30297_);
  and (_30300_, _30299_, _07231_);
  and (_30301_, _30300_, _30296_);
  nor (_30302_, _11244_, _13046_);
  or (_30303_, _30302_, _30212_);
  and (_30304_, _30303_, _06535_);
  or (_30306_, _30304_, _06559_);
  or (_30307_, _30306_, _30301_);
  or (_30308_, _30222_, _07240_);
  and (_30309_, _30308_, _05933_);
  and (_30310_, _30309_, _30307_);
  and (_30311_, _30219_, _05932_);
  or (_30312_, _30311_, _06566_);
  or (_30313_, _30312_, _30310_);
  and (_30314_, _15296_, _07876_);
  or (_30315_, _30212_, _06570_);
  or (_30317_, _30315_, _30314_);
  and (_30318_, _30317_, _01320_);
  and (_30319_, _30318_, _30313_);
  or (_43005_, _30319_, _30211_);
  and (_30320_, _13046_, \oc8051_golden_model_1.P2 [5]);
  and (_30321_, _15330_, _07876_);
  or (_30322_, _30321_, _30320_);
  or (_30323_, _30322_, _06286_);
  and (_30324_, _07876_, \oc8051_golden_model_1.ACC [5]);
  or (_30325_, _30324_, _30320_);
  and (_30326_, _30325_, _07143_);
  and (_30327_, _07144_, \oc8051_golden_model_1.P2 [5]);
  or (_30328_, _30327_, _06285_);
  or (_30329_, _30328_, _30326_);
  and (_30330_, _30329_, _06282_);
  and (_30331_, _30330_, _30323_);
  and (_30332_, _13051_, \oc8051_golden_model_1.P2 [5]);
  and (_30333_, _15315_, _08614_);
  or (_30334_, _30333_, _30332_);
  and (_30335_, _30334_, _06281_);
  or (_30338_, _30335_, _06354_);
  or (_30339_, _30338_, _30331_);
  and (_30340_, _09419_, _07876_);
  or (_30341_, _30340_, _30320_);
  or (_30342_, _30341_, _07169_);
  and (_30343_, _30342_, _30339_);
  or (_30344_, _30343_, _06345_);
  or (_30345_, _30325_, _06346_);
  and (_30346_, _30345_, _06278_);
  and (_30347_, _30346_, _30344_);
  and (_30349_, _15342_, _08614_);
  or (_30350_, _30349_, _30332_);
  and (_30351_, _30350_, _06277_);
  or (_30352_, _30351_, _06270_);
  or (_30353_, _30352_, _30347_);
  or (_30354_, _30332_, _15349_);
  and (_30355_, _30354_, _30334_);
  or (_30356_, _30355_, _06271_);
  and (_30357_, _30356_, _06267_);
  and (_30358_, _30357_, _30353_);
  or (_30360_, _30332_, _15365_);
  and (_30361_, _30360_, _06266_);
  and (_30362_, _30361_, _30334_);
  or (_30363_, _30362_, _06259_);
  or (_30364_, _30363_, _30358_);
  or (_30365_, _30341_, _06260_);
  and (_30366_, _30365_, _30364_);
  or (_30367_, _30366_, _09486_);
  and (_30368_, _09436_, _07876_);
  or (_30369_, _30320_, _06258_);
  or (_30371_, _30369_, _30368_);
  and (_30372_, _30371_, _06251_);
  and (_30373_, _30372_, _30367_);
  and (_30374_, _15421_, _07876_);
  or (_30375_, _30374_, _30320_);
  and (_30376_, _30375_, _05972_);
  or (_30377_, _30376_, _10080_);
  or (_30378_, _30377_, _30373_);
  and (_30379_, _15313_, _07876_);
  or (_30380_, _30320_, _09025_);
  or (_30382_, _30380_, _30379_);
  and (_30383_, _08913_, _07876_);
  or (_30384_, _30383_, _30320_);
  or (_30385_, _30384_, _06216_);
  and (_30386_, _30385_, _09030_);
  and (_30387_, _30386_, _30382_);
  and (_30388_, _30387_, _30378_);
  and (_30389_, _12536_, _07876_);
  or (_30390_, _30389_, _30320_);
  and (_30391_, _30390_, _06524_);
  or (_30393_, _30391_, _30388_);
  and (_30394_, _30393_, _07219_);
  or (_30395_, _30320_, _08231_);
  and (_30396_, _30384_, _06426_);
  and (_30397_, _30396_, _30395_);
  or (_30398_, _30397_, _30394_);
  and (_30399_, _30398_, _07217_);
  and (_30400_, _30325_, _06532_);
  and (_30401_, _30400_, _30395_);
  or (_30402_, _30401_, _06437_);
  or (_30404_, _30402_, _30399_);
  and (_30405_, _15310_, _07876_);
  or (_30406_, _30320_, _07229_);
  or (_30407_, _30406_, _30405_);
  and (_30408_, _30407_, _07231_);
  and (_30409_, _30408_, _30404_);
  nor (_30410_, _11241_, _13046_);
  or (_30411_, _30410_, _30320_);
  and (_30412_, _30411_, _06535_);
  or (_30413_, _30412_, _06559_);
  or (_30415_, _30413_, _30409_);
  or (_30416_, _30322_, _07240_);
  and (_30417_, _30416_, _05933_);
  and (_30418_, _30417_, _30415_);
  and (_30419_, _30350_, _05932_);
  or (_30420_, _30419_, _06566_);
  or (_30421_, _30420_, _30418_);
  and (_30422_, _15493_, _07876_);
  or (_30423_, _30320_, _06570_);
  or (_30424_, _30423_, _30422_);
  and (_30426_, _30424_, _01320_);
  and (_30427_, _30426_, _30421_);
  nor (_30428_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_30429_, _30428_, _00000_);
  or (_43006_, _30429_, _30427_);
  and (_30430_, _13046_, \oc8051_golden_model_1.P2 [6]);
  and (_30431_, _15521_, _07876_);
  or (_30432_, _30431_, _30430_);
  or (_30433_, _30432_, _06286_);
  and (_30434_, _07876_, \oc8051_golden_model_1.ACC [6]);
  or (_30436_, _30434_, _30430_);
  and (_30437_, _30436_, _07143_);
  and (_30438_, _07144_, \oc8051_golden_model_1.P2 [6]);
  or (_30439_, _30438_, _06285_);
  or (_30440_, _30439_, _30437_);
  and (_30441_, _30440_, _06282_);
  and (_30442_, _30441_, _30433_);
  and (_30443_, _13051_, \oc8051_golden_model_1.P2 [6]);
  and (_30444_, _15535_, _08614_);
  or (_30445_, _30444_, _30443_);
  and (_30447_, _30445_, _06281_);
  or (_30448_, _30447_, _06354_);
  or (_30449_, _30448_, _30442_);
  and (_30450_, _09418_, _07876_);
  or (_30451_, _30450_, _30430_);
  or (_30452_, _30451_, _07169_);
  and (_30453_, _30452_, _30449_);
  or (_30454_, _30453_, _06345_);
  or (_30455_, _30436_, _06346_);
  and (_30456_, _30455_, _06278_);
  and (_30458_, _30456_, _30454_);
  and (_30459_, _15544_, _08614_);
  or (_30460_, _30459_, _30443_);
  and (_30461_, _30460_, _06277_);
  or (_30462_, _30461_, _06270_);
  or (_30463_, _30462_, _30458_);
  or (_30464_, _30443_, _15551_);
  and (_30465_, _30464_, _30445_);
  or (_30466_, _30465_, _06271_);
  and (_30467_, _30466_, _06267_);
  and (_30469_, _30467_, _30463_);
  and (_30470_, _15568_, _08614_);
  or (_30471_, _30470_, _30443_);
  and (_30472_, _30471_, _06266_);
  or (_30473_, _30472_, _06259_);
  or (_30474_, _30473_, _30469_);
  or (_30475_, _30451_, _06260_);
  and (_30476_, _30475_, _30474_);
  or (_30477_, _30476_, _09486_);
  and (_30478_, _09435_, _07876_);
  or (_30480_, _30430_, _06258_);
  or (_30481_, _30480_, _30478_);
  and (_30482_, _30481_, _06251_);
  and (_30483_, _30482_, _30477_);
  and (_30484_, _15623_, _07876_);
  or (_30485_, _30484_, _30430_);
  and (_30486_, _30485_, _05972_);
  or (_30487_, _30486_, _10080_);
  or (_30488_, _30487_, _30483_);
  and (_30489_, _15517_, _07876_);
  or (_30491_, _30430_, _09025_);
  or (_30492_, _30491_, _30489_);
  and (_30493_, _08845_, _07876_);
  or (_30494_, _30493_, _30430_);
  or (_30495_, _30494_, _06216_);
  and (_30496_, _30495_, _09030_);
  and (_30497_, _30496_, _30492_);
  and (_30498_, _30497_, _30488_);
  and (_30499_, _11239_, _07876_);
  or (_30500_, _30499_, _30430_);
  and (_30502_, _30500_, _06524_);
  or (_30503_, _30502_, _30498_);
  and (_30504_, _30503_, _07219_);
  or (_30505_, _30430_, _08128_);
  and (_30506_, _30494_, _06426_);
  and (_30507_, _30506_, _30505_);
  or (_30508_, _30507_, _30504_);
  and (_30509_, _30508_, _07217_);
  and (_30510_, _30436_, _06532_);
  and (_30511_, _30510_, _30505_);
  or (_30513_, _30511_, _06437_);
  or (_30514_, _30513_, _30509_);
  and (_30515_, _15514_, _07876_);
  or (_30516_, _30430_, _07229_);
  or (_30517_, _30516_, _30515_);
  and (_30518_, _30517_, _07231_);
  and (_30519_, _30518_, _30514_);
  nor (_30520_, _11238_, _13046_);
  or (_30521_, _30520_, _30430_);
  and (_30522_, _30521_, _06535_);
  or (_30524_, _30522_, _06559_);
  or (_30525_, _30524_, _30519_);
  or (_30526_, _30432_, _07240_);
  and (_30527_, _30526_, _05933_);
  and (_30528_, _30527_, _30525_);
  and (_30529_, _30460_, _05932_);
  or (_30530_, _30529_, _06566_);
  or (_30531_, _30530_, _30528_);
  and (_30532_, _15695_, _07876_);
  or (_30533_, _30430_, _06570_);
  or (_30535_, _30533_, _30532_);
  and (_30536_, _30535_, _01320_);
  and (_30537_, _30536_, _30531_);
  nor (_30538_, \oc8051_golden_model_1.P2 [6], rst);
  nor (_30539_, _30538_, _00000_);
  or (_43007_, _30539_, _30537_);
  and (_30540_, _07885_, \oc8051_golden_model_1.ACC [0]);
  and (_30541_, _30540_, _08374_);
  and (_30542_, _13148_, \oc8051_golden_model_1.P3 [0]);
  or (_30543_, _30542_, _07217_);
  or (_30545_, _30543_, _30541_);
  and (_30546_, _07885_, _07135_);
  or (_30547_, _30546_, _30542_);
  or (_30548_, _30547_, _06260_);
  nor (_30549_, _08374_, _13148_);
  or (_30550_, _30549_, _30542_);
  or (_30551_, _30550_, _06286_);
  or (_30552_, _30540_, _30542_);
  and (_30553_, _30552_, _07143_);
  and (_30554_, _07144_, \oc8051_golden_model_1.P3 [0]);
  or (_30556_, _30554_, _06285_);
  or (_30557_, _30556_, _30553_);
  and (_30558_, _30557_, _06282_);
  and (_30559_, _30558_, _30551_);
  and (_30560_, _13153_, \oc8051_golden_model_1.P3 [0]);
  and (_30561_, _14326_, _08607_);
  or (_30562_, _30561_, _30560_);
  and (_30563_, _30562_, _06281_);
  or (_30564_, _30563_, _30559_);
  and (_30565_, _30564_, _07169_);
  and (_30567_, _30547_, _06354_);
  or (_30568_, _30567_, _06345_);
  or (_30569_, _30568_, _30565_);
  or (_30570_, _30552_, _06346_);
  and (_30571_, _30570_, _06278_);
  and (_30572_, _30571_, _30569_);
  and (_30573_, _30542_, _06277_);
  or (_30574_, _30573_, _06270_);
  or (_30575_, _30574_, _30572_);
  or (_30576_, _30550_, _06271_);
  and (_30578_, _30576_, _06267_);
  and (_30579_, _30578_, _30575_);
  and (_30580_, _14358_, _08607_);
  or (_30581_, _30580_, _30560_);
  and (_30582_, _30581_, _06266_);
  or (_30583_, _30582_, _06259_);
  or (_30584_, _30583_, _30579_);
  and (_30585_, _30584_, _30548_);
  or (_30586_, _30585_, _09486_);
  and (_30587_, _09384_, _07885_);
  or (_30589_, _30542_, _06258_);
  or (_30590_, _30589_, _30587_);
  and (_30591_, _30590_, _06251_);
  and (_30592_, _30591_, _30586_);
  and (_30593_, _14413_, _07885_);
  or (_30594_, _30593_, _30542_);
  and (_30595_, _30594_, _05972_);
  or (_30596_, _30595_, _30592_);
  or (_30597_, _30596_, _10080_);
  and (_30598_, _14311_, _07885_);
  or (_30600_, _30542_, _09025_);
  or (_30601_, _30600_, _30598_);
  and (_30602_, _07885_, _08929_);
  or (_30603_, _30602_, _30542_);
  or (_30604_, _30603_, _06216_);
  and (_30605_, _30604_, _09030_);
  and (_30606_, _30605_, _30601_);
  and (_30607_, _30606_, _30597_);
  nor (_30608_, _12532_, _13148_);
  or (_30609_, _30608_, _30542_);
  nor (_30611_, _30541_, _09030_);
  and (_30612_, _30611_, _30609_);
  or (_30613_, _30612_, _30607_);
  and (_30614_, _30613_, _07219_);
  nand (_30615_, _30603_, _06426_);
  nor (_30616_, _30615_, _30549_);
  or (_30617_, _30616_, _06532_);
  or (_30618_, _30617_, _30614_);
  and (_30619_, _30618_, _30545_);
  or (_30620_, _30619_, _06437_);
  and (_30622_, _14307_, _07885_);
  or (_30623_, _30622_, _30542_);
  or (_30624_, _30623_, _07229_);
  and (_30625_, _30624_, _07231_);
  and (_30626_, _30625_, _30620_);
  and (_30627_, _30609_, _06535_);
  or (_30628_, _30627_, _06559_);
  or (_30629_, _30628_, _30626_);
  or (_30630_, _30550_, _07240_);
  and (_30631_, _30630_, _30629_);
  or (_30633_, _30631_, _05932_);
  or (_30634_, _30542_, _05933_);
  and (_30635_, _30634_, _30633_);
  or (_30636_, _30635_, _06566_);
  or (_30637_, _30550_, _06570_);
  and (_30638_, _30637_, _01320_);
  and (_30639_, _30638_, _30636_);
  nor (_30640_, \oc8051_golden_model_1.P3 [0], rst);
  nor (_30641_, _30640_, _00000_);
  or (_43009_, _30641_, _30639_);
  and (_30643_, _13148_, \oc8051_golden_model_1.P3 [1]);
  nor (_30644_, _11252_, _13148_);
  or (_30645_, _30644_, _30643_);
  or (_30646_, _30645_, _07231_);
  and (_30647_, _07885_, _09422_);
  or (_30648_, _30647_, _30643_);
  or (_30649_, _30648_, _07169_);
  or (_30650_, _07885_, \oc8051_golden_model_1.P3 [1]);
  and (_30651_, _14520_, _07885_);
  not (_30652_, _30651_);
  and (_30654_, _30652_, _30650_);
  or (_30655_, _30654_, _06286_);
  and (_30656_, _07885_, \oc8051_golden_model_1.ACC [1]);
  or (_30657_, _30656_, _30643_);
  and (_30658_, _30657_, _07143_);
  and (_30659_, _07144_, \oc8051_golden_model_1.P3 [1]);
  or (_30660_, _30659_, _06285_);
  or (_30661_, _30660_, _30658_);
  and (_30662_, _30661_, _06282_);
  and (_30663_, _30662_, _30655_);
  and (_30665_, _13153_, \oc8051_golden_model_1.P3 [1]);
  and (_30666_, _14508_, _08607_);
  or (_30667_, _30666_, _30665_);
  and (_30668_, _30667_, _06281_);
  or (_30669_, _30668_, _06354_);
  or (_30670_, _30669_, _30663_);
  and (_30671_, _30670_, _30649_);
  or (_30672_, _30671_, _06345_);
  or (_30673_, _30657_, _06346_);
  and (_30674_, _30673_, _06278_);
  and (_30676_, _30674_, _30672_);
  and (_30677_, _14511_, _08607_);
  or (_30678_, _30677_, _30665_);
  and (_30679_, _30678_, _06277_);
  or (_30680_, _30679_, _06270_);
  or (_30681_, _30680_, _30676_);
  and (_30682_, _30666_, _14507_);
  or (_30683_, _30665_, _06271_);
  or (_30684_, _30683_, _30682_);
  and (_30685_, _30684_, _06267_);
  and (_30687_, _30685_, _30681_);
  or (_30688_, _30665_, _14551_);
  and (_30689_, _30688_, _06266_);
  and (_30690_, _30689_, _30667_);
  or (_30691_, _30690_, _06259_);
  or (_30692_, _30691_, _30687_);
  or (_30693_, _30648_, _06260_);
  and (_30694_, _30693_, _30692_);
  or (_30695_, _30694_, _09486_);
  and (_30696_, _09339_, _07885_);
  or (_30698_, _30643_, _06258_);
  or (_30699_, _30698_, _30696_);
  and (_30700_, _30699_, _06251_);
  and (_30701_, _30700_, _30695_);
  and (_30702_, _14607_, _07885_);
  or (_30703_, _30702_, _30643_);
  and (_30704_, _30703_, _05972_);
  or (_30705_, _30704_, _30701_);
  and (_30706_, _30705_, _06399_);
  or (_30707_, _14505_, _13148_);
  and (_30709_, _30707_, _06398_);
  nand (_30710_, _07885_, _07031_);
  and (_30711_, _30710_, _06215_);
  or (_30712_, _30711_, _30709_);
  and (_30713_, _30712_, _30650_);
  or (_30714_, _30713_, _06524_);
  or (_30715_, _30714_, _30706_);
  and (_30716_, _11253_, _07885_);
  or (_30717_, _30716_, _30643_);
  or (_30718_, _30717_, _09030_);
  and (_30720_, _30718_, _07219_);
  and (_30721_, _30720_, _30715_);
  or (_30722_, _14503_, _13148_);
  and (_30723_, _30650_, _06426_);
  and (_30724_, _30723_, _30722_);
  or (_30725_, _30724_, _06532_);
  or (_30726_, _30725_, _30721_);
  and (_30727_, _30656_, _08325_);
  or (_30728_, _30643_, _07217_);
  or (_30729_, _30728_, _30727_);
  and (_30731_, _30729_, _07229_);
  and (_30732_, _30731_, _30726_);
  or (_30733_, _30710_, _08325_);
  and (_30734_, _30650_, _06437_);
  and (_30735_, _30734_, _30733_);
  or (_30736_, _30735_, _06535_);
  or (_30737_, _30736_, _30732_);
  and (_30738_, _30737_, _30646_);
  or (_30739_, _30738_, _06559_);
  or (_30740_, _30654_, _07240_);
  and (_30742_, _30740_, _05933_);
  and (_30743_, _30742_, _30739_);
  and (_30744_, _30678_, _05932_);
  or (_30745_, _30744_, _06566_);
  or (_30746_, _30745_, _30743_);
  or (_30747_, _30643_, _06570_);
  or (_30748_, _30747_, _30651_);
  and (_30749_, _30748_, _01320_);
  and (_30750_, _30749_, _30746_);
  nor (_30751_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_30753_, _30751_, _00000_);
  or (_43010_, _30753_, _30750_);
  and (_30754_, _13148_, \oc8051_golden_model_1.P3 [2]);
  and (_30755_, _07885_, _08662_);
  or (_30756_, _30755_, _30754_);
  or (_30757_, _30756_, _06260_);
  or (_30758_, _30756_, _07169_);
  and (_30759_, _14703_, _07885_);
  or (_30760_, _30759_, _30754_);
  or (_30761_, _30760_, _06286_);
  and (_30763_, _07885_, \oc8051_golden_model_1.ACC [2]);
  or (_30764_, _30763_, _30754_);
  and (_30765_, _30764_, _07143_);
  and (_30766_, _07144_, \oc8051_golden_model_1.P3 [2]);
  or (_30767_, _30766_, _06285_);
  or (_30768_, _30767_, _30765_);
  and (_30769_, _30768_, _06282_);
  and (_30770_, _30769_, _30761_);
  and (_30771_, _13153_, \oc8051_golden_model_1.P3 [2]);
  and (_30772_, _14716_, _08607_);
  or (_30774_, _30772_, _30771_);
  and (_30775_, _30774_, _06281_);
  or (_30776_, _30775_, _06354_);
  or (_30777_, _30776_, _30770_);
  and (_30778_, _30777_, _30758_);
  or (_30779_, _30778_, _06345_);
  or (_30780_, _30764_, _06346_);
  and (_30781_, _30780_, _06278_);
  and (_30782_, _30781_, _30779_);
  and (_30783_, _14699_, _08607_);
  or (_30785_, _30783_, _30771_);
  and (_30786_, _30785_, _06277_);
  or (_30787_, _30786_, _06270_);
  or (_30788_, _30787_, _30782_);
  and (_30789_, _30772_, _14731_);
  or (_30790_, _30771_, _06271_);
  or (_30791_, _30790_, _30789_);
  and (_30792_, _30791_, _06267_);
  and (_30793_, _30792_, _30788_);
  and (_30794_, _14749_, _08607_);
  or (_30796_, _30794_, _30771_);
  and (_30797_, _30796_, _06266_);
  or (_30798_, _30797_, _06259_);
  or (_30799_, _30798_, _30793_);
  and (_30800_, _30799_, _30757_);
  or (_30801_, _30800_, _09486_);
  and (_30802_, _09293_, _07885_);
  or (_30803_, _30754_, _06258_);
  or (_30804_, _30803_, _30802_);
  and (_30805_, _30804_, _06251_);
  and (_30807_, _30805_, _30801_);
  and (_30808_, _14804_, _07885_);
  or (_30809_, _30754_, _30808_);
  and (_30810_, _30809_, _05972_);
  or (_30811_, _30810_, _30807_);
  or (_30812_, _30811_, _10080_);
  and (_30813_, _14697_, _07885_);
  or (_30814_, _30754_, _09025_);
  or (_30815_, _30814_, _30813_);
  and (_30816_, _07885_, _08980_);
  or (_30818_, _30816_, _30754_);
  or (_30819_, _30818_, _06216_);
  and (_30820_, _30819_, _09030_);
  and (_30821_, _30820_, _30815_);
  and (_30822_, _30821_, _30812_);
  and (_30823_, _11250_, _07885_);
  or (_30824_, _30823_, _30754_);
  and (_30825_, _30824_, _06524_);
  or (_30826_, _30825_, _30822_);
  and (_30827_, _30826_, _07219_);
  or (_30829_, _30754_, _08424_);
  and (_30830_, _30818_, _06426_);
  and (_30831_, _30830_, _30829_);
  or (_30832_, _30831_, _30827_);
  and (_30833_, _30832_, _07217_);
  and (_30834_, _30764_, _06532_);
  and (_30835_, _30834_, _30829_);
  or (_30836_, _30835_, _06437_);
  or (_30837_, _30836_, _30833_);
  and (_30838_, _14694_, _07885_);
  or (_30840_, _30754_, _07229_);
  or (_30841_, _30840_, _30838_);
  and (_30842_, _30841_, _07231_);
  and (_30843_, _30842_, _30837_);
  nor (_30844_, _11249_, _13148_);
  or (_30845_, _30844_, _30754_);
  and (_30846_, _30845_, _06535_);
  or (_30847_, _30846_, _06559_);
  or (_30848_, _30847_, _30843_);
  or (_30849_, _30760_, _07240_);
  and (_30851_, _30849_, _05933_);
  and (_30852_, _30851_, _30848_);
  and (_30853_, _30785_, _05932_);
  or (_30854_, _30853_, _06566_);
  or (_30855_, _30854_, _30852_);
  and (_30856_, _14873_, _07885_);
  or (_30857_, _30754_, _06570_);
  or (_30858_, _30857_, _30856_);
  and (_30859_, _30858_, _01320_);
  and (_30860_, _30859_, _30855_);
  nor (_30862_, \oc8051_golden_model_1.P3 [2], rst);
  nor (_30863_, _30862_, _00000_);
  or (_43011_, _30863_, _30860_);
  nor (_30864_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_30865_, _30864_, _00000_);
  and (_30866_, _13148_, \oc8051_golden_model_1.P3 [3]);
  and (_30867_, _07885_, _09421_);
  or (_30868_, _30867_, _30866_);
  or (_30869_, _30868_, _06260_);
  and (_30870_, _14900_, _07885_);
  or (_30872_, _30870_, _30866_);
  or (_30873_, _30872_, _06286_);
  and (_30874_, _07885_, \oc8051_golden_model_1.ACC [3]);
  or (_30875_, _30874_, _30866_);
  and (_30876_, _30875_, _07143_);
  and (_30877_, _07144_, \oc8051_golden_model_1.P3 [3]);
  or (_30878_, _30877_, _06285_);
  or (_30879_, _30878_, _30876_);
  and (_30880_, _30879_, _06282_);
  and (_30881_, _30880_, _30873_);
  and (_30883_, _13153_, \oc8051_golden_model_1.P3 [3]);
  and (_30884_, _14897_, _08607_);
  or (_30885_, _30884_, _30883_);
  and (_30886_, _30885_, _06281_);
  or (_30887_, _30886_, _06354_);
  or (_30888_, _30887_, _30881_);
  or (_30889_, _30868_, _07169_);
  and (_30890_, _30889_, _30888_);
  or (_30891_, _30890_, _06345_);
  or (_30892_, _30875_, _06346_);
  and (_30894_, _30892_, _06278_);
  and (_30895_, _30894_, _30891_);
  and (_30896_, _14895_, _08607_);
  or (_30897_, _30896_, _30883_);
  and (_30898_, _30897_, _06277_);
  or (_30899_, _30898_, _06270_);
  or (_30900_, _30899_, _30895_);
  or (_30901_, _30883_, _14926_);
  and (_30902_, _30901_, _30885_);
  or (_30903_, _30902_, _06271_);
  and (_30905_, _30903_, _06267_);
  and (_30906_, _30905_, _30900_);
  and (_30907_, _14943_, _08607_);
  or (_30908_, _30907_, _30883_);
  and (_30909_, _30908_, _06266_);
  or (_30910_, _30909_, _06259_);
  or (_30911_, _30910_, _30906_);
  and (_30912_, _30911_, _30869_);
  or (_30913_, _30912_, _09486_);
  and (_30914_, _09247_, _07885_);
  or (_30916_, _30866_, _06258_);
  or (_30917_, _30916_, _30914_);
  and (_30918_, _30917_, _06251_);
  and (_30919_, _30918_, _30913_);
  and (_30920_, _14998_, _07885_);
  or (_30921_, _30866_, _30920_);
  and (_30922_, _30921_, _05972_);
  or (_30923_, _30922_, _30919_);
  or (_30924_, _30923_, _10080_);
  and (_30925_, _14893_, _07885_);
  or (_30927_, _30866_, _09025_);
  or (_30928_, _30927_, _30925_);
  and (_30929_, _07885_, _08809_);
  or (_30930_, _30929_, _30866_);
  or (_30931_, _30930_, _06216_);
  and (_30932_, _30931_, _09030_);
  and (_30933_, _30932_, _30928_);
  and (_30934_, _30933_, _30924_);
  and (_30935_, _12529_, _07885_);
  or (_30936_, _30935_, _30866_);
  and (_30938_, _30936_, _06524_);
  or (_30939_, _30938_, _30934_);
  and (_30940_, _30939_, _07219_);
  or (_30941_, _30866_, _08280_);
  and (_30942_, _30930_, _06426_);
  and (_30943_, _30942_, _30941_);
  or (_30944_, _30943_, _30940_);
  and (_30945_, _30944_, _07217_);
  and (_30946_, _30875_, _06532_);
  and (_30947_, _30946_, _30941_);
  or (_30949_, _30947_, _06437_);
  or (_30950_, _30949_, _30945_);
  and (_30951_, _14890_, _07885_);
  or (_30952_, _30866_, _07229_);
  or (_30953_, _30952_, _30951_);
  and (_30954_, _30953_, _07231_);
  and (_30955_, _30954_, _30950_);
  nor (_30956_, _11247_, _13148_);
  or (_30957_, _30956_, _30866_);
  and (_30958_, _30957_, _06535_);
  or (_30960_, _30958_, _06559_);
  or (_30961_, _30960_, _30955_);
  or (_30962_, _30872_, _07240_);
  and (_30963_, _30962_, _05933_);
  and (_30964_, _30963_, _30961_);
  and (_30965_, _30897_, _05932_);
  or (_30966_, _30965_, _06566_);
  or (_30967_, _30966_, _30964_);
  and (_30968_, _15068_, _07885_);
  or (_30969_, _30866_, _06570_);
  or (_30971_, _30969_, _30968_);
  and (_30972_, _30971_, _01320_);
  and (_30973_, _30972_, _30967_);
  or (_43012_, _30973_, _30865_);
  and (_30974_, _13148_, \oc8051_golden_model_1.P3 [4]);
  and (_30975_, _09420_, _07885_);
  or (_30976_, _30975_, _30974_);
  or (_30977_, _30976_, _06260_);
  and (_30978_, _13153_, \oc8051_golden_model_1.P3 [4]);
  and (_30979_, _15145_, _08607_);
  or (_30981_, _30979_, _30978_);
  and (_30982_, _30981_, _06277_);
  and (_30983_, _15133_, _07885_);
  or (_30984_, _30983_, _30974_);
  or (_30985_, _30984_, _06286_);
  and (_30986_, _07885_, \oc8051_golden_model_1.ACC [4]);
  or (_30987_, _30986_, _30974_);
  and (_30988_, _30987_, _07143_);
  and (_30989_, _07144_, \oc8051_golden_model_1.P3 [4]);
  or (_30990_, _30989_, _06285_);
  or (_30992_, _30990_, _30988_);
  and (_30993_, _30992_, _06282_);
  and (_30994_, _30993_, _30985_);
  and (_30995_, _15116_, _08607_);
  or (_30996_, _30995_, _30978_);
  and (_30997_, _30996_, _06281_);
  or (_30998_, _30997_, _06354_);
  or (_30999_, _30998_, _30994_);
  or (_31000_, _30976_, _07169_);
  and (_31001_, _31000_, _30999_);
  or (_31003_, _31001_, _06345_);
  or (_31004_, _30987_, _06346_);
  and (_31005_, _31004_, _06278_);
  and (_31006_, _31005_, _31003_);
  or (_31007_, _31006_, _30982_);
  and (_31008_, _31007_, _06271_);
  and (_31009_, _15153_, _08607_);
  or (_31010_, _31009_, _30978_);
  and (_31011_, _31010_, _06270_);
  or (_31012_, _31011_, _31008_);
  and (_31014_, _31012_, _06267_);
  and (_31015_, _15170_, _08607_);
  or (_31016_, _31015_, _30978_);
  and (_31017_, _31016_, _06266_);
  or (_31018_, _31017_, _06259_);
  or (_31019_, _31018_, _31014_);
  and (_31020_, _31019_, _30977_);
  or (_31021_, _31020_, _09486_);
  and (_31022_, _09437_, _07885_);
  or (_31023_, _30974_, _06258_);
  or (_31025_, _31023_, _31022_);
  and (_31026_, _31025_, _06251_);
  and (_31027_, _31026_, _31021_);
  and (_31028_, _15226_, _07885_);
  or (_31029_, _31028_, _30974_);
  and (_31030_, _31029_, _05972_);
  or (_31031_, _31030_, _10080_);
  or (_31032_, _31031_, _31027_);
  and (_31033_, _15114_, _07885_);
  or (_31034_, _30974_, _09025_);
  or (_31036_, _31034_, _31033_);
  and (_31037_, _08919_, _07885_);
  or (_31038_, _31037_, _30974_);
  or (_31039_, _31038_, _06216_);
  and (_31040_, _31039_, _09030_);
  and (_31041_, _31040_, _31036_);
  and (_31042_, _31041_, _31032_);
  and (_31043_, _11245_, _07885_);
  or (_31044_, _31043_, _30974_);
  and (_31045_, _31044_, _06524_);
  or (_31048_, _31045_, _31042_);
  and (_31049_, _31048_, _07219_);
  or (_31050_, _30974_, _08528_);
  and (_31051_, _31038_, _06426_);
  and (_31052_, _31051_, _31050_);
  or (_31053_, _31052_, _31049_);
  and (_31054_, _31053_, _07217_);
  and (_31055_, _30987_, _06532_);
  and (_31056_, _31055_, _31050_);
  or (_31057_, _31056_, _06437_);
  or (_31059_, _31057_, _31054_);
  and (_31060_, _15111_, _07885_);
  or (_31061_, _30974_, _07229_);
  or (_31062_, _31061_, _31060_);
  and (_31063_, _31062_, _07231_);
  and (_31064_, _31063_, _31059_);
  nor (_31065_, _11244_, _13148_);
  or (_31066_, _31065_, _30974_);
  and (_31067_, _31066_, _06535_);
  or (_31068_, _31067_, _06559_);
  or (_31071_, _31068_, _31064_);
  or (_31072_, _30984_, _07240_);
  and (_31073_, _31072_, _05933_);
  and (_31074_, _31073_, _31071_);
  and (_31075_, _30981_, _05932_);
  or (_31076_, _31075_, _06566_);
  or (_31077_, _31076_, _31074_);
  and (_31078_, _15296_, _07885_);
  or (_31079_, _30974_, _06570_);
  or (_31080_, _31079_, _31078_);
  and (_31082_, _31080_, _01320_);
  and (_31083_, _31082_, _31077_);
  nor (_31084_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_31085_, _31084_, _00000_);
  or (_43013_, _31085_, _31083_);
  nor (_31086_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_31087_, _31086_, _00000_);
  and (_31088_, _13148_, \oc8051_golden_model_1.P3 [5]);
  and (_31089_, _15330_, _07885_);
  or (_31090_, _31089_, _31088_);
  or (_31093_, _31090_, _06286_);
  and (_31094_, _07885_, \oc8051_golden_model_1.ACC [5]);
  or (_31095_, _31094_, _31088_);
  and (_31096_, _31095_, _07143_);
  and (_31097_, _07144_, \oc8051_golden_model_1.P3 [5]);
  or (_31098_, _31097_, _06285_);
  or (_31099_, _31098_, _31096_);
  and (_31100_, _31099_, _06282_);
  and (_31101_, _31100_, _31093_);
  and (_31102_, _13153_, \oc8051_golden_model_1.P3 [5]);
  and (_31104_, _15315_, _08607_);
  or (_31105_, _31104_, _31102_);
  and (_31106_, _31105_, _06281_);
  or (_31107_, _31106_, _06354_);
  or (_31108_, _31107_, _31101_);
  and (_31109_, _09419_, _07885_);
  or (_31110_, _31109_, _31088_);
  or (_31111_, _31110_, _07169_);
  and (_31112_, _31111_, _31108_);
  or (_31113_, _31112_, _06345_);
  or (_31116_, _31095_, _06346_);
  and (_31117_, _31116_, _06278_);
  and (_31118_, _31117_, _31113_);
  and (_31119_, _15342_, _08607_);
  or (_31120_, _31119_, _31102_);
  and (_31121_, _31120_, _06277_);
  or (_31122_, _31121_, _06270_);
  or (_31123_, _31122_, _31118_);
  or (_31124_, _31102_, _15349_);
  and (_31125_, _31124_, _31105_);
  or (_31127_, _31125_, _06271_);
  and (_31128_, _31127_, _06267_);
  and (_31129_, _31128_, _31123_);
  or (_31130_, _31102_, _15365_);
  and (_31131_, _31130_, _06266_);
  and (_31132_, _31131_, _31105_);
  or (_31133_, _31132_, _06259_);
  or (_31134_, _31133_, _31129_);
  or (_31135_, _31110_, _06260_);
  and (_31136_, _31135_, _31134_);
  or (_31138_, _31136_, _09486_);
  and (_31139_, _09436_, _07885_);
  or (_31140_, _31088_, _06258_);
  or (_31141_, _31140_, _31139_);
  and (_31142_, _31141_, _06251_);
  and (_31143_, _31142_, _31138_);
  and (_31144_, _15421_, _07885_);
  or (_31145_, _31144_, _31088_);
  and (_31146_, _31145_, _05972_);
  or (_31147_, _31146_, _10080_);
  or (_31149_, _31147_, _31143_);
  and (_31150_, _15313_, _07885_);
  or (_31151_, _31088_, _09025_);
  or (_31152_, _31151_, _31150_);
  and (_31153_, _08913_, _07885_);
  or (_31154_, _31153_, _31088_);
  or (_31155_, _31154_, _06216_);
  and (_31156_, _31155_, _09030_);
  and (_31157_, _31156_, _31152_);
  and (_31158_, _31157_, _31149_);
  and (_31159_, _12536_, _07885_);
  or (_31160_, _31159_, _31088_);
  and (_31161_, _31160_, _06524_);
  or (_31162_, _31161_, _31158_);
  and (_31163_, _31162_, _07219_);
  or (_31164_, _31088_, _08231_);
  and (_31165_, _31154_, _06426_);
  and (_31166_, _31165_, _31164_);
  or (_31167_, _31166_, _31163_);
  and (_31168_, _31167_, _07217_);
  and (_31171_, _31095_, _06532_);
  and (_31172_, _31171_, _31164_);
  or (_31173_, _31172_, _06437_);
  or (_31174_, _31173_, _31168_);
  and (_31175_, _15310_, _07885_);
  or (_31176_, _31088_, _07229_);
  or (_31177_, _31176_, _31175_);
  and (_31178_, _31177_, _07231_);
  and (_31179_, _31178_, _31174_);
  nor (_31180_, _11241_, _13148_);
  or (_31181_, _31180_, _31088_);
  and (_31182_, _31181_, _06535_);
  or (_31183_, _31182_, _06559_);
  or (_31184_, _31183_, _31179_);
  or (_31185_, _31090_, _07240_);
  and (_31186_, _31185_, _05933_);
  and (_31187_, _31186_, _31184_);
  and (_31188_, _31120_, _05932_);
  or (_31189_, _31188_, _06566_);
  or (_31190_, _31189_, _31187_);
  and (_31193_, _15493_, _07885_);
  or (_31194_, _31088_, _06570_);
  or (_31195_, _31194_, _31193_);
  and (_31196_, _31195_, _01320_);
  and (_31197_, _31196_, _31190_);
  or (_43014_, _31197_, _31087_);
  and (_31198_, _13148_, \oc8051_golden_model_1.P3 [6]);
  and (_31199_, _15521_, _07885_);
  or (_31200_, _31199_, _31198_);
  or (_31201_, _31200_, _06286_);
  and (_31202_, _07885_, \oc8051_golden_model_1.ACC [6]);
  or (_31203_, _31202_, _31198_);
  and (_31204_, _31203_, _07143_);
  and (_31205_, _07144_, \oc8051_golden_model_1.P3 [6]);
  or (_31206_, _31205_, _06285_);
  or (_31207_, _31206_, _31204_);
  and (_31208_, _31207_, _06282_);
  and (_31209_, _31208_, _31201_);
  and (_31210_, _13153_, \oc8051_golden_model_1.P3 [6]);
  and (_31211_, _15535_, _08607_);
  or (_31214_, _31211_, _31210_);
  and (_31215_, _31214_, _06281_);
  or (_31216_, _31215_, _06354_);
  or (_31217_, _31216_, _31209_);
  and (_31218_, _09418_, _07885_);
  or (_31219_, _31218_, _31198_);
  or (_31220_, _31219_, _07169_);
  and (_31221_, _31220_, _31217_);
  or (_31222_, _31221_, _06345_);
  or (_31223_, _31203_, _06346_);
  and (_31224_, _31223_, _06278_);
  and (_31225_, _31224_, _31222_);
  and (_31226_, _15544_, _08607_);
  or (_31227_, _31226_, _31210_);
  and (_31228_, _31227_, _06277_);
  or (_31229_, _31228_, _06270_);
  or (_31230_, _31229_, _31225_);
  or (_31231_, _31210_, _15551_);
  and (_31232_, _31231_, _31214_);
  or (_31233_, _31232_, _06271_);
  and (_31236_, _31233_, _06267_);
  and (_31237_, _31236_, _31230_);
  and (_31238_, _15568_, _08607_);
  or (_31239_, _31238_, _31210_);
  and (_31240_, _31239_, _06266_);
  or (_31241_, _31240_, _06259_);
  or (_31242_, _31241_, _31237_);
  or (_31243_, _31219_, _06260_);
  and (_31244_, _31243_, _31242_);
  or (_31245_, _31244_, _09486_);
  and (_31246_, _09435_, _07885_);
  or (_31247_, _31198_, _06258_);
  or (_31248_, _31247_, _31246_);
  and (_31249_, _31248_, _06251_);
  and (_31250_, _31249_, _31245_);
  and (_31251_, _15623_, _07885_);
  or (_31252_, _31251_, _31198_);
  and (_31253_, _31252_, _05972_);
  or (_31254_, _31253_, _10080_);
  or (_31255_, _31254_, _31250_);
  and (_31258_, _15517_, _07885_);
  or (_31259_, _31198_, _09025_);
  or (_31260_, _31259_, _31258_);
  and (_31261_, _08845_, _07885_);
  or (_31262_, _31261_, _31198_);
  or (_31263_, _31262_, _06216_);
  and (_31264_, _31263_, _09030_);
  and (_31265_, _31264_, _31260_);
  and (_31266_, _31265_, _31255_);
  and (_31267_, _11239_, _07885_);
  or (_31268_, _31267_, _31198_);
  and (_31269_, _31268_, _06524_);
  or (_31270_, _31269_, _31266_);
  and (_31271_, _31270_, _07219_);
  or (_31272_, _31198_, _08128_);
  and (_31273_, _31262_, _06426_);
  and (_31274_, _31273_, _31272_);
  or (_31275_, _31274_, _31271_);
  and (_31276_, _31275_, _07217_);
  and (_31277_, _31203_, _06532_);
  and (_31280_, _31277_, _31272_);
  or (_31281_, _31280_, _06437_);
  or (_31282_, _31281_, _31276_);
  and (_31283_, _15514_, _07885_);
  or (_31284_, _31198_, _07229_);
  or (_31285_, _31284_, _31283_);
  and (_31286_, _31285_, _07231_);
  and (_31287_, _31286_, _31282_);
  nor (_31288_, _11238_, _13148_);
  or (_31289_, _31288_, _31198_);
  and (_31290_, _31289_, _06535_);
  or (_31291_, _31290_, _06559_);
  or (_31292_, _31291_, _31287_);
  or (_31293_, _31200_, _07240_);
  and (_31294_, _31293_, _05933_);
  and (_31295_, _31294_, _31292_);
  and (_31296_, _31227_, _05932_);
  or (_31297_, _31296_, _06566_);
  or (_31298_, _31297_, _31295_);
  and (_31299_, _15695_, _07885_);
  or (_31302_, _31198_, _06570_);
  or (_31303_, _31302_, _31299_);
  and (_31304_, _31303_, _01320_);
  and (_31305_, _31304_, _31298_);
  nor (_31306_, \oc8051_golden_model_1.P3 [6], rst);
  nor (_31307_, _31306_, _00000_);
  or (_43015_, _31307_, _31305_);
  nand (_31308_, _11254_, _07946_);
  not (_31309_, \oc8051_golden_model_1.P0 [0]);
  nor (_31310_, _07946_, _31309_);
  nor (_31311_, _31310_, _07217_);
  nand (_31312_, _31311_, _31308_);
  and (_31313_, _07946_, _07135_);
  or (_31314_, _31313_, _31310_);
  or (_31315_, _31314_, _06260_);
  nor (_31316_, _08374_, _13250_);
  or (_31317_, _31316_, _31310_);
  or (_31318_, _31317_, _06286_);
  and (_31319_, _07946_, \oc8051_golden_model_1.ACC [0]);
  or (_31320_, _31319_, _31310_);
  and (_31323_, _31320_, _07143_);
  nor (_31324_, _07143_, _31309_);
  or (_31325_, _31324_, _06285_);
  or (_31326_, _31325_, _31323_);
  and (_31327_, _31326_, _06282_);
  and (_31328_, _31327_, _31318_);
  nor (_31329_, _07939_, _31309_);
  and (_31330_, _14326_, _07939_);
  or (_31331_, _31330_, _31329_);
  and (_31332_, _31331_, _06281_);
  or (_31333_, _31332_, _31328_);
  and (_31334_, _31333_, _07169_);
  and (_31335_, _31314_, _06354_);
  or (_31336_, _31335_, _06345_);
  or (_31337_, _31336_, _31334_);
  or (_31338_, _31320_, _06346_);
  and (_31339_, _31338_, _06278_);
  and (_31340_, _31339_, _31337_);
  and (_31341_, _31310_, _06277_);
  or (_31342_, _31341_, _06270_);
  or (_31345_, _31342_, _31340_);
  or (_31346_, _31317_, _06271_);
  and (_31347_, _31346_, _06267_);
  and (_31348_, _31347_, _31345_);
  and (_31349_, _14358_, _07939_);
  or (_31350_, _31349_, _31329_);
  and (_31351_, _31350_, _06266_);
  or (_31352_, _31351_, _06259_);
  or (_31353_, _31352_, _31348_);
  and (_31354_, _31353_, _31315_);
  or (_31355_, _31354_, _09486_);
  and (_31356_, _09384_, _07946_);
  or (_31357_, _31310_, _06258_);
  or (_31358_, _31357_, _31356_);
  and (_31359_, _31358_, _06251_);
  and (_31360_, _31359_, _31355_);
  and (_31361_, _14413_, _07946_);
  or (_31362_, _31361_, _31310_);
  and (_31363_, _31362_, _05972_);
  or (_31364_, _31363_, _31360_);
  or (_31367_, _31364_, _10080_);
  and (_31368_, _14311_, _07946_);
  or (_31369_, _31310_, _09025_);
  or (_31370_, _31369_, _31368_);
  and (_31371_, _07946_, _08929_);
  or (_31372_, _31371_, _31310_);
  or (_31373_, _31372_, _06216_);
  and (_31374_, _31373_, _09030_);
  and (_31375_, _31374_, _31370_);
  and (_31376_, _31375_, _31367_);
  nor (_31377_, _12532_, _13250_);
  or (_31378_, _31377_, _31310_);
  and (_31379_, _31308_, _06524_);
  and (_31380_, _31379_, _31378_);
  or (_31381_, _31380_, _31376_);
  and (_31382_, _31381_, _07219_);
  nand (_31383_, _31372_, _06426_);
  nor (_31384_, _31383_, _31316_);
  or (_31385_, _31384_, _06532_);
  or (_31386_, _31385_, _31382_);
  and (_31389_, _31386_, _31312_);
  or (_31390_, _31389_, _06437_);
  and (_31391_, _14307_, _07946_);
  or (_31392_, _31391_, _31310_);
  or (_31393_, _31392_, _07229_);
  and (_31394_, _31393_, _07231_);
  and (_31395_, _31394_, _31390_);
  and (_31396_, _31378_, _06535_);
  or (_31397_, _31396_, _06559_);
  or (_31398_, _31397_, _31395_);
  or (_31399_, _31317_, _07240_);
  and (_31400_, _31399_, _31398_);
  or (_31401_, _31400_, _05932_);
  or (_31402_, _31310_, _05933_);
  and (_31403_, _31402_, _31401_);
  or (_31404_, _31403_, _06566_);
  or (_31405_, _31317_, _06570_);
  and (_31406_, _31405_, _01320_);
  and (_31407_, _31406_, _31404_);
  nor (_31408_, \oc8051_golden_model_1.P0 [0], rst);
  nor (_31411_, _31408_, _00000_);
  or (_43017_, _31411_, _31407_);
  not (_31412_, \oc8051_golden_model_1.P0 [1]);
  nor (_31413_, _07946_, _31412_);
  nor (_31414_, _11252_, _13250_);
  or (_31415_, _31414_, _31413_);
  or (_31416_, _31415_, _07231_);
  and (_31417_, _07946_, _09422_);
  or (_31418_, _31417_, _31413_);
  or (_31419_, _31418_, _07169_);
  or (_31420_, _07946_, \oc8051_golden_model_1.P0 [1]);
  and (_31421_, _14520_, _07946_);
  not (_31422_, _31421_);
  and (_31423_, _31422_, _31420_);
  or (_31424_, _31423_, _06286_);
  and (_31425_, _07946_, \oc8051_golden_model_1.ACC [1]);
  or (_31426_, _31425_, _31413_);
  and (_31427_, _31426_, _07143_);
  nor (_31428_, _07143_, _31412_);
  or (_31429_, _31428_, _06285_);
  or (_31432_, _31429_, _31427_);
  and (_31433_, _31432_, _06282_);
  and (_31434_, _31433_, _31424_);
  nor (_31435_, _07939_, _31412_);
  and (_31436_, _14508_, _07939_);
  or (_31437_, _31436_, _31435_);
  and (_31438_, _31437_, _06281_);
  or (_31439_, _31438_, _06354_);
  or (_31440_, _31439_, _31434_);
  and (_31441_, _31440_, _31419_);
  or (_31442_, _31441_, _06345_);
  or (_31443_, _31426_, _06346_);
  and (_31444_, _31443_, _06278_);
  and (_31445_, _31444_, _31442_);
  and (_31446_, _14511_, _07939_);
  or (_31447_, _31446_, _31435_);
  and (_31448_, _31447_, _06277_);
  or (_31449_, _31448_, _06270_);
  or (_31450_, _31449_, _31445_);
  and (_31451_, _31436_, _14507_);
  or (_31454_, _31435_, _06271_);
  or (_31455_, _31454_, _31451_);
  and (_31456_, _31455_, _06267_);
  and (_31457_, _31456_, _31450_);
  or (_31458_, _31435_, _14551_);
  and (_31459_, _31458_, _06266_);
  and (_31460_, _31459_, _31437_);
  or (_31461_, _31460_, _06259_);
  or (_31462_, _31461_, _31457_);
  or (_31463_, _31418_, _06260_);
  and (_31464_, _31463_, _31462_);
  or (_31465_, _31464_, _09486_);
  and (_31466_, _09339_, _07946_);
  or (_31467_, _31413_, _06258_);
  or (_31468_, _31467_, _31466_);
  and (_31469_, _31468_, _06251_);
  and (_31470_, _31469_, _31465_);
  and (_31471_, _14607_, _07946_);
  or (_31472_, _31471_, _31413_);
  and (_31473_, _31472_, _05972_);
  or (_31476_, _31473_, _31470_);
  and (_31477_, _31476_, _06399_);
  or (_31478_, _14505_, _13250_);
  and (_31479_, _31478_, _06398_);
  nand (_31480_, _07946_, _07031_);
  and (_31481_, _31480_, _06215_);
  or (_31482_, _31481_, _31479_);
  and (_31483_, _31482_, _31420_);
  or (_31484_, _31483_, _06524_);
  or (_31485_, _31484_, _31477_);
  nand (_31486_, _11251_, _07946_);
  and (_31487_, _31486_, _31415_);
  or (_31488_, _31487_, _09030_);
  and (_31489_, _31488_, _07219_);
  and (_31490_, _31489_, _31485_);
  or (_31491_, _14503_, _13250_);
  and (_31492_, _31420_, _06426_);
  and (_31493_, _31492_, _31491_);
  or (_31494_, _31493_, _06532_);
  or (_31495_, _31494_, _31490_);
  nor (_31498_, _31413_, _07217_);
  nand (_31499_, _31498_, _31486_);
  and (_31500_, _31499_, _07229_);
  and (_31501_, _31500_, _31495_);
  or (_31502_, _31480_, _08325_);
  and (_31503_, _31420_, _06437_);
  and (_31504_, _31503_, _31502_);
  or (_31505_, _31504_, _06535_);
  or (_31506_, _31505_, _31501_);
  and (_31507_, _31506_, _31416_);
  or (_31508_, _31507_, _06559_);
  or (_31509_, _31423_, _07240_);
  and (_31510_, _31509_, _05933_);
  and (_31511_, _31510_, _31508_);
  and (_31512_, _31447_, _05932_);
  or (_31513_, _31512_, _06566_);
  or (_31514_, _31513_, _31511_);
  or (_31515_, _31413_, _06570_);
  or (_31516_, _31515_, _31421_);
  and (_31517_, _31516_, _01320_);
  and (_31520_, _31517_, _31514_);
  nor (_31521_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_31522_, _31521_, _00000_);
  or (_43018_, _31522_, _31520_);
  and (_31523_, _13250_, \oc8051_golden_model_1.P0 [2]);
  and (_31524_, _07946_, _08662_);
  or (_31525_, _31524_, _31523_);
  or (_31526_, _31525_, _06260_);
  or (_31527_, _31525_, _07169_);
  and (_31528_, _14703_, _07946_);
  or (_31529_, _31528_, _31523_);
  or (_31530_, _31529_, _06286_);
  and (_31531_, _07946_, \oc8051_golden_model_1.ACC [2]);
  or (_31532_, _31531_, _31523_);
  and (_31533_, _31532_, _07143_);
  and (_31534_, _07144_, \oc8051_golden_model_1.P0 [2]);
  or (_31535_, _31534_, _06285_);
  or (_31536_, _31535_, _31533_);
  and (_31537_, _31536_, _06282_);
  and (_31538_, _31537_, _31530_);
  and (_31541_, _13255_, \oc8051_golden_model_1.P0 [2]);
  and (_31542_, _14716_, _07939_);
  or (_31543_, _31542_, _31541_);
  and (_31544_, _31543_, _06281_);
  or (_31545_, _31544_, _06354_);
  or (_31546_, _31545_, _31538_);
  and (_31547_, _31546_, _31527_);
  or (_31548_, _31547_, _06345_);
  or (_31549_, _31532_, _06346_);
  and (_31550_, _31549_, _06278_);
  and (_31551_, _31550_, _31548_);
  and (_31552_, _14699_, _07939_);
  or (_31553_, _31552_, _31541_);
  and (_31554_, _31553_, _06277_);
  or (_31555_, _31554_, _06270_);
  or (_31556_, _31555_, _31551_);
  and (_31557_, _31542_, _14731_);
  or (_31558_, _31541_, _06271_);
  or (_31559_, _31558_, _31557_);
  and (_31560_, _31559_, _06267_);
  and (_31563_, _31560_, _31556_);
  and (_31564_, _14749_, _07939_);
  or (_31565_, _31564_, _31541_);
  and (_31566_, _31565_, _06266_);
  or (_31567_, _31566_, _06259_);
  or (_31568_, _31567_, _31563_);
  and (_31569_, _31568_, _31526_);
  or (_31570_, _31569_, _09486_);
  and (_31571_, _09293_, _07946_);
  or (_31572_, _31523_, _06258_);
  or (_31573_, _31572_, _31571_);
  and (_31574_, _31573_, _06251_);
  and (_31575_, _31574_, _31570_);
  and (_31576_, _14804_, _07946_);
  or (_31577_, _31523_, _31576_);
  and (_31578_, _31577_, _05972_);
  or (_31579_, _31578_, _31575_);
  or (_31580_, _31579_, _10080_);
  and (_31581_, _14697_, _07946_);
  or (_31582_, _31523_, _09025_);
  or (_31585_, _31582_, _31581_);
  and (_31586_, _07946_, _08980_);
  or (_31587_, _31586_, _31523_);
  or (_31588_, _31587_, _06216_);
  and (_31589_, _31588_, _09030_);
  and (_31590_, _31589_, _31585_);
  and (_31591_, _31590_, _31580_);
  and (_31592_, _11250_, _07946_);
  or (_31593_, _31592_, _31523_);
  and (_31594_, _31593_, _06524_);
  or (_31595_, _31594_, _31591_);
  and (_31596_, _31595_, _07219_);
  or (_31597_, _31523_, _08424_);
  and (_31598_, _31587_, _06426_);
  and (_31599_, _31598_, _31597_);
  or (_31600_, _31599_, _31596_);
  and (_31601_, _31600_, _07217_);
  and (_31602_, _31532_, _06532_);
  and (_31603_, _31602_, _31597_);
  or (_31604_, _31603_, _06437_);
  or (_31607_, _31604_, _31601_);
  and (_31608_, _14694_, _07946_);
  or (_31609_, _31523_, _07229_);
  or (_31610_, _31609_, _31608_);
  and (_31611_, _31610_, _07231_);
  and (_31612_, _31611_, _31607_);
  nor (_31613_, _11249_, _13250_);
  or (_31614_, _31613_, _31523_);
  and (_31615_, _31614_, _06535_);
  or (_31616_, _31615_, _06559_);
  or (_31617_, _31616_, _31612_);
  or (_31618_, _31529_, _07240_);
  and (_31619_, _31618_, _05933_);
  and (_31620_, _31619_, _31617_);
  and (_31621_, _31553_, _05932_);
  or (_31622_, _31621_, _06566_);
  or (_31623_, _31622_, _31620_);
  and (_31624_, _14873_, _07946_);
  or (_31625_, _31523_, _06570_);
  or (_31626_, _31625_, _31624_);
  and (_31629_, _31626_, _01320_);
  and (_31630_, _31629_, _31623_);
  nor (_31631_, \oc8051_golden_model_1.P0 [2], rst);
  nor (_31632_, _31631_, _00000_);
  or (_43019_, _31632_, _31630_);
  and (_31633_, _13250_, \oc8051_golden_model_1.P0 [3]);
  and (_31634_, _07946_, _09421_);
  or (_31635_, _31634_, _31633_);
  or (_31636_, _31635_, _06260_);
  and (_31637_, _14900_, _07946_);
  or (_31638_, _31637_, _31633_);
  or (_31639_, _31638_, _06286_);
  and (_31640_, _07946_, \oc8051_golden_model_1.ACC [3]);
  or (_31641_, _31640_, _31633_);
  and (_31642_, _31641_, _07143_);
  and (_31643_, _07144_, \oc8051_golden_model_1.P0 [3]);
  or (_31644_, _31643_, _06285_);
  or (_31645_, _31644_, _31642_);
  and (_31646_, _31645_, _06282_);
  and (_31647_, _31646_, _31639_);
  and (_31650_, _13255_, \oc8051_golden_model_1.P0 [3]);
  and (_31651_, _14897_, _07939_);
  or (_31652_, _31651_, _31650_);
  and (_31653_, _31652_, _06281_);
  or (_31654_, _31653_, _06354_);
  or (_31655_, _31654_, _31647_);
  or (_31656_, _31635_, _07169_);
  and (_31657_, _31656_, _31655_);
  or (_31658_, _31657_, _06345_);
  or (_31659_, _31641_, _06346_);
  and (_31660_, _31659_, _06278_);
  and (_31661_, _31660_, _31658_);
  and (_31662_, _14895_, _07939_);
  or (_31663_, _31662_, _31650_);
  and (_31664_, _31663_, _06277_);
  or (_31665_, _31664_, _06270_);
  or (_31666_, _31665_, _31661_);
  or (_31667_, _31650_, _14926_);
  and (_31668_, _31667_, _31652_);
  or (_31669_, _31668_, _06271_);
  and (_31672_, _31669_, _06267_);
  and (_31673_, _31672_, _31666_);
  and (_31674_, _14943_, _07939_);
  or (_31675_, _31674_, _31650_);
  and (_31676_, _31675_, _06266_);
  or (_31677_, _31676_, _06259_);
  or (_31678_, _31677_, _31673_);
  and (_31679_, _31678_, _31636_);
  or (_31680_, _31679_, _09486_);
  and (_31681_, _09247_, _07946_);
  or (_31682_, _31633_, _06258_);
  or (_31683_, _31682_, _31681_);
  and (_31684_, _31683_, _06251_);
  and (_31685_, _31684_, _31680_);
  and (_31686_, _14998_, _07946_);
  or (_31687_, _31633_, _31686_);
  and (_31688_, _31687_, _05972_);
  or (_31689_, _31688_, _31685_);
  or (_31690_, _31689_, _10080_);
  and (_31691_, _14893_, _07946_);
  or (_31694_, _31633_, _09025_);
  or (_31695_, _31694_, _31691_);
  and (_31696_, _07946_, _08809_);
  or (_31697_, _31696_, _31633_);
  or (_31698_, _31697_, _06216_);
  and (_31699_, _31698_, _09030_);
  and (_31700_, _31699_, _31695_);
  and (_31701_, _31700_, _31690_);
  and (_31702_, _12529_, _07946_);
  or (_31703_, _31702_, _31633_);
  and (_31704_, _31703_, _06524_);
  or (_31705_, _31704_, _31701_);
  and (_31706_, _31705_, _07219_);
  or (_31707_, _31633_, _08280_);
  and (_31708_, _31697_, _06426_);
  and (_31709_, _31708_, _31707_);
  or (_31710_, _31709_, _31706_);
  and (_31711_, _31710_, _07217_);
  and (_31712_, _31641_, _06532_);
  and (_31713_, _31712_, _31707_);
  or (_31716_, _31713_, _06437_);
  or (_31717_, _31716_, _31711_);
  and (_31718_, _14890_, _07946_);
  or (_31719_, _31633_, _07229_);
  or (_31720_, _31719_, _31718_);
  and (_31721_, _31720_, _07231_);
  and (_31722_, _31721_, _31717_);
  nor (_31723_, _11247_, _13250_);
  or (_31724_, _31723_, _31633_);
  and (_31725_, _31724_, _06535_);
  or (_31726_, _31725_, _06559_);
  or (_31727_, _31726_, _31722_);
  or (_31728_, _31638_, _07240_);
  and (_31729_, _31728_, _05933_);
  and (_31730_, _31729_, _31727_);
  and (_31731_, _31663_, _05932_);
  or (_31732_, _31731_, _06566_);
  or (_31733_, _31732_, _31730_);
  and (_31734_, _15068_, _07946_);
  or (_31735_, _31633_, _06570_);
  or (_31738_, _31735_, _31734_);
  and (_31739_, _31738_, _01320_);
  and (_31740_, _31739_, _31733_);
  nor (_31741_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_31742_, _31741_, _00000_);
  or (_43021_, _31742_, _31740_);
  nor (_31743_, \oc8051_golden_model_1.P0 [4], rst);
  nor (_31744_, _31743_, _00000_);
  and (_31745_, _13250_, \oc8051_golden_model_1.P0 [4]);
  and (_31746_, _09420_, _07946_);
  or (_31747_, _31746_, _31745_);
  or (_31748_, _31747_, _06260_);
  and (_31749_, _13255_, \oc8051_golden_model_1.P0 [4]);
  and (_31750_, _15145_, _07939_);
  or (_31751_, _31750_, _31749_);
  and (_31752_, _31751_, _06277_);
  and (_31753_, _15133_, _07946_);
  or (_31754_, _31753_, _31745_);
  or (_31755_, _31754_, _06286_);
  and (_31756_, _07946_, \oc8051_golden_model_1.ACC [4]);
  or (_31759_, _31756_, _31745_);
  and (_31760_, _31759_, _07143_);
  and (_31761_, _07144_, \oc8051_golden_model_1.P0 [4]);
  or (_31762_, _31761_, _06285_);
  or (_31763_, _31762_, _31760_);
  and (_31764_, _31763_, _06282_);
  and (_31765_, _31764_, _31755_);
  and (_31766_, _15116_, _07939_);
  or (_31767_, _31766_, _31749_);
  and (_31768_, _31767_, _06281_);
  or (_31770_, _31768_, _06354_);
  or (_31771_, _31770_, _31765_);
  or (_31772_, _31747_, _07169_);
  and (_31773_, _31772_, _31771_);
  or (_31774_, _31773_, _06345_);
  or (_31775_, _31759_, _06346_);
  and (_31776_, _31775_, _06278_);
  and (_31777_, _31776_, _31774_);
  or (_31778_, _31777_, _31752_);
  and (_31779_, _31778_, _06271_);
  and (_31781_, _15153_, _07939_);
  or (_31782_, _31781_, _31749_);
  and (_31783_, _31782_, _06270_);
  or (_31784_, _31783_, _31779_);
  and (_31785_, _31784_, _06267_);
  and (_31786_, _15170_, _07939_);
  or (_31787_, _31786_, _31749_);
  and (_31788_, _31787_, _06266_);
  or (_31789_, _31788_, _06259_);
  or (_31790_, _31789_, _31785_);
  and (_31792_, _31790_, _31748_);
  or (_31793_, _31792_, _09486_);
  and (_31794_, _09437_, _07946_);
  or (_31795_, _31745_, _06258_);
  or (_31796_, _31795_, _31794_);
  and (_31797_, _31796_, _06251_);
  and (_31798_, _31797_, _31793_);
  and (_31799_, _15226_, _07946_);
  or (_31800_, _31799_, _31745_);
  and (_31801_, _31800_, _05972_);
  or (_31803_, _31801_, _10080_);
  or (_31804_, _31803_, _31798_);
  and (_31805_, _15114_, _07946_);
  or (_31806_, _31745_, _09025_);
  or (_31807_, _31806_, _31805_);
  and (_31808_, _08919_, _07946_);
  or (_31809_, _31808_, _31745_);
  or (_31810_, _31809_, _06216_);
  and (_31811_, _31810_, _09030_);
  and (_31812_, _31811_, _31807_);
  and (_31814_, _31812_, _31804_);
  and (_31815_, _11245_, _07946_);
  or (_31816_, _31815_, _31745_);
  and (_31817_, _31816_, _06524_);
  or (_31818_, _31817_, _31814_);
  and (_31819_, _31818_, _07219_);
  or (_31820_, _31745_, _08528_);
  and (_31821_, _31809_, _06426_);
  and (_31822_, _31821_, _31820_);
  or (_31823_, _31822_, _31819_);
  and (_31825_, _31823_, _07217_);
  and (_31826_, _31759_, _06532_);
  and (_31827_, _31826_, _31820_);
  or (_31828_, _31827_, _06437_);
  or (_31829_, _31828_, _31825_);
  and (_31830_, _15111_, _07946_);
  or (_31831_, _31745_, _07229_);
  or (_31832_, _31831_, _31830_);
  and (_31833_, _31832_, _07231_);
  and (_31834_, _31833_, _31829_);
  nor (_31836_, _11244_, _13250_);
  or (_31837_, _31836_, _31745_);
  and (_31838_, _31837_, _06535_);
  or (_31839_, _31838_, _06559_);
  or (_31840_, _31839_, _31834_);
  or (_31841_, _31754_, _07240_);
  and (_31842_, _31841_, _05933_);
  and (_31843_, _31842_, _31840_);
  and (_31844_, _31751_, _05932_);
  or (_31845_, _31844_, _06566_);
  or (_31847_, _31845_, _31843_);
  and (_31848_, _15296_, _07946_);
  or (_31849_, _31745_, _06570_);
  or (_31850_, _31849_, _31848_);
  and (_31851_, _31850_, _01320_);
  and (_31852_, _31851_, _31847_);
  or (_43022_, _31852_, _31744_);
  and (_31853_, _13250_, \oc8051_golden_model_1.P0 [5]);
  and (_31854_, _15330_, _07946_);
  or (_31855_, _31854_, _31853_);
  or (_31857_, _31855_, _06286_);
  and (_31858_, _07946_, \oc8051_golden_model_1.ACC [5]);
  or (_31859_, _31858_, _31853_);
  and (_31860_, _31859_, _07143_);
  and (_31861_, _07144_, \oc8051_golden_model_1.P0 [5]);
  or (_31862_, _31861_, _06285_);
  or (_31863_, _31862_, _31860_);
  and (_31864_, _31863_, _06282_);
  and (_31865_, _31864_, _31857_);
  and (_31866_, _13255_, \oc8051_golden_model_1.P0 [5]);
  and (_31868_, _15315_, _07939_);
  or (_31869_, _31868_, _31866_);
  and (_31870_, _31869_, _06281_);
  or (_31871_, _31870_, _06354_);
  or (_31872_, _31871_, _31865_);
  and (_31873_, _09419_, _07946_);
  or (_31874_, _31873_, _31853_);
  or (_31875_, _31874_, _07169_);
  and (_31876_, _31875_, _31872_);
  or (_31877_, _31876_, _06345_);
  or (_31879_, _31859_, _06346_);
  and (_31880_, _31879_, _06278_);
  and (_31881_, _31880_, _31877_);
  and (_31882_, _15342_, _07939_);
  or (_31883_, _31882_, _31866_);
  and (_31884_, _31883_, _06277_);
  or (_31885_, _31884_, _06270_);
  or (_31886_, _31885_, _31881_);
  or (_31887_, _31866_, _15349_);
  and (_31888_, _31887_, _31869_);
  or (_31890_, _31888_, _06271_);
  and (_31891_, _31890_, _06267_);
  and (_31892_, _31891_, _31886_);
  or (_31893_, _31866_, _15365_);
  and (_31894_, _31893_, _06266_);
  and (_31895_, _31894_, _31869_);
  or (_31896_, _31895_, _06259_);
  or (_31897_, _31896_, _31892_);
  or (_31898_, _31874_, _06260_);
  and (_31899_, _31898_, _31897_);
  or (_31901_, _31899_, _09486_);
  and (_31902_, _09436_, _07946_);
  or (_31903_, _31853_, _06258_);
  or (_31904_, _31903_, _31902_);
  and (_31905_, _31904_, _06251_);
  and (_31906_, _31905_, _31901_);
  and (_31907_, _15421_, _07946_);
  or (_31908_, _31907_, _31853_);
  and (_31909_, _31908_, _05972_);
  or (_31910_, _31909_, _10080_);
  or (_31912_, _31910_, _31906_);
  and (_31913_, _15313_, _07946_);
  or (_31914_, _31853_, _09025_);
  or (_31915_, _31914_, _31913_);
  and (_31916_, _08913_, _07946_);
  or (_31917_, _31916_, _31853_);
  or (_31918_, _31917_, _06216_);
  and (_31919_, _31918_, _09030_);
  and (_31920_, _31919_, _31915_);
  and (_31921_, _31920_, _31912_);
  and (_31923_, _12536_, _07946_);
  or (_31924_, _31923_, _31853_);
  and (_31925_, _31924_, _06524_);
  or (_31926_, _31925_, _31921_);
  and (_31927_, _31926_, _07219_);
  or (_31928_, _31853_, _08231_);
  and (_31929_, _31917_, _06426_);
  and (_31930_, _31929_, _31928_);
  or (_31931_, _31930_, _31927_);
  and (_31932_, _31931_, _07217_);
  and (_31934_, _31859_, _06532_);
  and (_31935_, _31934_, _31928_);
  or (_31936_, _31935_, _06437_);
  or (_31937_, _31936_, _31932_);
  and (_31938_, _15310_, _07946_);
  or (_31939_, _31853_, _07229_);
  or (_31940_, _31939_, _31938_);
  and (_31941_, _31940_, _07231_);
  and (_31942_, _31941_, _31937_);
  nor (_31943_, _11241_, _13250_);
  or (_31945_, _31943_, _31853_);
  and (_31946_, _31945_, _06535_);
  or (_31947_, _31946_, _06559_);
  or (_31948_, _31947_, _31942_);
  or (_31949_, _31855_, _07240_);
  and (_31950_, _31949_, _05933_);
  and (_31951_, _31950_, _31948_);
  and (_31952_, _31883_, _05932_);
  or (_31953_, _31952_, _06566_);
  or (_31954_, _31953_, _31951_);
  and (_31956_, _15493_, _07946_);
  or (_31957_, _31853_, _06570_);
  or (_31958_, _31957_, _31956_);
  and (_31959_, _31958_, _01320_);
  and (_31960_, _31959_, _31954_);
  nor (_31961_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_31962_, _31961_, _00000_);
  or (_43023_, _31962_, _31960_);
  and (_31963_, _13250_, \oc8051_golden_model_1.P0 [6]);
  and (_31964_, _15521_, _07946_);
  or (_31966_, _31964_, _31963_);
  or (_31967_, _31966_, _06286_);
  and (_31968_, _07946_, \oc8051_golden_model_1.ACC [6]);
  or (_31969_, _31968_, _31963_);
  and (_31970_, _31969_, _07143_);
  and (_31971_, _07144_, \oc8051_golden_model_1.P0 [6]);
  or (_31972_, _31971_, _06285_);
  or (_31973_, _31972_, _31970_);
  and (_31974_, _31973_, _06282_);
  and (_31975_, _31974_, _31967_);
  and (_31977_, _13255_, \oc8051_golden_model_1.P0 [6]);
  and (_31978_, _15535_, _07939_);
  or (_31979_, _31978_, _31977_);
  and (_31980_, _31979_, _06281_);
  or (_31981_, _31980_, _06354_);
  or (_31982_, _31981_, _31975_);
  and (_31983_, _09418_, _07946_);
  or (_31984_, _31983_, _31963_);
  or (_31985_, _31984_, _07169_);
  and (_31986_, _31985_, _31982_);
  or (_31988_, _31986_, _06345_);
  or (_31989_, _31969_, _06346_);
  and (_31990_, _31989_, _06278_);
  and (_31991_, _31990_, _31988_);
  and (_31992_, _15544_, _07939_);
  or (_31993_, _31992_, _31977_);
  and (_31994_, _31993_, _06277_);
  or (_31995_, _31994_, _06270_);
  or (_31996_, _31995_, _31991_);
  or (_31997_, _31977_, _15551_);
  and (_31999_, _31997_, _31979_);
  or (_32000_, _31999_, _06271_);
  and (_32001_, _32000_, _06267_);
  and (_32002_, _32001_, _31996_);
  and (_32003_, _15568_, _07939_);
  or (_32004_, _32003_, _31977_);
  and (_32005_, _32004_, _06266_);
  or (_32006_, _32005_, _06259_);
  or (_32007_, _32006_, _32002_);
  or (_32008_, _31984_, _06260_);
  and (_32010_, _32008_, _32007_);
  or (_32011_, _32010_, _09486_);
  and (_32012_, _09435_, _07946_);
  or (_32013_, _31963_, _06258_);
  or (_32014_, _32013_, _32012_);
  and (_32015_, _32014_, _06251_);
  and (_32016_, _32015_, _32011_);
  and (_32017_, _15623_, _07946_);
  or (_32018_, _32017_, _31963_);
  and (_32019_, _32018_, _05972_);
  or (_32020_, _32019_, _10080_);
  or (_32021_, _32020_, _32016_);
  and (_32022_, _15517_, _07946_);
  or (_32023_, _31963_, _09025_);
  or (_32024_, _32023_, _32022_);
  and (_32025_, _08845_, _07946_);
  or (_32026_, _32025_, _31963_);
  or (_32027_, _32026_, _06216_);
  and (_32028_, _32027_, _09030_);
  and (_32029_, _32028_, _32024_);
  and (_32031_, _32029_, _32021_);
  and (_32032_, _11239_, _07946_);
  or (_32033_, _32032_, _31963_);
  and (_32034_, _32033_, _06524_);
  or (_32035_, _32034_, _32031_);
  and (_32036_, _32035_, _07219_);
  or (_32037_, _31963_, _08128_);
  and (_32038_, _32026_, _06426_);
  and (_32039_, _32038_, _32037_);
  or (_32040_, _32039_, _32036_);
  and (_32042_, _32040_, _07217_);
  and (_32043_, _31969_, _06532_);
  and (_32044_, _32043_, _32037_);
  or (_32045_, _32044_, _06437_);
  or (_32046_, _32045_, _32042_);
  and (_32047_, _15514_, _07946_);
  or (_32048_, _31963_, _07229_);
  or (_32049_, _32048_, _32047_);
  and (_32050_, _32049_, _07231_);
  and (_32051_, _32050_, _32046_);
  nor (_32053_, _11238_, _13250_);
  or (_32054_, _32053_, _31963_);
  and (_32055_, _32054_, _06535_);
  or (_32056_, _32055_, _06559_);
  or (_32057_, _32056_, _32051_);
  or (_32058_, _31966_, _07240_);
  and (_32059_, _32058_, _05933_);
  and (_32060_, _32059_, _32057_);
  and (_32061_, _31993_, _05932_);
  or (_32062_, _32061_, _06566_);
  or (_32064_, _32062_, _32060_);
  and (_32065_, _15695_, _07946_);
  or (_32066_, _31963_, _06570_);
  or (_32067_, _32066_, _32065_);
  and (_32068_, _32067_, _01320_);
  and (_32069_, _32068_, _32064_);
  nor (_32070_, \oc8051_golden_model_1.P0 [6], rst);
  nor (_32071_, _32070_, _00000_);
  or (_43024_, _32071_, _32069_);
  nor (_32072_, \oc8051_golden_model_1.P1 [0], rst);
  nor (_32074_, _32072_, _00000_);
  nand (_32075_, _11254_, _07961_);
  and (_32076_, _13354_, \oc8051_golden_model_1.P1 [0]);
  nor (_32077_, _32076_, _07217_);
  nand (_32078_, _32077_, _32075_);
  and (_32079_, _07961_, _07135_);
  or (_32080_, _32079_, _32076_);
  or (_32081_, _32080_, _06260_);
  nor (_32082_, _08374_, _13354_);
  or (_32083_, _32082_, _32076_);
  or (_32085_, _32083_, _06286_);
  and (_32086_, _07961_, \oc8051_golden_model_1.ACC [0]);
  or (_32087_, _32086_, _32076_);
  and (_32088_, _32087_, _07143_);
  and (_32089_, _07144_, \oc8051_golden_model_1.P1 [0]);
  or (_32090_, _32089_, _06285_);
  or (_32091_, _32090_, _32088_);
  and (_32092_, _32091_, _06282_);
  and (_32093_, _32092_, _32085_);
  and (_32094_, _13359_, \oc8051_golden_model_1.P1 [0]);
  and (_32096_, _14326_, _08603_);
  or (_32097_, _32096_, _32094_);
  and (_32098_, _32097_, _06281_);
  or (_32099_, _32098_, _32093_);
  and (_32100_, _32099_, _07169_);
  and (_32101_, _32080_, _06354_);
  or (_32102_, _32101_, _06345_);
  or (_32103_, _32102_, _32100_);
  or (_32104_, _32087_, _06346_);
  and (_32105_, _32104_, _06278_);
  and (_32107_, _32105_, _32103_);
  and (_32108_, _32076_, _06277_);
  or (_32109_, _32108_, _06270_);
  or (_32110_, _32109_, _32107_);
  or (_32111_, _32083_, _06271_);
  and (_32112_, _32111_, _06267_);
  and (_32113_, _32112_, _32110_);
  and (_32114_, _14358_, _08603_);
  or (_32115_, _32114_, _32094_);
  and (_32116_, _32115_, _06266_);
  or (_32118_, _32116_, _06259_);
  or (_32119_, _32118_, _32113_);
  and (_32120_, _32119_, _32081_);
  or (_32121_, _32120_, _09486_);
  and (_32122_, _09384_, _07961_);
  or (_32123_, _32076_, _06258_);
  or (_32124_, _32123_, _32122_);
  and (_32125_, _32124_, _06251_);
  and (_32126_, _32125_, _32121_);
  and (_32127_, _14413_, _07961_);
  or (_32129_, _32127_, _32076_);
  and (_32130_, _32129_, _05972_);
  or (_32131_, _32130_, _32126_);
  or (_32132_, _32131_, _10080_);
  and (_32133_, _14311_, _07961_);
  or (_32134_, _32076_, _09025_);
  or (_32135_, _32134_, _32133_);
  and (_32136_, _07961_, _08929_);
  or (_32137_, _32136_, _32076_);
  or (_32138_, _32137_, _06216_);
  and (_32140_, _32138_, _09030_);
  and (_32141_, _32140_, _32135_);
  and (_32142_, _32141_, _32132_);
  nor (_32143_, _12532_, _13354_);
  or (_32144_, _32143_, _32076_);
  and (_32145_, _32075_, _06524_);
  and (_32146_, _32145_, _32144_);
  or (_32147_, _32146_, _32142_);
  and (_32148_, _32147_, _07219_);
  nand (_32149_, _32137_, _06426_);
  nor (_32151_, _32149_, _32082_);
  or (_32152_, _32151_, _06532_);
  or (_32153_, _32152_, _32148_);
  and (_32154_, _32153_, _32078_);
  or (_32155_, _32154_, _06437_);
  and (_32156_, _14307_, _07961_);
  or (_32157_, _32076_, _07229_);
  or (_32158_, _32157_, _32156_);
  and (_32159_, _32158_, _07231_);
  and (_32160_, _32159_, _32155_);
  and (_32162_, _32144_, _06535_);
  or (_32163_, _32162_, _06559_);
  or (_32164_, _32163_, _32160_);
  or (_32165_, _32083_, _07240_);
  and (_32166_, _32165_, _32164_);
  or (_32167_, _32166_, _05932_);
  or (_32168_, _32076_, _05933_);
  and (_32169_, _32168_, _32167_);
  or (_32170_, _32169_, _06566_);
  or (_32171_, _32083_, _06570_);
  and (_32173_, _32171_, _01320_);
  and (_32174_, _32173_, _32170_);
  or (_43026_, _32174_, _32074_);
  and (_32175_, _13354_, \oc8051_golden_model_1.P1 [1]);
  and (_32176_, _07961_, _09422_);
  or (_32177_, _32176_, _32175_);
  or (_32178_, _32177_, _07169_);
  or (_32179_, _07961_, \oc8051_golden_model_1.P1 [1]);
  and (_32180_, _14520_, _07961_);
  not (_32181_, _32180_);
  and (_32183_, _32181_, _32179_);
  or (_32184_, _32183_, _06286_);
  and (_32185_, _07961_, \oc8051_golden_model_1.ACC [1]);
  or (_32186_, _32185_, _32175_);
  and (_32187_, _32186_, _07143_);
  and (_32188_, _07144_, \oc8051_golden_model_1.P1 [1]);
  or (_32189_, _32188_, _06285_);
  or (_32190_, _32189_, _32187_);
  and (_32191_, _32190_, _06282_);
  and (_32192_, _32191_, _32184_);
  and (_32194_, _13359_, \oc8051_golden_model_1.P1 [1]);
  and (_32195_, _14508_, _08603_);
  or (_32196_, _32195_, _32194_);
  and (_32197_, _32196_, _06281_);
  or (_32198_, _32197_, _06354_);
  or (_32199_, _32198_, _32192_);
  and (_32200_, _32199_, _32178_);
  or (_32201_, _32200_, _06345_);
  or (_32202_, _32186_, _06346_);
  and (_32203_, _32202_, _06278_);
  and (_32205_, _32203_, _32201_);
  and (_32206_, _14511_, _08603_);
  or (_32207_, _32206_, _32194_);
  and (_32208_, _32207_, _06277_);
  or (_32209_, _32208_, _06270_);
  or (_32210_, _32209_, _32205_);
  and (_32211_, _32195_, _14507_);
  or (_32212_, _32194_, _06271_);
  or (_32213_, _32212_, _32211_);
  and (_32214_, _32213_, _06267_);
  and (_32216_, _32214_, _32210_);
  or (_32217_, _32194_, _14551_);
  and (_32218_, _32217_, _06266_);
  and (_32219_, _32218_, _32196_);
  or (_32220_, _32219_, _06259_);
  or (_32221_, _32220_, _32216_);
  or (_32222_, _32177_, _06260_);
  and (_32223_, _32222_, _32221_);
  or (_32224_, _32223_, _09486_);
  and (_32225_, _09339_, _07961_);
  or (_32227_, _32175_, _06258_);
  or (_32228_, _32227_, _32225_);
  and (_32229_, _32228_, _06251_);
  and (_32230_, _32229_, _32224_);
  and (_32231_, _14607_, _07961_);
  or (_32232_, _32231_, _32175_);
  and (_32233_, _32232_, _05972_);
  or (_32234_, _32233_, _32230_);
  and (_32235_, _32234_, _06399_);
  or (_32236_, _14505_, _13354_);
  and (_32238_, _32179_, _06398_);
  and (_32239_, _32238_, _32236_);
  nand (_32240_, _07961_, _07031_);
  and (_32241_, _32240_, _06215_);
  and (_32242_, _32241_, _32179_);
  or (_32243_, _32242_, _06524_);
  or (_32244_, _32243_, _32239_);
  or (_32245_, _32244_, _32235_);
  and (_32246_, _11253_, _07961_);
  or (_32247_, _32246_, _32175_);
  or (_32249_, _32247_, _09030_);
  and (_32250_, _32249_, _07219_);
  and (_32251_, _32250_, _32245_);
  or (_32252_, _14503_, _13354_);
  and (_32253_, _32179_, _06426_);
  and (_32254_, _32253_, _32252_);
  or (_32255_, _32254_, _06532_);
  or (_32256_, _32255_, _32251_);
  and (_32257_, _32185_, _08325_);
  or (_32258_, _32175_, _07217_);
  or (_32260_, _32258_, _32257_);
  and (_32261_, _32260_, _07229_);
  and (_32262_, _32261_, _32256_);
  or (_32263_, _32240_, _08325_);
  and (_32264_, _32179_, _06437_);
  and (_32265_, _32264_, _32263_);
  or (_32266_, _32265_, _06535_);
  or (_32267_, _32266_, _32262_);
  nor (_32268_, _11252_, _13354_);
  or (_32269_, _32268_, _32175_);
  or (_32271_, _32269_, _07231_);
  and (_32272_, _32271_, _32267_);
  or (_32273_, _32272_, _06559_);
  or (_32274_, _32183_, _07240_);
  and (_32275_, _32274_, _05933_);
  and (_32276_, _32275_, _32273_);
  and (_32277_, _32207_, _05932_);
  or (_32278_, _32277_, _06566_);
  or (_32279_, _32278_, _32276_);
  or (_32280_, _32175_, _06570_);
  or (_32282_, _32280_, _32180_);
  and (_32283_, _32282_, _01320_);
  and (_32284_, _32283_, _32279_);
  nor (_32285_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_32286_, _32285_, _00000_);
  or (_43027_, _32286_, _32284_);
  nor (_32287_, \oc8051_golden_model_1.P1 [2], rst);
  nor (_32288_, _32287_, _00000_);
  and (_32289_, _13354_, \oc8051_golden_model_1.P1 [2]);
  and (_32290_, _07961_, _08662_);
  or (_32292_, _32290_, _32289_);
  or (_32293_, _32292_, _06260_);
  or (_32294_, _32292_, _07169_);
  and (_32295_, _14703_, _07961_);
  or (_32296_, _32295_, _32289_);
  or (_32297_, _32296_, _06286_);
  and (_32298_, _07961_, \oc8051_golden_model_1.ACC [2]);
  or (_32299_, _32298_, _32289_);
  and (_32300_, _32299_, _07143_);
  and (_32301_, _07144_, \oc8051_golden_model_1.P1 [2]);
  or (_32303_, _32301_, _06285_);
  or (_32304_, _32303_, _32300_);
  and (_32305_, _32304_, _06282_);
  and (_32306_, _32305_, _32297_);
  and (_32307_, _13359_, \oc8051_golden_model_1.P1 [2]);
  and (_32308_, _14716_, _08603_);
  or (_32309_, _32308_, _32307_);
  and (_32310_, _32309_, _06281_);
  or (_32311_, _32310_, _06354_);
  or (_32312_, _32311_, _32306_);
  and (_32314_, _32312_, _32294_);
  or (_32315_, _32314_, _06345_);
  or (_32316_, _32299_, _06346_);
  and (_32317_, _32316_, _06278_);
  and (_32318_, _32317_, _32315_);
  and (_32319_, _14699_, _08603_);
  or (_32320_, _32319_, _32307_);
  and (_32321_, _32320_, _06277_);
  or (_32322_, _32321_, _06270_);
  or (_32323_, _32322_, _32318_);
  and (_32325_, _32308_, _14731_);
  or (_32326_, _32307_, _06271_);
  or (_32327_, _32326_, _32325_);
  and (_32328_, _32327_, _06267_);
  and (_32329_, _32328_, _32323_);
  and (_32330_, _14749_, _08603_);
  or (_32331_, _32330_, _32307_);
  and (_32332_, _32331_, _06266_);
  or (_32333_, _32332_, _06259_);
  or (_32334_, _32333_, _32329_);
  and (_32336_, _32334_, _32293_);
  or (_32337_, _32336_, _09486_);
  and (_32338_, _09293_, _07961_);
  or (_32339_, _32289_, _06258_);
  or (_32340_, _32339_, _32338_);
  and (_32341_, _32340_, _06251_);
  and (_32342_, _32341_, _32337_);
  and (_32343_, _14804_, _07961_);
  or (_32344_, _32289_, _32343_);
  and (_32345_, _32344_, _05972_);
  or (_32347_, _32345_, _32342_);
  or (_32348_, _32347_, _10080_);
  and (_32349_, _14697_, _07961_);
  or (_32350_, _32289_, _09025_);
  or (_32351_, _32350_, _32349_);
  and (_32352_, _07961_, _08980_);
  or (_32353_, _32352_, _32289_);
  or (_32354_, _32353_, _06216_);
  and (_32355_, _32354_, _09030_);
  and (_32356_, _32355_, _32351_);
  and (_32358_, _32356_, _32348_);
  and (_32359_, _11250_, _07961_);
  or (_32360_, _32359_, _32289_);
  and (_32361_, _32360_, _06524_);
  or (_32362_, _32361_, _32358_);
  and (_32363_, _32362_, _07219_);
  or (_32364_, _32289_, _08424_);
  and (_32365_, _32353_, _06426_);
  and (_32366_, _32365_, _32364_);
  or (_32367_, _32366_, _32363_);
  and (_32369_, _32367_, _07217_);
  and (_32370_, _32299_, _06532_);
  and (_32371_, _32370_, _32364_);
  or (_32372_, _32371_, _06437_);
  or (_32373_, _32372_, _32369_);
  and (_32374_, _14694_, _07961_);
  or (_32375_, _32289_, _07229_);
  or (_32376_, _32375_, _32374_);
  and (_32377_, _32376_, _07231_);
  and (_32378_, _32377_, _32373_);
  nor (_32380_, _11249_, _13354_);
  or (_32381_, _32380_, _32289_);
  and (_32382_, _32381_, _06535_);
  or (_32383_, _32382_, _06559_);
  or (_32384_, _32383_, _32378_);
  or (_32385_, _32296_, _07240_);
  and (_32386_, _32385_, _05933_);
  and (_32387_, _32386_, _32384_);
  and (_32388_, _32320_, _05932_);
  or (_32389_, _32388_, _06566_);
  or (_32391_, _32389_, _32387_);
  and (_32392_, _14873_, _07961_);
  or (_32393_, _32289_, _06570_);
  or (_32394_, _32393_, _32392_);
  and (_32395_, _32394_, _01320_);
  and (_32396_, _32395_, _32391_);
  or (_43028_, _32396_, _32288_);
  and (_32397_, _13354_, \oc8051_golden_model_1.P1 [3]);
  and (_32398_, _07961_, _09421_);
  or (_32399_, _32398_, _32397_);
  or (_32401_, _32399_, _06260_);
  and (_32402_, _14900_, _07961_);
  or (_32403_, _32402_, _32397_);
  or (_32404_, _32403_, _06286_);
  and (_32405_, _07961_, \oc8051_golden_model_1.ACC [3]);
  or (_32406_, _32405_, _32397_);
  and (_32407_, _32406_, _07143_);
  and (_32408_, _07144_, \oc8051_golden_model_1.P1 [3]);
  or (_32409_, _32408_, _06285_);
  or (_32410_, _32409_, _32407_);
  and (_32412_, _32410_, _06282_);
  and (_32413_, _32412_, _32404_);
  and (_32414_, _13359_, \oc8051_golden_model_1.P1 [3]);
  and (_32415_, _14897_, _08603_);
  or (_32416_, _32415_, _32414_);
  and (_32417_, _32416_, _06281_);
  or (_32418_, _32417_, _06354_);
  or (_32419_, _32418_, _32413_);
  or (_32420_, _32399_, _07169_);
  and (_32421_, _32420_, _32419_);
  or (_32423_, _32421_, _06345_);
  or (_32424_, _32406_, _06346_);
  and (_32425_, _32424_, _06278_);
  and (_32426_, _32425_, _32423_);
  and (_32427_, _14895_, _08603_);
  or (_32428_, _32427_, _32414_);
  and (_32429_, _32428_, _06277_);
  or (_32430_, _32429_, _06270_);
  or (_32431_, _32430_, _32426_);
  or (_32432_, _32414_, _14926_);
  and (_32434_, _32432_, _32416_);
  or (_32435_, _32434_, _06271_);
  and (_32436_, _32435_, _06267_);
  and (_32437_, _32436_, _32431_);
  and (_32438_, _14943_, _08603_);
  or (_32439_, _32438_, _32414_);
  and (_32440_, _32439_, _06266_);
  or (_32441_, _32440_, _06259_);
  or (_32442_, _32441_, _32437_);
  and (_32443_, _32442_, _32401_);
  or (_32445_, _32443_, _09486_);
  and (_32446_, _09247_, _07961_);
  or (_32447_, _32397_, _06258_);
  or (_32448_, _32447_, _32446_);
  and (_32449_, _32448_, _06251_);
  and (_32450_, _32449_, _32445_);
  and (_32451_, _14998_, _07961_);
  or (_32452_, _32397_, _32451_);
  and (_32453_, _32452_, _05972_);
  or (_32454_, _32453_, _32450_);
  or (_32456_, _32454_, _10080_);
  and (_32457_, _14893_, _07961_);
  or (_32458_, _32397_, _09025_);
  or (_32459_, _32458_, _32457_);
  and (_32460_, _07961_, _08809_);
  or (_32461_, _32460_, _32397_);
  or (_32462_, _32461_, _06216_);
  and (_32463_, _32462_, _09030_);
  and (_32464_, _32463_, _32459_);
  and (_32465_, _32464_, _32456_);
  and (_32467_, _12529_, _07961_);
  or (_32468_, _32467_, _32397_);
  and (_32469_, _32468_, _06524_);
  or (_32470_, _32469_, _32465_);
  and (_32471_, _32470_, _07219_);
  or (_32472_, _32397_, _08280_);
  and (_32473_, _32461_, _06426_);
  and (_32474_, _32473_, _32472_);
  or (_32475_, _32474_, _32471_);
  and (_32476_, _32475_, _07217_);
  and (_32478_, _32406_, _06532_);
  and (_32479_, _32478_, _32472_);
  or (_32480_, _32479_, _06437_);
  or (_32481_, _32480_, _32476_);
  and (_32482_, _14890_, _07961_);
  or (_32483_, _32397_, _07229_);
  or (_32484_, _32483_, _32482_);
  and (_32485_, _32484_, _07231_);
  and (_32486_, _32485_, _32481_);
  nor (_32487_, _11247_, _13354_);
  or (_32489_, _32487_, _32397_);
  and (_32490_, _32489_, _06535_);
  or (_32491_, _32490_, _06559_);
  or (_32492_, _32491_, _32486_);
  or (_32493_, _32403_, _07240_);
  and (_32494_, _32493_, _05933_);
  and (_32495_, _32494_, _32492_);
  and (_32496_, _32428_, _05932_);
  or (_32497_, _32496_, _06566_);
  or (_32498_, _32497_, _32495_);
  and (_32500_, _15068_, _07961_);
  or (_32501_, _32397_, _06570_);
  or (_32502_, _32501_, _32500_);
  and (_32503_, _32502_, _01320_);
  and (_32504_, _32503_, _32498_);
  nor (_32505_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_32506_, _32505_, _00000_);
  or (_43029_, _32506_, _32504_);
  nor (_32507_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_32508_, _32507_, _00000_);
  and (_32510_, _13354_, \oc8051_golden_model_1.P1 [4]);
  and (_32511_, _09420_, _07961_);
  or (_32512_, _32511_, _32510_);
  or (_32513_, _32512_, _06260_);
  and (_32514_, _13359_, \oc8051_golden_model_1.P1 [4]);
  and (_32515_, _15145_, _08603_);
  or (_32516_, _32515_, _32514_);
  and (_32517_, _32516_, _06277_);
  and (_32518_, _15133_, _07961_);
  or (_32519_, _32518_, _32510_);
  or (_32521_, _32519_, _06286_);
  and (_32522_, _07961_, \oc8051_golden_model_1.ACC [4]);
  or (_32523_, _32522_, _32510_);
  and (_32524_, _32523_, _07143_);
  and (_32525_, _07144_, \oc8051_golden_model_1.P1 [4]);
  or (_32526_, _32525_, _06285_);
  or (_32527_, _32526_, _32524_);
  and (_32528_, _32527_, _06282_);
  and (_32529_, _32528_, _32521_);
  and (_32530_, _15116_, _08603_);
  or (_32532_, _32530_, _32514_);
  and (_32533_, _32532_, _06281_);
  or (_32534_, _32533_, _06354_);
  or (_32535_, _32534_, _32529_);
  or (_32536_, _32512_, _07169_);
  and (_32537_, _32536_, _32535_);
  or (_32538_, _32537_, _06345_);
  or (_32539_, _32523_, _06346_);
  and (_32540_, _32539_, _06278_);
  and (_32541_, _32540_, _32538_);
  or (_32543_, _32541_, _32517_);
  and (_32544_, _32543_, _06271_);
  or (_32545_, _32514_, _15152_);
  and (_32546_, _32532_, _06270_);
  and (_32547_, _32546_, _32545_);
  or (_32548_, _32547_, _32544_);
  and (_32549_, _32548_, _06267_);
  and (_32550_, _15170_, _08603_);
  or (_32551_, _32550_, _32514_);
  and (_32552_, _32551_, _06266_);
  or (_32554_, _32552_, _06259_);
  or (_32555_, _32554_, _32549_);
  and (_32556_, _32555_, _32513_);
  or (_32557_, _32556_, _09486_);
  and (_32558_, _09437_, _07961_);
  or (_32559_, _32510_, _06258_);
  or (_32560_, _32559_, _32558_);
  and (_32561_, _32560_, _06251_);
  and (_32562_, _32561_, _32557_);
  and (_32563_, _15226_, _07961_);
  or (_32565_, _32563_, _32510_);
  and (_32566_, _32565_, _05972_);
  or (_32567_, _32566_, _10080_);
  or (_32568_, _32567_, _32562_);
  and (_32569_, _15114_, _07961_);
  or (_32570_, _32510_, _09025_);
  or (_32571_, _32570_, _32569_);
  and (_32572_, _08919_, _07961_);
  or (_32573_, _32572_, _32510_);
  or (_32574_, _32573_, _06216_);
  and (_32576_, _32574_, _09030_);
  and (_32577_, _32576_, _32571_);
  and (_32578_, _32577_, _32568_);
  and (_32579_, _11245_, _07961_);
  or (_32580_, _32579_, _32510_);
  and (_32581_, _32580_, _06524_);
  or (_32582_, _32581_, _32578_);
  and (_32583_, _32582_, _07219_);
  or (_32584_, _32510_, _08528_);
  and (_32585_, _32573_, _06426_);
  and (_32587_, _32585_, _32584_);
  or (_32588_, _32587_, _32583_);
  and (_32589_, _32588_, _07217_);
  and (_32590_, _32523_, _06532_);
  and (_32591_, _32590_, _32584_);
  or (_32592_, _32591_, _06437_);
  or (_32593_, _32592_, _32589_);
  and (_32594_, _15111_, _07961_);
  or (_32595_, _32510_, _07229_);
  or (_32596_, _32595_, _32594_);
  and (_32597_, _32596_, _07231_);
  and (_32598_, _32597_, _32593_);
  nor (_32599_, _11244_, _13354_);
  or (_32600_, _32599_, _32510_);
  and (_32601_, _32600_, _06535_);
  or (_32602_, _32601_, _06559_);
  or (_32603_, _32602_, _32598_);
  or (_32604_, _32519_, _07240_);
  and (_32605_, _32604_, _05933_);
  and (_32606_, _32605_, _32603_);
  and (_32608_, _32516_, _05932_);
  or (_32609_, _32608_, _06566_);
  or (_32610_, _32609_, _32606_);
  and (_32611_, _15296_, _07961_);
  or (_32612_, _32510_, _06570_);
  or (_32613_, _32612_, _32611_);
  and (_32614_, _32613_, _01320_);
  and (_32615_, _32614_, _32610_);
  or (_43030_, _32615_, _32508_);
  and (_32616_, _13354_, \oc8051_golden_model_1.P1 [5]);
  and (_32618_, _15330_, _07961_);
  or (_32619_, _32618_, _32616_);
  or (_32620_, _32619_, _06286_);
  and (_32621_, _07961_, \oc8051_golden_model_1.ACC [5]);
  or (_32622_, _32621_, _32616_);
  and (_32623_, _32622_, _07143_);
  and (_32624_, _07144_, \oc8051_golden_model_1.P1 [5]);
  or (_32625_, _32624_, _06285_);
  or (_32626_, _32625_, _32623_);
  and (_32627_, _32626_, _06282_);
  and (_32629_, _32627_, _32620_);
  and (_32630_, _13359_, \oc8051_golden_model_1.P1 [5]);
  and (_32631_, _15315_, _08603_);
  or (_32632_, _32631_, _32630_);
  and (_32633_, _32632_, _06281_);
  or (_32634_, _32633_, _06354_);
  or (_32635_, _32634_, _32629_);
  and (_32636_, _09419_, _07961_);
  or (_32637_, _32636_, _32616_);
  or (_32638_, _32637_, _07169_);
  and (_32640_, _32638_, _32635_);
  or (_32641_, _32640_, _06345_);
  or (_32642_, _32622_, _06346_);
  and (_32643_, _32642_, _06278_);
  and (_32644_, _32643_, _32641_);
  and (_32645_, _15342_, _08603_);
  or (_32646_, _32645_, _32630_);
  and (_32647_, _32646_, _06277_);
  or (_32648_, _32647_, _06270_);
  or (_32649_, _32648_, _32644_);
  or (_32651_, _32630_, _15349_);
  and (_32652_, _32651_, _32632_);
  or (_32653_, _32652_, _06271_);
  and (_32654_, _32653_, _06267_);
  and (_32655_, _32654_, _32649_);
  or (_32656_, _32630_, _15365_);
  and (_32657_, _32656_, _06266_);
  and (_32658_, _32657_, _32632_);
  or (_32659_, _32658_, _06259_);
  or (_32660_, _32659_, _32655_);
  or (_32662_, _32637_, _06260_);
  and (_32663_, _32662_, _32660_);
  or (_32664_, _32663_, _09486_);
  and (_32665_, _09436_, _07961_);
  or (_32666_, _32616_, _06258_);
  or (_32667_, _32666_, _32665_);
  and (_32668_, _32667_, _06251_);
  and (_32669_, _32668_, _32664_);
  and (_32670_, _15421_, _07961_);
  or (_32671_, _32670_, _32616_);
  and (_32673_, _32671_, _05972_);
  or (_32674_, _32673_, _10080_);
  or (_32675_, _32674_, _32669_);
  and (_32676_, _15313_, _07961_);
  or (_32677_, _32616_, _09025_);
  or (_32678_, _32677_, _32676_);
  and (_32679_, _08913_, _07961_);
  or (_32680_, _32679_, _32616_);
  or (_32681_, _32680_, _06216_);
  and (_32682_, _32681_, _09030_);
  and (_32684_, _32682_, _32678_);
  and (_32685_, _32684_, _32675_);
  and (_32686_, _12536_, _07961_);
  or (_32687_, _32686_, _32616_);
  and (_32688_, _32687_, _06524_);
  or (_32689_, _32688_, _32685_);
  and (_32690_, _32689_, _07219_);
  or (_32691_, _32616_, _08231_);
  and (_32692_, _32680_, _06426_);
  and (_32693_, _32692_, _32691_);
  or (_32695_, _32693_, _32690_);
  and (_32696_, _32695_, _07217_);
  and (_32697_, _32622_, _06532_);
  and (_32698_, _32697_, _32691_);
  or (_32699_, _32698_, _06437_);
  or (_32700_, _32699_, _32696_);
  and (_32701_, _15310_, _07961_);
  or (_32702_, _32616_, _07229_);
  or (_32703_, _32702_, _32701_);
  and (_32704_, _32703_, _07231_);
  and (_32706_, _32704_, _32700_);
  nor (_32707_, _11241_, _13354_);
  or (_32708_, _32707_, _32616_);
  and (_32709_, _32708_, _06535_);
  or (_32710_, _32709_, _06559_);
  or (_32711_, _32710_, _32706_);
  or (_32712_, _32619_, _07240_);
  and (_32713_, _32712_, _05933_);
  and (_32714_, _32713_, _32711_);
  and (_32715_, _32646_, _05932_);
  or (_32717_, _32715_, _06566_);
  or (_32718_, _32717_, _32714_);
  and (_32719_, _15493_, _07961_);
  or (_32720_, _32616_, _06570_);
  or (_32721_, _32720_, _32719_);
  and (_32722_, _32721_, _01320_);
  and (_32723_, _32722_, _32718_);
  nor (_32724_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_32725_, _32724_, _00000_);
  or (_43031_, _32725_, _32723_);
  and (_32727_, _13354_, \oc8051_golden_model_1.P1 [6]);
  and (_32728_, _15521_, _07961_);
  or (_32729_, _32728_, _32727_);
  or (_32730_, _32729_, _06286_);
  and (_32731_, _07961_, \oc8051_golden_model_1.ACC [6]);
  or (_32732_, _32731_, _32727_);
  and (_32733_, _32732_, _07143_);
  and (_32734_, _07144_, \oc8051_golden_model_1.P1 [6]);
  or (_32735_, _32734_, _06285_);
  or (_32736_, _32735_, _32733_);
  and (_32738_, _32736_, _06282_);
  and (_32739_, _32738_, _32730_);
  and (_32740_, _13359_, \oc8051_golden_model_1.P1 [6]);
  and (_32741_, _15535_, _08603_);
  or (_32742_, _32741_, _32740_);
  and (_32743_, _32742_, _06281_);
  or (_32744_, _32743_, _06354_);
  or (_32745_, _32744_, _32739_);
  and (_32746_, _09418_, _07961_);
  or (_32747_, _32746_, _32727_);
  or (_32749_, _32747_, _07169_);
  and (_32750_, _32749_, _32745_);
  or (_32751_, _32750_, _06345_);
  or (_32752_, _32732_, _06346_);
  and (_32753_, _32752_, _06278_);
  and (_32754_, _32753_, _32751_);
  and (_32755_, _15544_, _08603_);
  or (_32756_, _32755_, _32740_);
  and (_32757_, _32756_, _06277_);
  or (_32758_, _32757_, _06270_);
  or (_32760_, _32758_, _32754_);
  or (_32761_, _32740_, _15551_);
  and (_32762_, _32761_, _32742_);
  or (_32763_, _32762_, _06271_);
  and (_32764_, _32763_, _06267_);
  and (_32765_, _32764_, _32760_);
  and (_32766_, _15568_, _08603_);
  or (_32767_, _32766_, _32740_);
  and (_32768_, _32767_, _06266_);
  or (_32769_, _32768_, _06259_);
  or (_32771_, _32769_, _32765_);
  or (_32772_, _32747_, _06260_);
  and (_32773_, _32772_, _32771_);
  or (_32774_, _32773_, _09486_);
  and (_32775_, _09435_, _07961_);
  or (_32776_, _32727_, _06258_);
  or (_32777_, _32776_, _32775_);
  and (_32778_, _32777_, _06251_);
  and (_32779_, _32778_, _32774_);
  and (_32780_, _15623_, _07961_);
  or (_32782_, _32780_, _32727_);
  and (_32783_, _32782_, _05972_);
  or (_32784_, _32783_, _10080_);
  or (_32785_, _32784_, _32779_);
  and (_32786_, _15517_, _07961_);
  or (_32787_, _32727_, _09025_);
  or (_32788_, _32787_, _32786_);
  and (_32789_, _08845_, _07961_);
  or (_32790_, _32789_, _32727_);
  or (_32791_, _32790_, _06216_);
  and (_32793_, _32791_, _09030_);
  and (_32794_, _32793_, _32788_);
  and (_32795_, _32794_, _32785_);
  and (_32796_, _11239_, _07961_);
  or (_32797_, _32796_, _32727_);
  and (_32798_, _32797_, _06524_);
  or (_32799_, _32798_, _32795_);
  and (_32800_, _32799_, _07219_);
  or (_32801_, _32727_, _08128_);
  and (_32802_, _32790_, _06426_);
  and (_32804_, _32802_, _32801_);
  or (_32805_, _32804_, _32800_);
  and (_32806_, _32805_, _07217_);
  and (_32807_, _32732_, _06532_);
  and (_32808_, _32807_, _32801_);
  or (_32809_, _32808_, _06437_);
  or (_32810_, _32809_, _32806_);
  and (_32811_, _15514_, _07961_);
  or (_32812_, _32727_, _07229_);
  or (_32813_, _32812_, _32811_);
  and (_32815_, _32813_, _07231_);
  and (_32816_, _32815_, _32810_);
  nor (_32817_, _11238_, _13354_);
  or (_32818_, _32817_, _32727_);
  and (_32819_, _32818_, _06535_);
  or (_32820_, _32819_, _06559_);
  or (_32821_, _32820_, _32816_);
  or (_32822_, _32729_, _07240_);
  and (_32823_, _32822_, _05933_);
  and (_32824_, _32823_, _32821_);
  and (_32826_, _32756_, _05932_);
  or (_32827_, _32826_, _06566_);
  or (_32828_, _32827_, _32824_);
  and (_32829_, _15695_, _07961_);
  or (_32830_, _32727_, _06570_);
  or (_32831_, _32830_, _32829_);
  and (_32832_, _32831_, _01320_);
  and (_32833_, _32832_, _32828_);
  nor (_32834_, \oc8051_golden_model_1.P1 [6], rst);
  nor (_32835_, _32834_, _00000_);
  or (_43032_, _32835_, _32833_);
  and (_32837_, _01324_, \oc8051_golden_model_1.IP [0]);
  and (_32838_, _07937_, \oc8051_golden_model_1.ACC [0]);
  and (_32839_, _32838_, _08374_);
  and (_32840_, _13455_, \oc8051_golden_model_1.IP [0]);
  or (_32841_, _32840_, _07217_);
  or (_32842_, _32841_, _32839_);
  and (_32843_, _07937_, _07135_);
  or (_32844_, _32843_, _32840_);
  or (_32845_, _32844_, _06260_);
  nor (_32847_, _08374_, _13455_);
  or (_32848_, _32847_, _32840_);
  and (_32849_, _32848_, _06285_);
  and (_32850_, _07144_, \oc8051_golden_model_1.IP [0]);
  or (_32851_, _32838_, _32840_);
  and (_32852_, _32851_, _07143_);
  or (_32853_, _32852_, _32850_);
  and (_32854_, _32853_, _06286_);
  or (_32855_, _32854_, _06281_);
  or (_32856_, _32855_, _32849_);
  and (_32858_, _14326_, _08589_);
  and (_32859_, _13460_, \oc8051_golden_model_1.IP [0]);
  or (_32860_, _32859_, _06282_);
  or (_32861_, _32860_, _32858_);
  and (_32862_, _32861_, _07169_);
  and (_32863_, _32862_, _32856_);
  and (_32864_, _32844_, _06354_);
  or (_32865_, _32864_, _06345_);
  or (_32866_, _32865_, _32863_);
  or (_32867_, _32851_, _06346_);
  and (_32869_, _32867_, _06278_);
  and (_32870_, _32869_, _32866_);
  and (_32871_, _32840_, _06277_);
  or (_32872_, _32871_, _06270_);
  or (_32873_, _32872_, _32870_);
  or (_32874_, _32848_, _06271_);
  and (_32875_, _32874_, _06267_);
  and (_32876_, _32875_, _32873_);
  and (_32877_, _14358_, _08589_);
  or (_32878_, _32877_, _32859_);
  and (_32880_, _32878_, _06266_);
  or (_32881_, _32880_, _06259_);
  or (_32882_, _32881_, _32876_);
  and (_32883_, _32882_, _32845_);
  or (_32884_, _32883_, _09486_);
  and (_32885_, _09384_, _07937_);
  or (_32886_, _32840_, _06258_);
  or (_32887_, _32886_, _32885_);
  and (_32888_, _32887_, _06251_);
  and (_32889_, _32888_, _32884_);
  and (_32891_, _14413_, _07937_);
  or (_32892_, _32891_, _32840_);
  and (_32893_, _32892_, _05972_);
  or (_32894_, _32893_, _32889_);
  or (_32895_, _32894_, _10080_);
  and (_32896_, _14311_, _07937_);
  or (_32897_, _32840_, _09025_);
  or (_32898_, _32897_, _32896_);
  and (_32899_, _07937_, _08929_);
  or (_32900_, _32899_, _32840_);
  or (_32902_, _32900_, _06216_);
  and (_32903_, _32902_, _09030_);
  and (_32904_, _32903_, _32898_);
  and (_32905_, _32904_, _32895_);
  nor (_32906_, _12532_, _13455_);
  or (_32907_, _32906_, _32840_);
  nor (_32908_, _32839_, _09030_);
  and (_32909_, _32908_, _32907_);
  or (_32910_, _32909_, _32905_);
  and (_32911_, _32910_, _07219_);
  nand (_32913_, _32900_, _06426_);
  nor (_32914_, _32913_, _32847_);
  or (_32915_, _32914_, _06532_);
  or (_32916_, _32915_, _32911_);
  and (_32917_, _32916_, _32842_);
  or (_32918_, _32917_, _06437_);
  and (_32919_, _14307_, _07937_);
  or (_32920_, _32919_, _32840_);
  or (_32921_, _32920_, _07229_);
  and (_32922_, _32921_, _07231_);
  and (_32924_, _32922_, _32918_);
  and (_32925_, _32907_, _06535_);
  or (_32926_, _32925_, _06559_);
  or (_32927_, _32926_, _32924_);
  or (_32928_, _32848_, _07240_);
  and (_32929_, _32928_, _32927_);
  or (_32930_, _32929_, _05932_);
  or (_32931_, _32840_, _05933_);
  and (_32932_, _32931_, _32930_);
  or (_32933_, _32932_, _06566_);
  or (_32935_, _32848_, _06570_);
  and (_32936_, _32935_, _01320_);
  and (_32937_, _32936_, _32933_);
  or (_32938_, _32937_, _32837_);
  and (_43034_, _32938_, _42355_);
  not (_32939_, \oc8051_golden_model_1.IP [1]);
  nor (_32940_, _01320_, _32939_);
  nor (_32941_, _07937_, _32939_);
  and (_32942_, _07937_, _09422_);
  or (_32943_, _32942_, _32941_);
  or (_32945_, _32943_, _07169_);
  or (_32946_, _07937_, \oc8051_golden_model_1.IP [1]);
  and (_32947_, _14520_, _07937_);
  not (_32948_, _32947_);
  and (_32949_, _32948_, _32946_);
  or (_32950_, _32949_, _06286_);
  and (_32951_, _07937_, \oc8051_golden_model_1.ACC [1]);
  or (_32952_, _32951_, _32941_);
  and (_32953_, _32952_, _07143_);
  nor (_32954_, _07143_, _32939_);
  or (_32956_, _32954_, _06285_);
  or (_32957_, _32956_, _32953_);
  and (_32958_, _32957_, _06282_);
  and (_32959_, _32958_, _32950_);
  nor (_32960_, _08589_, _32939_);
  and (_32961_, _14508_, _08589_);
  or (_32962_, _32961_, _32960_);
  and (_32963_, _32962_, _06281_);
  or (_32964_, _32963_, _06354_);
  or (_32965_, _32964_, _32959_);
  and (_32967_, _32965_, _32945_);
  or (_32968_, _32967_, _06345_);
  or (_32969_, _32952_, _06346_);
  and (_32970_, _32969_, _06278_);
  and (_32971_, _32970_, _32968_);
  and (_32972_, _14511_, _08589_);
  or (_32973_, _32972_, _32960_);
  and (_32974_, _32973_, _06277_);
  or (_32975_, _32974_, _06270_);
  or (_32976_, _32975_, _32971_);
  and (_32978_, _32961_, _14507_);
  or (_32979_, _32960_, _06271_);
  or (_32980_, _32979_, _32978_);
  and (_32981_, _32980_, _06267_);
  and (_32982_, _32981_, _32976_);
  or (_32983_, _32960_, _14551_);
  and (_32984_, _32983_, _06266_);
  and (_32985_, _32984_, _32962_);
  or (_32986_, _32985_, _06259_);
  or (_32987_, _32986_, _32982_);
  or (_32989_, _32943_, _06260_);
  and (_32990_, _32989_, _32987_);
  or (_32991_, _32990_, _09486_);
  and (_32992_, _09339_, _07937_);
  or (_32993_, _32941_, _06258_);
  or (_32994_, _32993_, _32992_);
  and (_32995_, _32994_, _06251_);
  and (_32996_, _32995_, _32991_);
  and (_32997_, _14607_, _07937_);
  or (_32998_, _32997_, _32941_);
  and (_33000_, _32998_, _05972_);
  or (_33001_, _33000_, _32996_);
  and (_33002_, _33001_, _06399_);
  or (_33003_, _14505_, _13455_);
  and (_33004_, _32946_, _06398_);
  and (_33005_, _33004_, _33003_);
  nand (_33006_, _07937_, _07031_);
  and (_33007_, _33006_, _06215_);
  and (_33008_, _33007_, _32946_);
  or (_33009_, _33008_, _06524_);
  or (_33011_, _33009_, _33005_);
  or (_33012_, _33011_, _33002_);
  nor (_33013_, _11252_, _13455_);
  or (_33014_, _33013_, _32941_);
  nand (_33015_, _11251_, _07937_);
  and (_33016_, _33015_, _33014_);
  or (_33017_, _33016_, _09030_);
  and (_33018_, _33017_, _07219_);
  and (_33019_, _33018_, _33012_);
  or (_33020_, _14503_, _13455_);
  and (_33022_, _32946_, _06426_);
  and (_33023_, _33022_, _33020_);
  or (_33024_, _33023_, _06532_);
  or (_33025_, _33024_, _33019_);
  nor (_33026_, _32941_, _07217_);
  nand (_33027_, _33026_, _33015_);
  and (_33028_, _33027_, _07229_);
  and (_33029_, _33028_, _33025_);
  or (_33030_, _33006_, _08325_);
  and (_33031_, _32946_, _06437_);
  and (_33033_, _33031_, _33030_);
  or (_33034_, _33033_, _06535_);
  or (_33035_, _33034_, _33029_);
  or (_33036_, _33014_, _07231_);
  and (_33037_, _33036_, _33035_);
  or (_33038_, _33037_, _06559_);
  or (_33039_, _32949_, _07240_);
  and (_33040_, _33039_, _05933_);
  and (_33041_, _33040_, _33038_);
  and (_33042_, _32973_, _05932_);
  or (_33044_, _33042_, _06566_);
  or (_33045_, _33044_, _33041_);
  or (_33046_, _32941_, _06570_);
  or (_33047_, _33046_, _32947_);
  and (_33048_, _33047_, _01320_);
  and (_33049_, _33048_, _33045_);
  or (_33050_, _33049_, _32940_);
  and (_43035_, _33050_, _42355_);
  and (_33051_, _01324_, \oc8051_golden_model_1.IP [2]);
  and (_33052_, _13455_, \oc8051_golden_model_1.IP [2]);
  and (_33054_, _07937_, _08662_);
  or (_33055_, _33054_, _33052_);
  or (_33056_, _33055_, _06260_);
  or (_33057_, _33055_, _07169_);
  and (_33058_, _14703_, _07937_);
  or (_33059_, _33058_, _33052_);
  or (_33060_, _33059_, _06286_);
  and (_33061_, _07937_, \oc8051_golden_model_1.ACC [2]);
  or (_33062_, _33061_, _33052_);
  and (_33063_, _33062_, _07143_);
  and (_33065_, _07144_, \oc8051_golden_model_1.IP [2]);
  or (_33066_, _33065_, _06285_);
  or (_33067_, _33066_, _33063_);
  and (_33068_, _33067_, _06282_);
  and (_33069_, _33068_, _33060_);
  and (_33070_, _13460_, \oc8051_golden_model_1.IP [2]);
  and (_33071_, _14716_, _08589_);
  or (_33072_, _33071_, _33070_);
  and (_33073_, _33072_, _06281_);
  or (_33074_, _33073_, _06354_);
  or (_33076_, _33074_, _33069_);
  and (_33077_, _33076_, _33057_);
  or (_33078_, _33077_, _06345_);
  or (_33079_, _33062_, _06346_);
  and (_33080_, _33079_, _06278_);
  and (_33081_, _33080_, _33078_);
  and (_33082_, _14699_, _08589_);
  or (_33083_, _33082_, _33070_);
  and (_33084_, _33083_, _06277_);
  or (_33085_, _33084_, _06270_);
  or (_33087_, _33085_, _33081_);
  and (_33088_, _33071_, _14731_);
  or (_33089_, _33070_, _06271_);
  or (_33090_, _33089_, _33088_);
  and (_33091_, _33090_, _06267_);
  and (_33092_, _33091_, _33087_);
  and (_33093_, _14749_, _08589_);
  or (_33094_, _33093_, _33070_);
  and (_33095_, _33094_, _06266_);
  or (_33096_, _33095_, _06259_);
  or (_33098_, _33096_, _33092_);
  and (_33099_, _33098_, _33056_);
  or (_33100_, _33099_, _09486_);
  and (_33101_, _09293_, _07937_);
  or (_33102_, _33052_, _06258_);
  or (_33103_, _33102_, _33101_);
  and (_33104_, _33103_, _06251_);
  and (_33105_, _33104_, _33100_);
  and (_33106_, _14804_, _07937_);
  or (_33107_, _33052_, _33106_);
  and (_33109_, _33107_, _05972_);
  or (_33110_, _33109_, _33105_);
  or (_33111_, _33110_, _10080_);
  and (_33112_, _14697_, _07937_);
  or (_33113_, _33052_, _09025_);
  or (_33114_, _33113_, _33112_);
  and (_33115_, _07937_, _08980_);
  or (_33116_, _33115_, _33052_);
  or (_33117_, _33116_, _06216_);
  and (_33118_, _33117_, _09030_);
  and (_33120_, _33118_, _33114_);
  and (_33121_, _33120_, _33111_);
  and (_33122_, _11250_, _07937_);
  or (_33123_, _33122_, _33052_);
  and (_33124_, _33123_, _06524_);
  or (_33125_, _33124_, _33121_);
  and (_33126_, _33125_, _07219_);
  or (_33127_, _33052_, _08424_);
  and (_33128_, _33116_, _06426_);
  and (_33129_, _33128_, _33127_);
  or (_33131_, _33129_, _33126_);
  and (_33132_, _33131_, _07217_);
  and (_33133_, _33062_, _06532_);
  and (_33134_, _33133_, _33127_);
  or (_33135_, _33134_, _06437_);
  or (_33136_, _33135_, _33132_);
  and (_33137_, _14694_, _07937_);
  or (_33138_, _33052_, _07229_);
  or (_33139_, _33138_, _33137_);
  and (_33140_, _33139_, _07231_);
  and (_33142_, _33140_, _33136_);
  nor (_33143_, _11249_, _13455_);
  or (_33144_, _33143_, _33052_);
  and (_33145_, _33144_, _06535_);
  or (_33146_, _33145_, _06559_);
  or (_33147_, _33146_, _33142_);
  or (_33148_, _33059_, _07240_);
  and (_33149_, _33148_, _05933_);
  and (_33150_, _33149_, _33147_);
  and (_33151_, _33083_, _05932_);
  or (_33153_, _33151_, _06566_);
  or (_33154_, _33153_, _33150_);
  and (_33155_, _14873_, _07937_);
  or (_33156_, _33052_, _06570_);
  or (_33157_, _33156_, _33155_);
  and (_33158_, _33157_, _01320_);
  and (_33159_, _33158_, _33154_);
  or (_33160_, _33159_, _33051_);
  and (_43036_, _33160_, _42355_);
  and (_33161_, _01324_, \oc8051_golden_model_1.IP [3]);
  and (_33163_, _13455_, \oc8051_golden_model_1.IP [3]);
  and (_33164_, _07937_, _09421_);
  or (_33165_, _33164_, _33163_);
  or (_33166_, _33165_, _06260_);
  and (_33167_, _14900_, _07937_);
  or (_33168_, _33167_, _33163_);
  or (_33169_, _33168_, _06286_);
  and (_33170_, _07937_, \oc8051_golden_model_1.ACC [3]);
  or (_33171_, _33170_, _33163_);
  and (_33172_, _33171_, _07143_);
  and (_33174_, _07144_, \oc8051_golden_model_1.IP [3]);
  or (_33175_, _33174_, _06285_);
  or (_33176_, _33175_, _33172_);
  and (_33177_, _33176_, _06282_);
  and (_33178_, _33177_, _33169_);
  and (_33179_, _13460_, \oc8051_golden_model_1.IP [3]);
  and (_33180_, _14897_, _08589_);
  or (_33181_, _33180_, _33179_);
  and (_33182_, _33181_, _06281_);
  or (_33183_, _33182_, _06354_);
  or (_33185_, _33183_, _33178_);
  or (_33186_, _33165_, _07169_);
  and (_33187_, _33186_, _33185_);
  or (_33188_, _33187_, _06345_);
  or (_33189_, _33171_, _06346_);
  and (_33190_, _33189_, _06278_);
  and (_33191_, _33190_, _33188_);
  and (_33192_, _14895_, _08589_);
  or (_33193_, _33192_, _33179_);
  and (_33194_, _33193_, _06277_);
  or (_33196_, _33194_, _06270_);
  or (_33197_, _33196_, _33191_);
  or (_33198_, _33179_, _14926_);
  and (_33199_, _33198_, _33181_);
  or (_33200_, _33199_, _06271_);
  and (_33201_, _33200_, _06267_);
  and (_33202_, _33201_, _33197_);
  and (_33203_, _14943_, _08589_);
  or (_33204_, _33203_, _33179_);
  and (_33205_, _33204_, _06266_);
  or (_33207_, _33205_, _06259_);
  or (_33208_, _33207_, _33202_);
  and (_33209_, _33208_, _33166_);
  or (_33210_, _33209_, _09486_);
  and (_33211_, _09247_, _07937_);
  or (_33212_, _33163_, _06258_);
  or (_33213_, _33212_, _33211_);
  and (_33214_, _33213_, _06251_);
  and (_33215_, _33214_, _33210_);
  and (_33216_, _14998_, _07937_);
  or (_33218_, _33163_, _33216_);
  and (_33219_, _33218_, _05972_);
  or (_33220_, _33219_, _33215_);
  or (_33221_, _33220_, _10080_);
  and (_33222_, _14893_, _07937_);
  or (_33223_, _33163_, _09025_);
  or (_33224_, _33223_, _33222_);
  and (_33225_, _07937_, _08809_);
  or (_33226_, _33225_, _33163_);
  or (_33227_, _33226_, _06216_);
  and (_33229_, _33227_, _09030_);
  and (_33230_, _33229_, _33224_);
  and (_33231_, _33230_, _33221_);
  and (_33232_, _12529_, _07937_);
  or (_33233_, _33232_, _33163_);
  and (_33234_, _33233_, _06524_);
  or (_33235_, _33234_, _33231_);
  and (_33236_, _33235_, _07219_);
  or (_33237_, _33163_, _08280_);
  and (_33238_, _33226_, _06426_);
  and (_33240_, _33238_, _33237_);
  or (_33241_, _33240_, _33236_);
  and (_33242_, _33241_, _07217_);
  and (_33243_, _33171_, _06532_);
  and (_33244_, _33243_, _33237_);
  or (_33245_, _33244_, _06437_);
  or (_33246_, _33245_, _33242_);
  and (_33247_, _14890_, _07937_);
  or (_33248_, _33163_, _07229_);
  or (_33249_, _33248_, _33247_);
  and (_33251_, _33249_, _07231_);
  and (_33252_, _33251_, _33246_);
  nor (_33253_, _11247_, _13455_);
  or (_33254_, _33253_, _33163_);
  and (_33255_, _33254_, _06535_);
  or (_33256_, _33255_, _06559_);
  or (_33257_, _33256_, _33252_);
  or (_33258_, _33168_, _07240_);
  and (_33259_, _33258_, _05933_);
  and (_33260_, _33259_, _33257_);
  and (_33262_, _33193_, _05932_);
  or (_33263_, _33262_, _06566_);
  or (_33264_, _33263_, _33260_);
  and (_33265_, _15068_, _07937_);
  or (_33266_, _33163_, _06570_);
  or (_33267_, _33266_, _33265_);
  and (_33268_, _33267_, _01320_);
  and (_33269_, _33268_, _33264_);
  or (_33270_, _33269_, _33161_);
  and (_43037_, _33270_, _42355_);
  and (_33272_, _01324_, \oc8051_golden_model_1.IP [4]);
  and (_33273_, _13455_, \oc8051_golden_model_1.IP [4]);
  and (_33274_, _09420_, _07937_);
  or (_33275_, _33274_, _33273_);
  or (_33276_, _33275_, _06260_);
  and (_33277_, _13460_, \oc8051_golden_model_1.IP [4]);
  and (_33278_, _15145_, _08589_);
  or (_33279_, _33278_, _33277_);
  and (_33280_, _33279_, _06277_);
  and (_33281_, _15133_, _07937_);
  or (_33283_, _33281_, _33273_);
  or (_33284_, _33283_, _06286_);
  and (_33285_, _07937_, \oc8051_golden_model_1.ACC [4]);
  or (_33286_, _33285_, _33273_);
  and (_33287_, _33286_, _07143_);
  and (_33288_, _07144_, \oc8051_golden_model_1.IP [4]);
  or (_33289_, _33288_, _06285_);
  or (_33290_, _33289_, _33287_);
  and (_33291_, _33290_, _06282_);
  and (_33292_, _33291_, _33284_);
  and (_33294_, _15116_, _08589_);
  or (_33295_, _33294_, _33277_);
  and (_33296_, _33295_, _06281_);
  or (_33297_, _33296_, _06354_);
  or (_33298_, _33297_, _33292_);
  or (_33299_, _33275_, _07169_);
  and (_33300_, _33299_, _33298_);
  or (_33301_, _33300_, _06345_);
  or (_33302_, _33286_, _06346_);
  and (_33303_, _33302_, _06278_);
  and (_33305_, _33303_, _33301_);
  or (_33306_, _33305_, _33280_);
  and (_33307_, _33306_, _06271_);
  or (_33308_, _33277_, _15152_);
  and (_33309_, _33308_, _06270_);
  and (_33310_, _33309_, _33295_);
  or (_33311_, _33310_, _33307_);
  and (_33312_, _33311_, _06267_);
  and (_33313_, _15170_, _08589_);
  or (_33314_, _33313_, _33277_);
  and (_33315_, _33314_, _06266_);
  or (_33316_, _33315_, _06259_);
  or (_33317_, _33316_, _33312_);
  and (_33318_, _33317_, _33276_);
  or (_33319_, _33318_, _09486_);
  and (_33320_, _09437_, _07937_);
  or (_33321_, _33273_, _06258_);
  or (_33322_, _33321_, _33320_);
  and (_33323_, _33322_, _06251_);
  and (_33324_, _33323_, _33319_);
  and (_33326_, _15226_, _07937_);
  or (_33327_, _33326_, _33273_);
  and (_33328_, _33327_, _05972_);
  or (_33329_, _33328_, _10080_);
  or (_33330_, _33329_, _33324_);
  and (_33331_, _15114_, _07937_);
  or (_33332_, _33273_, _09025_);
  or (_33333_, _33332_, _33331_);
  and (_33334_, _08919_, _07937_);
  or (_33335_, _33334_, _33273_);
  or (_33337_, _33335_, _06216_);
  and (_33338_, _33337_, _09030_);
  and (_33339_, _33338_, _33333_);
  and (_33340_, _33339_, _33330_);
  and (_33341_, _11245_, _07937_);
  or (_33342_, _33341_, _33273_);
  and (_33343_, _33342_, _06524_);
  or (_33344_, _33343_, _33340_);
  and (_33345_, _33344_, _07219_);
  or (_33346_, _33273_, _08528_);
  and (_33348_, _33335_, _06426_);
  and (_33349_, _33348_, _33346_);
  or (_33350_, _33349_, _33345_);
  and (_33351_, _33350_, _07217_);
  and (_33352_, _33286_, _06532_);
  and (_33353_, _33352_, _33346_);
  or (_33354_, _33353_, _06437_);
  or (_33355_, _33354_, _33351_);
  and (_33356_, _15111_, _07937_);
  or (_33357_, _33273_, _07229_);
  or (_33359_, _33357_, _33356_);
  and (_33360_, _33359_, _07231_);
  and (_33361_, _33360_, _33355_);
  nor (_33362_, _11244_, _13455_);
  or (_33363_, _33362_, _33273_);
  and (_33364_, _33363_, _06535_);
  or (_33365_, _33364_, _06559_);
  or (_33366_, _33365_, _33361_);
  or (_33367_, _33283_, _07240_);
  and (_33368_, _33367_, _05933_);
  and (_33370_, _33368_, _33366_);
  and (_33371_, _33279_, _05932_);
  or (_33372_, _33371_, _06566_);
  or (_33373_, _33372_, _33370_);
  and (_33374_, _15296_, _07937_);
  or (_33375_, _33273_, _06570_);
  or (_33376_, _33375_, _33374_);
  and (_33377_, _33376_, _01320_);
  and (_33378_, _33377_, _33373_);
  or (_33379_, _33378_, _33272_);
  and (_43038_, _33379_, _42355_);
  and (_33381_, _01324_, \oc8051_golden_model_1.IP [5]);
  and (_33382_, _13455_, \oc8051_golden_model_1.IP [5]);
  and (_33383_, _15330_, _07937_);
  or (_33384_, _33383_, _33382_);
  or (_33385_, _33384_, _06286_);
  and (_33386_, _07937_, \oc8051_golden_model_1.ACC [5]);
  or (_33387_, _33386_, _33382_);
  and (_33388_, _33387_, _07143_);
  and (_33389_, _07144_, \oc8051_golden_model_1.IP [5]);
  or (_33391_, _33389_, _06285_);
  or (_33392_, _33391_, _33388_);
  and (_33393_, _33392_, _06282_);
  and (_33394_, _33393_, _33385_);
  and (_33395_, _13460_, \oc8051_golden_model_1.IP [5]);
  and (_33396_, _15315_, _08589_);
  or (_33397_, _33396_, _33395_);
  and (_33398_, _33397_, _06281_);
  or (_33399_, _33398_, _06354_);
  or (_33400_, _33399_, _33394_);
  and (_33402_, _09419_, _07937_);
  or (_33403_, _33402_, _33382_);
  or (_33404_, _33403_, _07169_);
  and (_33405_, _33404_, _33400_);
  or (_33406_, _33405_, _06345_);
  or (_33407_, _33387_, _06346_);
  and (_33408_, _33407_, _06278_);
  and (_33409_, _33408_, _33406_);
  and (_33410_, _15342_, _08589_);
  or (_33411_, _33410_, _33395_);
  and (_33413_, _33411_, _06277_);
  or (_33414_, _33413_, _06270_);
  or (_33415_, _33414_, _33409_);
  or (_33416_, _33395_, _15349_);
  and (_33417_, _33416_, _33397_);
  or (_33418_, _33417_, _06271_);
  and (_33419_, _33418_, _06267_);
  and (_33420_, _33419_, _33415_);
  or (_33421_, _33395_, _15365_);
  and (_33422_, _33421_, _06266_);
  and (_33424_, _33422_, _33397_);
  or (_33425_, _33424_, _06259_);
  or (_33426_, _33425_, _33420_);
  or (_33427_, _33403_, _06260_);
  and (_33428_, _33427_, _33426_);
  or (_33429_, _33428_, _09486_);
  and (_33430_, _09436_, _07937_);
  or (_33431_, _33382_, _06258_);
  or (_33432_, _33431_, _33430_);
  and (_33433_, _33432_, _06251_);
  and (_33435_, _33433_, _33429_);
  and (_33436_, _15421_, _07937_);
  or (_33437_, _33436_, _33382_);
  and (_33438_, _33437_, _05972_);
  or (_33439_, _33438_, _10080_);
  or (_33440_, _33439_, _33435_);
  and (_33441_, _15313_, _07937_);
  or (_33442_, _33382_, _09025_);
  or (_33443_, _33442_, _33441_);
  and (_33444_, _08913_, _07937_);
  or (_33446_, _33444_, _33382_);
  or (_33447_, _33446_, _06216_);
  and (_33448_, _33447_, _09030_);
  and (_33449_, _33448_, _33443_);
  and (_33450_, _33449_, _33440_);
  and (_33451_, _12536_, _07937_);
  or (_33452_, _33451_, _33382_);
  and (_33453_, _33452_, _06524_);
  or (_33454_, _33453_, _33450_);
  and (_33455_, _33454_, _07219_);
  or (_33457_, _33382_, _08231_);
  and (_33458_, _33446_, _06426_);
  and (_33459_, _33458_, _33457_);
  or (_33460_, _33459_, _33455_);
  and (_33461_, _33460_, _07217_);
  and (_33462_, _33387_, _06532_);
  and (_33463_, _33462_, _33457_);
  or (_33464_, _33463_, _06437_);
  or (_33465_, _33464_, _33461_);
  and (_33466_, _15310_, _07937_);
  or (_33468_, _33382_, _07229_);
  or (_33469_, _33468_, _33466_);
  and (_33470_, _33469_, _07231_);
  and (_33471_, _33470_, _33465_);
  nor (_33472_, _11241_, _13455_);
  or (_33473_, _33472_, _33382_);
  and (_33474_, _33473_, _06535_);
  or (_33475_, _33474_, _06559_);
  or (_33476_, _33475_, _33471_);
  or (_33477_, _33384_, _07240_);
  and (_33479_, _33477_, _05933_);
  and (_33480_, _33479_, _33476_);
  and (_33481_, _33411_, _05932_);
  or (_33482_, _33481_, _06566_);
  or (_33483_, _33482_, _33480_);
  and (_33484_, _15493_, _07937_);
  or (_33485_, _33382_, _06570_);
  or (_33486_, _33485_, _33484_);
  and (_33487_, _33486_, _01320_);
  and (_33488_, _33487_, _33483_);
  or (_33490_, _33488_, _33381_);
  and (_43040_, _33490_, _42355_);
  and (_33491_, _01324_, \oc8051_golden_model_1.IP [6]);
  and (_33492_, _13455_, \oc8051_golden_model_1.IP [6]);
  and (_33493_, _15521_, _07937_);
  or (_33494_, _33493_, _33492_);
  or (_33495_, _33494_, _06286_);
  and (_33496_, _07937_, \oc8051_golden_model_1.ACC [6]);
  or (_33497_, _33496_, _33492_);
  and (_33498_, _33497_, _07143_);
  and (_33500_, _07144_, \oc8051_golden_model_1.IP [6]);
  or (_33501_, _33500_, _06285_);
  or (_33502_, _33501_, _33498_);
  and (_33503_, _33502_, _06282_);
  and (_33504_, _33503_, _33495_);
  and (_33505_, _13460_, \oc8051_golden_model_1.IP [6]);
  and (_33506_, _15535_, _08589_);
  or (_33507_, _33506_, _33505_);
  and (_33508_, _33507_, _06281_);
  or (_33509_, _33508_, _06354_);
  or (_33511_, _33509_, _33504_);
  and (_33512_, _09418_, _07937_);
  or (_33513_, _33512_, _33492_);
  or (_33514_, _33513_, _07169_);
  and (_33515_, _33514_, _33511_);
  or (_33516_, _33515_, _06345_);
  or (_33517_, _33497_, _06346_);
  and (_33518_, _33517_, _06278_);
  and (_33519_, _33518_, _33516_);
  and (_33520_, _15544_, _08589_);
  or (_33522_, _33520_, _33505_);
  and (_33523_, _33522_, _06277_);
  or (_33524_, _33523_, _06270_);
  or (_33525_, _33524_, _33519_);
  or (_33526_, _33505_, _15551_);
  and (_33527_, _33526_, _33507_);
  or (_33528_, _33527_, _06271_);
  and (_33529_, _33528_, _06267_);
  and (_33530_, _33529_, _33525_);
  and (_33531_, _15568_, _08589_);
  or (_33533_, _33531_, _33505_);
  and (_33534_, _33533_, _06266_);
  or (_33535_, _33534_, _06259_);
  or (_33536_, _33535_, _33530_);
  or (_33537_, _33513_, _06260_);
  and (_33538_, _33537_, _33536_);
  or (_33539_, _33538_, _09486_);
  and (_33540_, _09435_, _07937_);
  or (_33541_, _33492_, _06258_);
  or (_33542_, _33541_, _33540_);
  and (_33544_, _33542_, _06251_);
  and (_33545_, _33544_, _33539_);
  and (_33546_, _15623_, _07937_);
  or (_33547_, _33546_, _33492_);
  and (_33548_, _33547_, _05972_);
  or (_33549_, _33548_, _10080_);
  or (_33550_, _33549_, _33545_);
  and (_33551_, _15517_, _07937_);
  or (_33552_, _33492_, _09025_);
  or (_33553_, _33552_, _33551_);
  and (_33555_, _08845_, _07937_);
  or (_33556_, _33555_, _33492_);
  or (_33557_, _33556_, _06216_);
  and (_33558_, _33557_, _09030_);
  and (_33559_, _33558_, _33553_);
  and (_33560_, _33559_, _33550_);
  and (_33561_, _11239_, _07937_);
  or (_33562_, _33561_, _33492_);
  and (_33563_, _33562_, _06524_);
  or (_33564_, _33563_, _33560_);
  and (_33566_, _33564_, _07219_);
  or (_33567_, _33492_, _08128_);
  and (_33568_, _33556_, _06426_);
  and (_33569_, _33568_, _33567_);
  or (_33570_, _33569_, _33566_);
  and (_33571_, _33570_, _07217_);
  and (_33572_, _33497_, _06532_);
  and (_33573_, _33572_, _33567_);
  or (_33574_, _33573_, _06437_);
  or (_33575_, _33574_, _33571_);
  and (_33577_, _15514_, _07937_);
  or (_33578_, _33492_, _07229_);
  or (_33579_, _33578_, _33577_);
  and (_33580_, _33579_, _07231_);
  and (_33581_, _33580_, _33575_);
  nor (_33582_, _11238_, _13455_);
  or (_33583_, _33582_, _33492_);
  and (_33584_, _33583_, _06535_);
  or (_33585_, _33584_, _06559_);
  or (_33586_, _33585_, _33581_);
  or (_33588_, _33494_, _07240_);
  and (_33589_, _33588_, _05933_);
  and (_33590_, _33589_, _33586_);
  and (_33591_, _33522_, _05932_);
  or (_33592_, _33591_, _06566_);
  or (_33593_, _33592_, _33590_);
  and (_33594_, _15695_, _07937_);
  or (_33595_, _33492_, _06570_);
  or (_33596_, _33595_, _33594_);
  and (_33597_, _33596_, _01320_);
  and (_33599_, _33597_, _33593_);
  or (_33600_, _33599_, _33491_);
  and (_43041_, _33600_, _42355_);
  and (_33601_, _01324_, \oc8051_golden_model_1.IE [0]);
  and (_33602_, _07881_, \oc8051_golden_model_1.ACC [0]);
  and (_33603_, _33602_, _08374_);
  and (_33604_, _13557_, \oc8051_golden_model_1.IE [0]);
  or (_33605_, _33604_, _07217_);
  or (_33606_, _33605_, _33603_);
  and (_33607_, _07881_, _07135_);
  or (_33609_, _33607_, _33604_);
  or (_33610_, _33609_, _06260_);
  nor (_33611_, _08374_, _13557_);
  or (_33612_, _33611_, _33604_);
  or (_33613_, _33612_, _06286_);
  or (_33614_, _33602_, _33604_);
  and (_33615_, _33614_, _07143_);
  and (_33616_, _07144_, \oc8051_golden_model_1.IE [0]);
  or (_33617_, _33616_, _06285_);
  or (_33618_, _33617_, _33615_);
  and (_33620_, _33618_, _06282_);
  and (_33621_, _33620_, _33613_);
  and (_33622_, _13562_, \oc8051_golden_model_1.IE [0]);
  and (_33623_, _14326_, _08609_);
  or (_33624_, _33623_, _33622_);
  and (_33625_, _33624_, _06281_);
  or (_33626_, _33625_, _33621_);
  and (_33627_, _33626_, _07169_);
  and (_33628_, _33609_, _06354_);
  or (_33629_, _33628_, _06345_);
  or (_33631_, _33629_, _33627_);
  or (_33632_, _33614_, _06346_);
  and (_33633_, _33632_, _06278_);
  and (_33634_, _33633_, _33631_);
  and (_33635_, _33604_, _06277_);
  or (_33636_, _33635_, _06270_);
  or (_33637_, _33636_, _33634_);
  or (_33638_, _33612_, _06271_);
  and (_33639_, _33638_, _06267_);
  and (_33640_, _33639_, _33637_);
  and (_33642_, _14358_, _08609_);
  or (_33643_, _33642_, _33622_);
  and (_33644_, _33643_, _06266_);
  or (_33645_, _33644_, _06259_);
  or (_33646_, _33645_, _33640_);
  and (_33647_, _33646_, _33610_);
  or (_33648_, _33647_, _09486_);
  and (_33649_, _09384_, _07881_);
  or (_33650_, _33604_, _06258_);
  or (_33651_, _33650_, _33649_);
  and (_33653_, _33651_, _06251_);
  and (_33654_, _33653_, _33648_);
  and (_33655_, _14413_, _07881_);
  or (_33656_, _33655_, _33604_);
  and (_33657_, _33656_, _05972_);
  or (_33658_, _33657_, _33654_);
  or (_33659_, _33658_, _10080_);
  and (_33660_, _14311_, _07881_);
  or (_33661_, _33604_, _09025_);
  or (_33662_, _33661_, _33660_);
  and (_33664_, _07881_, _08929_);
  or (_33665_, _33664_, _33604_);
  or (_33666_, _33665_, _06216_);
  and (_33667_, _33666_, _09030_);
  and (_33668_, _33667_, _33662_);
  and (_33669_, _33668_, _33659_);
  nor (_33670_, _12532_, _13557_);
  or (_33671_, _33670_, _33604_);
  nor (_33672_, _33603_, _09030_);
  and (_33673_, _33672_, _33671_);
  or (_33675_, _33673_, _33669_);
  and (_33676_, _33675_, _07219_);
  nand (_33677_, _33665_, _06426_);
  nor (_33678_, _33677_, _33611_);
  or (_33679_, _33678_, _06532_);
  or (_33680_, _33679_, _33676_);
  and (_33681_, _33680_, _33606_);
  or (_33682_, _33681_, _06437_);
  and (_33683_, _14307_, _07881_);
  or (_33684_, _33604_, _07229_);
  or (_33686_, _33684_, _33683_);
  and (_33687_, _33686_, _07231_);
  and (_33688_, _33687_, _33682_);
  and (_33689_, _33671_, _06535_);
  or (_33690_, _33689_, _06559_);
  or (_33691_, _33690_, _33688_);
  or (_33692_, _33612_, _07240_);
  and (_33693_, _33692_, _33691_);
  or (_33694_, _33693_, _05932_);
  or (_33695_, _33604_, _05933_);
  and (_33697_, _33695_, _33694_);
  or (_33698_, _33697_, _06566_);
  or (_33699_, _33612_, _06570_);
  and (_33700_, _33699_, _01320_);
  and (_33701_, _33700_, _33698_);
  or (_33702_, _33701_, _33601_);
  and (_43042_, _33702_, _42355_);
  not (_33703_, \oc8051_golden_model_1.IE [1]);
  nor (_33704_, _01320_, _33703_);
  nor (_33705_, _07881_, _33703_);
  and (_33707_, _07881_, _09422_);
  or (_33708_, _33707_, _33705_);
  and (_33709_, _33708_, _06354_);
  nor (_33710_, _08609_, _33703_);
  and (_33711_, _14508_, _08609_);
  or (_33712_, _33711_, _33710_);
  or (_33713_, _33712_, _06282_);
  or (_33714_, _07881_, \oc8051_golden_model_1.IE [1]);
  and (_33715_, _14520_, _07881_);
  not (_33716_, _33715_);
  and (_33718_, _33716_, _33714_);
  and (_33719_, _33718_, _06285_);
  nor (_33720_, _07143_, _33703_);
  and (_33721_, _07881_, \oc8051_golden_model_1.ACC [1]);
  or (_33722_, _33721_, _33705_);
  and (_33723_, _33722_, _07143_);
  or (_33724_, _33723_, _33720_);
  and (_33725_, _33724_, _06286_);
  or (_33726_, _33725_, _06281_);
  or (_33727_, _33726_, _33719_);
  and (_33729_, _33727_, _33713_);
  and (_33730_, _33729_, _07169_);
  or (_33731_, _33730_, _33709_);
  or (_33732_, _33731_, _06345_);
  or (_33733_, _33722_, _06346_);
  and (_33734_, _33733_, _06278_);
  and (_33735_, _33734_, _33732_);
  and (_33736_, _14511_, _08609_);
  or (_33737_, _33736_, _33710_);
  and (_33738_, _33737_, _06277_);
  or (_33740_, _33738_, _06270_);
  or (_33741_, _33740_, _33735_);
  or (_33742_, _33710_, _14507_);
  and (_33743_, _33742_, _33712_);
  or (_33744_, _33743_, _06271_);
  and (_33745_, _33744_, _06267_);
  and (_33746_, _33745_, _33741_);
  or (_33747_, _33710_, _14551_);
  and (_33748_, _33747_, _06266_);
  and (_33749_, _33748_, _33712_);
  or (_33751_, _33749_, _06259_);
  or (_33752_, _33751_, _33746_);
  or (_33753_, _33708_, _06260_);
  and (_33754_, _33753_, _33752_);
  or (_33755_, _33754_, _09486_);
  and (_33756_, _09339_, _07881_);
  or (_33757_, _33705_, _06258_);
  or (_33758_, _33757_, _33756_);
  and (_33759_, _33758_, _06251_);
  and (_33760_, _33759_, _33755_);
  and (_33762_, _14607_, _07881_);
  or (_33763_, _33762_, _33705_);
  and (_33764_, _33763_, _05972_);
  or (_33765_, _33764_, _33760_);
  and (_33766_, _33765_, _06399_);
  or (_33767_, _14505_, _13557_);
  and (_33768_, _33714_, _06398_);
  and (_33769_, _33768_, _33767_);
  nand (_33770_, _07881_, _07031_);
  and (_33771_, _33770_, _06215_);
  and (_33773_, _33771_, _33714_);
  or (_33774_, _33773_, _06524_);
  or (_33775_, _33774_, _33769_);
  or (_33776_, _33775_, _33766_);
  nor (_33777_, _11252_, _13557_);
  or (_33778_, _33777_, _33705_);
  nand (_33779_, _11251_, _07881_);
  and (_33780_, _33779_, _33778_);
  or (_33781_, _33780_, _09030_);
  and (_33782_, _33781_, _07219_);
  and (_33784_, _33782_, _33776_);
  or (_33785_, _14503_, _13557_);
  and (_33786_, _33714_, _06426_);
  and (_33787_, _33786_, _33785_);
  or (_33788_, _33787_, _06532_);
  or (_33789_, _33788_, _33784_);
  nor (_33790_, _33705_, _07217_);
  nand (_33791_, _33790_, _33779_);
  and (_33792_, _33791_, _07229_);
  and (_33793_, _33792_, _33789_);
  or (_33795_, _33770_, _08325_);
  and (_33796_, _33714_, _06437_);
  and (_33797_, _33796_, _33795_);
  or (_33798_, _33797_, _06535_);
  or (_33799_, _33798_, _33793_);
  or (_33800_, _33778_, _07231_);
  and (_33801_, _33800_, _33799_);
  or (_33802_, _33801_, _06559_);
  or (_33803_, _33718_, _07240_);
  and (_33804_, _33803_, _05933_);
  and (_33806_, _33804_, _33802_);
  and (_33807_, _33737_, _05932_);
  or (_33808_, _33807_, _06566_);
  or (_33809_, _33808_, _33806_);
  or (_33810_, _33705_, _06570_);
  or (_33811_, _33810_, _33715_);
  and (_33812_, _33811_, _01320_);
  and (_33813_, _33812_, _33809_);
  or (_33814_, _33813_, _33704_);
  and (_43044_, _33814_, _42355_);
  and (_33816_, _01324_, \oc8051_golden_model_1.IE [2]);
  and (_33817_, _13557_, \oc8051_golden_model_1.IE [2]);
  and (_33818_, _07881_, _08662_);
  or (_33819_, _33818_, _33817_);
  or (_33820_, _33819_, _06260_);
  and (_33821_, _33819_, _06354_);
  and (_33822_, _13562_, \oc8051_golden_model_1.IE [2]);
  and (_33823_, _14716_, _08609_);
  or (_33824_, _33823_, _33822_);
  or (_33825_, _33824_, _06282_);
  and (_33827_, _14703_, _07881_);
  or (_33828_, _33827_, _33817_);
  and (_33829_, _33828_, _06285_);
  and (_33830_, _07144_, \oc8051_golden_model_1.IE [2]);
  and (_33831_, _07881_, \oc8051_golden_model_1.ACC [2]);
  or (_33832_, _33831_, _33817_);
  and (_33833_, _33832_, _07143_);
  or (_33834_, _33833_, _33830_);
  and (_33835_, _33834_, _06286_);
  or (_33836_, _33835_, _06281_);
  or (_33838_, _33836_, _33829_);
  and (_33839_, _33838_, _33825_);
  and (_33840_, _33839_, _07169_);
  or (_33841_, _33840_, _33821_);
  or (_33842_, _33841_, _06345_);
  or (_33843_, _33832_, _06346_);
  and (_33844_, _33843_, _06278_);
  and (_33845_, _33844_, _33842_);
  and (_33846_, _14699_, _08609_);
  or (_33847_, _33846_, _33822_);
  and (_33849_, _33847_, _06277_);
  or (_33850_, _33849_, _06270_);
  or (_33851_, _33850_, _33845_);
  or (_33852_, _33822_, _14731_);
  and (_33853_, _33852_, _33824_);
  or (_33854_, _33853_, _06271_);
  and (_33855_, _33854_, _06267_);
  and (_33856_, _33855_, _33851_);
  and (_33857_, _14749_, _08609_);
  or (_33858_, _33857_, _33822_);
  and (_33860_, _33858_, _06266_);
  or (_33861_, _33860_, _06259_);
  or (_33862_, _33861_, _33856_);
  and (_33863_, _33862_, _33820_);
  or (_33864_, _33863_, _09486_);
  and (_33865_, _09293_, _07881_);
  or (_33866_, _33817_, _06258_);
  or (_33867_, _33866_, _33865_);
  and (_33868_, _33867_, _06251_);
  and (_33869_, _33868_, _33864_);
  and (_33871_, _14804_, _07881_);
  or (_33872_, _33817_, _33871_);
  and (_33873_, _33872_, _05972_);
  or (_33874_, _33873_, _33869_);
  or (_33875_, _33874_, _10080_);
  and (_33876_, _14697_, _07881_);
  or (_33877_, _33817_, _09025_);
  or (_33878_, _33877_, _33876_);
  and (_33879_, _07881_, _08980_);
  or (_33880_, _33879_, _33817_);
  or (_33882_, _33880_, _06216_);
  and (_33883_, _33882_, _09030_);
  and (_33884_, _33883_, _33878_);
  and (_33885_, _33884_, _33875_);
  and (_33886_, _11250_, _07881_);
  or (_33887_, _33886_, _33817_);
  and (_33888_, _33887_, _06524_);
  or (_33889_, _33888_, _33885_);
  and (_33890_, _33889_, _07219_);
  or (_33891_, _33817_, _08424_);
  and (_33893_, _33880_, _06426_);
  and (_33894_, _33893_, _33891_);
  or (_33895_, _33894_, _33890_);
  and (_33896_, _33895_, _07217_);
  and (_33897_, _33832_, _06532_);
  and (_33898_, _33897_, _33891_);
  or (_33899_, _33898_, _06437_);
  or (_33900_, _33899_, _33896_);
  and (_33901_, _14694_, _07881_);
  or (_33902_, _33817_, _07229_);
  or (_33904_, _33902_, _33901_);
  and (_33905_, _33904_, _07231_);
  and (_33906_, _33905_, _33900_);
  nor (_33907_, _11249_, _13557_);
  or (_33908_, _33907_, _33817_);
  and (_33909_, _33908_, _06535_);
  or (_33910_, _33909_, _06559_);
  or (_33911_, _33910_, _33906_);
  or (_33912_, _33828_, _07240_);
  and (_33913_, _33912_, _05933_);
  and (_33915_, _33913_, _33911_);
  and (_33916_, _33847_, _05932_);
  or (_33917_, _33916_, _06566_);
  or (_33918_, _33917_, _33915_);
  and (_33919_, _14873_, _07881_);
  or (_33920_, _33817_, _06570_);
  or (_33921_, _33920_, _33919_);
  and (_33922_, _33921_, _01320_);
  and (_33923_, _33922_, _33918_);
  or (_33924_, _33923_, _33816_);
  and (_43045_, _33924_, _42355_);
  and (_33926_, _01324_, \oc8051_golden_model_1.IE [3]);
  and (_33927_, _13557_, \oc8051_golden_model_1.IE [3]);
  and (_33928_, _07881_, _09421_);
  or (_33929_, _33928_, _33927_);
  or (_33930_, _33929_, _06260_);
  and (_33931_, _14900_, _07881_);
  or (_33932_, _33931_, _33927_);
  or (_33933_, _33932_, _06286_);
  and (_33934_, _07881_, \oc8051_golden_model_1.ACC [3]);
  or (_33936_, _33934_, _33927_);
  and (_33937_, _33936_, _07143_);
  and (_33938_, _07144_, \oc8051_golden_model_1.IE [3]);
  or (_33939_, _33938_, _06285_);
  or (_33940_, _33939_, _33937_);
  and (_33941_, _33940_, _06282_);
  and (_33942_, _33941_, _33933_);
  and (_33943_, _13562_, \oc8051_golden_model_1.IE [3]);
  and (_33944_, _14897_, _08609_);
  or (_33945_, _33944_, _33943_);
  and (_33947_, _33945_, _06281_);
  or (_33948_, _33947_, _06354_);
  or (_33949_, _33948_, _33942_);
  or (_33950_, _33929_, _07169_);
  and (_33951_, _33950_, _33949_);
  or (_33952_, _33951_, _06345_);
  or (_33953_, _33936_, _06346_);
  and (_33954_, _33953_, _06278_);
  and (_33955_, _33954_, _33952_);
  and (_33956_, _14895_, _08609_);
  or (_33958_, _33956_, _33943_);
  and (_33959_, _33958_, _06277_);
  or (_33960_, _33959_, _06270_);
  or (_33961_, _33960_, _33955_);
  or (_33962_, _33943_, _14926_);
  and (_33963_, _33962_, _33945_);
  or (_33964_, _33963_, _06271_);
  and (_33965_, _33964_, _06267_);
  and (_33966_, _33965_, _33961_);
  and (_33967_, _14943_, _08609_);
  or (_33969_, _33967_, _33943_);
  and (_33970_, _33969_, _06266_);
  or (_33971_, _33970_, _06259_);
  or (_33972_, _33971_, _33966_);
  and (_33973_, _33972_, _33930_);
  or (_33974_, _33973_, _09486_);
  and (_33975_, _09247_, _07881_);
  or (_33976_, _33927_, _06258_);
  or (_33977_, _33976_, _33975_);
  and (_33978_, _33977_, _06251_);
  and (_33980_, _33978_, _33974_);
  and (_33981_, _14998_, _07881_);
  or (_33982_, _33927_, _33981_);
  and (_33983_, _33982_, _05972_);
  or (_33984_, _33983_, _33980_);
  or (_33985_, _33984_, _10080_);
  and (_33986_, _14893_, _07881_);
  or (_33987_, _33927_, _09025_);
  or (_33988_, _33987_, _33986_);
  and (_33989_, _07881_, _08809_);
  or (_33991_, _33989_, _33927_);
  or (_33992_, _33991_, _06216_);
  and (_33993_, _33992_, _09030_);
  and (_33994_, _33993_, _33988_);
  and (_33995_, _33994_, _33985_);
  and (_33996_, _12529_, _07881_);
  or (_33997_, _33996_, _33927_);
  and (_33998_, _33997_, _06524_);
  or (_33999_, _33998_, _33995_);
  and (_34000_, _33999_, _07219_);
  or (_34002_, _33927_, _08280_);
  and (_34003_, _33991_, _06426_);
  and (_34004_, _34003_, _34002_);
  or (_34005_, _34004_, _34000_);
  and (_34006_, _34005_, _07217_);
  and (_34007_, _33936_, _06532_);
  and (_34008_, _34007_, _34002_);
  or (_34009_, _34008_, _06437_);
  or (_34010_, _34009_, _34006_);
  and (_34011_, _14890_, _07881_);
  or (_34013_, _33927_, _07229_);
  or (_34014_, _34013_, _34011_);
  and (_34015_, _34014_, _07231_);
  and (_34016_, _34015_, _34010_);
  nor (_34017_, _11247_, _13557_);
  or (_34018_, _34017_, _33927_);
  and (_34019_, _34018_, _06535_);
  or (_34020_, _34019_, _06559_);
  or (_34021_, _34020_, _34016_);
  or (_34022_, _33932_, _07240_);
  and (_34024_, _34022_, _05933_);
  and (_34025_, _34024_, _34021_);
  and (_34026_, _33958_, _05932_);
  or (_34027_, _34026_, _06566_);
  or (_34028_, _34027_, _34025_);
  and (_34029_, _15068_, _07881_);
  or (_34030_, _33927_, _06570_);
  or (_34031_, _34030_, _34029_);
  and (_34032_, _34031_, _01320_);
  and (_34033_, _34032_, _34028_);
  or (_34035_, _34033_, _33926_);
  and (_43046_, _34035_, _42355_);
  and (_34036_, _01324_, \oc8051_golden_model_1.IE [4]);
  and (_34037_, _13557_, \oc8051_golden_model_1.IE [4]);
  and (_34038_, _09420_, _07881_);
  or (_34039_, _34038_, _34037_);
  or (_34040_, _34039_, _06260_);
  and (_34041_, _13562_, \oc8051_golden_model_1.IE [4]);
  and (_34042_, _15145_, _08609_);
  or (_34043_, _34042_, _34041_);
  and (_34045_, _34043_, _06277_);
  and (_34046_, _15133_, _07881_);
  or (_34047_, _34046_, _34037_);
  or (_34048_, _34047_, _06286_);
  and (_34049_, _07881_, \oc8051_golden_model_1.ACC [4]);
  or (_34050_, _34049_, _34037_);
  and (_34051_, _34050_, _07143_);
  and (_34052_, _07144_, \oc8051_golden_model_1.IE [4]);
  or (_34053_, _34052_, _06285_);
  or (_34054_, _34053_, _34051_);
  and (_34056_, _34054_, _06282_);
  and (_34057_, _34056_, _34048_);
  and (_34058_, _15116_, _08609_);
  or (_34059_, _34058_, _34041_);
  and (_34060_, _34059_, _06281_);
  or (_34061_, _34060_, _06354_);
  or (_34062_, _34061_, _34057_);
  or (_34063_, _34039_, _07169_);
  and (_34064_, _34063_, _34062_);
  or (_34065_, _34064_, _06345_);
  or (_34067_, _34050_, _06346_);
  and (_34068_, _34067_, _06278_);
  and (_34069_, _34068_, _34065_);
  or (_34070_, _34069_, _34045_);
  and (_34071_, _34070_, _06271_);
  or (_34072_, _34041_, _15152_);
  and (_34073_, _34059_, _06270_);
  and (_34074_, _34073_, _34072_);
  or (_34075_, _34074_, _34071_);
  and (_34076_, _34075_, _06267_);
  and (_34078_, _15170_, _08609_);
  or (_34079_, _34078_, _34041_);
  and (_34080_, _34079_, _06266_);
  or (_34081_, _34080_, _06259_);
  or (_34082_, _34081_, _34076_);
  and (_34083_, _34082_, _34040_);
  or (_34084_, _34083_, _09486_);
  and (_34085_, _09437_, _07881_);
  or (_34086_, _34037_, _06258_);
  or (_34087_, _34086_, _34085_);
  and (_34089_, _34087_, _06251_);
  and (_34090_, _34089_, _34084_);
  and (_34091_, _15226_, _07881_);
  or (_34092_, _34091_, _34037_);
  and (_34093_, _34092_, _05972_);
  or (_34094_, _34093_, _10080_);
  or (_34095_, _34094_, _34090_);
  and (_34096_, _15114_, _07881_);
  or (_34097_, _34037_, _09025_);
  or (_34098_, _34097_, _34096_);
  and (_34099_, _08919_, _07881_);
  or (_34100_, _34099_, _34037_);
  or (_34101_, _34100_, _06216_);
  and (_34102_, _34101_, _09030_);
  and (_34103_, _34102_, _34098_);
  and (_34104_, _34103_, _34095_);
  and (_34105_, _11245_, _07881_);
  or (_34106_, _34105_, _34037_);
  and (_34107_, _34106_, _06524_);
  or (_34108_, _34107_, _34104_);
  and (_34110_, _34108_, _07219_);
  or (_34111_, _34037_, _08528_);
  and (_34112_, _34100_, _06426_);
  and (_34113_, _34112_, _34111_);
  or (_34114_, _34113_, _34110_);
  and (_34115_, _34114_, _07217_);
  and (_34116_, _34050_, _06532_);
  and (_34117_, _34116_, _34111_);
  or (_34118_, _34117_, _06437_);
  or (_34119_, _34118_, _34115_);
  and (_34121_, _15111_, _07881_);
  or (_34122_, _34037_, _07229_);
  or (_34123_, _34122_, _34121_);
  and (_34124_, _34123_, _07231_);
  and (_34125_, _34124_, _34119_);
  nor (_34126_, _11244_, _13557_);
  or (_34127_, _34126_, _34037_);
  and (_34128_, _34127_, _06535_);
  or (_34129_, _34128_, _06559_);
  or (_34130_, _34129_, _34125_);
  or (_34132_, _34047_, _07240_);
  and (_34133_, _34132_, _05933_);
  and (_34134_, _34133_, _34130_);
  and (_34135_, _34043_, _05932_);
  or (_34136_, _34135_, _06566_);
  or (_34137_, _34136_, _34134_);
  and (_34138_, _15296_, _07881_);
  or (_34139_, _34037_, _06570_);
  or (_34140_, _34139_, _34138_);
  and (_34141_, _34140_, _01320_);
  and (_34143_, _34141_, _34137_);
  or (_34144_, _34143_, _34036_);
  and (_43047_, _34144_, _42355_);
  and (_34145_, _01324_, \oc8051_golden_model_1.IE [5]);
  and (_34146_, _13557_, \oc8051_golden_model_1.IE [5]);
  and (_34147_, _15330_, _07881_);
  or (_34148_, _34147_, _34146_);
  or (_34149_, _34148_, _06286_);
  and (_34150_, _07881_, \oc8051_golden_model_1.ACC [5]);
  or (_34151_, _34150_, _34146_);
  and (_34153_, _34151_, _07143_);
  and (_34154_, _07144_, \oc8051_golden_model_1.IE [5]);
  or (_34155_, _34154_, _06285_);
  or (_34156_, _34155_, _34153_);
  and (_34157_, _34156_, _06282_);
  and (_34158_, _34157_, _34149_);
  and (_34159_, _13562_, \oc8051_golden_model_1.IE [5]);
  and (_34160_, _15315_, _08609_);
  or (_34161_, _34160_, _34159_);
  and (_34162_, _34161_, _06281_);
  or (_34164_, _34162_, _06354_);
  or (_34165_, _34164_, _34158_);
  and (_34166_, _09419_, _07881_);
  or (_34167_, _34166_, _34146_);
  or (_34168_, _34167_, _07169_);
  and (_34169_, _34168_, _34165_);
  or (_34170_, _34169_, _06345_);
  or (_34171_, _34151_, _06346_);
  and (_34172_, _34171_, _06278_);
  and (_34173_, _34172_, _34170_);
  and (_34175_, _15342_, _08609_);
  or (_34176_, _34175_, _34159_);
  and (_34177_, _34176_, _06277_);
  or (_34178_, _34177_, _06270_);
  or (_34179_, _34178_, _34173_);
  or (_34180_, _34159_, _15349_);
  and (_34181_, _34180_, _34161_);
  or (_34182_, _34181_, _06271_);
  and (_34184_, _34182_, _06267_);
  and (_34186_, _34184_, _34179_);
  or (_34189_, _34159_, _15365_);
  and (_34191_, _34189_, _06266_);
  and (_34193_, _34191_, _34161_);
  or (_34195_, _34193_, _06259_);
  or (_34197_, _34195_, _34186_);
  or (_34199_, _34167_, _06260_);
  and (_34201_, _34199_, _34197_);
  or (_34203_, _34201_, _09486_);
  and (_34204_, _09436_, _07881_);
  or (_34205_, _34146_, _06258_);
  or (_34207_, _34205_, _34204_);
  and (_34208_, _34207_, _06251_);
  and (_34209_, _34208_, _34203_);
  and (_34210_, _15421_, _07881_);
  or (_34211_, _34210_, _34146_);
  and (_34212_, _34211_, _05972_);
  or (_34213_, _34212_, _10080_);
  or (_34214_, _34213_, _34209_);
  and (_34215_, _15313_, _07881_);
  or (_34216_, _34146_, _09025_);
  or (_34218_, _34216_, _34215_);
  and (_34219_, _08913_, _07881_);
  or (_34220_, _34219_, _34146_);
  or (_34221_, _34220_, _06216_);
  and (_34222_, _34221_, _09030_);
  and (_34223_, _34222_, _34218_);
  and (_34224_, _34223_, _34214_);
  and (_34225_, _12536_, _07881_);
  or (_34226_, _34225_, _34146_);
  and (_34227_, _34226_, _06524_);
  or (_34229_, _34227_, _34224_);
  and (_34230_, _34229_, _07219_);
  or (_34231_, _34146_, _08231_);
  and (_34232_, _34220_, _06426_);
  and (_34233_, _34232_, _34231_);
  or (_34234_, _34233_, _34230_);
  and (_34235_, _34234_, _07217_);
  and (_34236_, _34151_, _06532_);
  and (_34237_, _34236_, _34231_);
  or (_34238_, _34237_, _06437_);
  or (_34240_, _34238_, _34235_);
  and (_34241_, _15310_, _07881_);
  or (_34242_, _34146_, _07229_);
  or (_34243_, _34242_, _34241_);
  and (_34244_, _34243_, _07231_);
  and (_34245_, _34244_, _34240_);
  nor (_34246_, _11241_, _13557_);
  or (_34247_, _34246_, _34146_);
  and (_34248_, _34247_, _06535_);
  or (_34249_, _34248_, _06559_);
  or (_34251_, _34249_, _34245_);
  or (_34252_, _34148_, _07240_);
  and (_34253_, _34252_, _05933_);
  and (_34254_, _34253_, _34251_);
  and (_34255_, _34176_, _05932_);
  or (_34256_, _34255_, _06566_);
  or (_34257_, _34256_, _34254_);
  and (_34258_, _15493_, _07881_);
  or (_34259_, _34146_, _06570_);
  or (_34260_, _34259_, _34258_);
  and (_34262_, _34260_, _01320_);
  and (_34263_, _34262_, _34257_);
  or (_34264_, _34263_, _34145_);
  and (_43048_, _34264_, _42355_);
  and (_34265_, _01324_, \oc8051_golden_model_1.IE [6]);
  and (_34266_, _13557_, \oc8051_golden_model_1.IE [6]);
  and (_34267_, _15521_, _07881_);
  or (_34268_, _34267_, _34266_);
  or (_34269_, _34268_, _06286_);
  and (_34270_, _07881_, \oc8051_golden_model_1.ACC [6]);
  or (_34272_, _34270_, _34266_);
  and (_34273_, _34272_, _07143_);
  and (_34274_, _07144_, \oc8051_golden_model_1.IE [6]);
  or (_34275_, _34274_, _06285_);
  or (_34276_, _34275_, _34273_);
  and (_34277_, _34276_, _06282_);
  and (_34278_, _34277_, _34269_);
  and (_34279_, _13562_, \oc8051_golden_model_1.IE [6]);
  and (_34280_, _15535_, _08609_);
  or (_34281_, _34280_, _34279_);
  and (_34283_, _34281_, _06281_);
  or (_34284_, _34283_, _06354_);
  or (_34285_, _34284_, _34278_);
  and (_34286_, _09418_, _07881_);
  or (_34287_, _34286_, _34266_);
  or (_34288_, _34287_, _07169_);
  and (_34289_, _34288_, _34285_);
  or (_34290_, _34289_, _06345_);
  or (_34291_, _34272_, _06346_);
  and (_34292_, _34291_, _06278_);
  and (_34294_, _34292_, _34290_);
  and (_34295_, _15544_, _08609_);
  or (_34296_, _34295_, _34279_);
  and (_34297_, _34296_, _06277_);
  or (_34298_, _34297_, _06270_);
  or (_34299_, _34298_, _34294_);
  or (_34300_, _34279_, _15551_);
  and (_34301_, _34300_, _34281_);
  or (_34302_, _34301_, _06271_);
  and (_34303_, _34302_, _06267_);
  and (_34305_, _34303_, _34299_);
  and (_34306_, _15568_, _08609_);
  or (_34307_, _34306_, _34279_);
  and (_34308_, _34307_, _06266_);
  or (_34309_, _34308_, _06259_);
  or (_34310_, _34309_, _34305_);
  or (_34311_, _34287_, _06260_);
  and (_34312_, _34311_, _34310_);
  or (_34313_, _34312_, _09486_);
  and (_34314_, _09435_, _07881_);
  or (_34316_, _34266_, _06258_);
  or (_34317_, _34316_, _34314_);
  and (_34318_, _34317_, _06251_);
  and (_34319_, _34318_, _34313_);
  and (_34320_, _15623_, _07881_);
  or (_34321_, _34320_, _34266_);
  and (_34322_, _34321_, _05972_);
  or (_34323_, _34322_, _10080_);
  or (_34324_, _34323_, _34319_);
  and (_34325_, _15517_, _07881_);
  or (_34327_, _34266_, _09025_);
  or (_34328_, _34327_, _34325_);
  and (_34329_, _08845_, _07881_);
  or (_34330_, _34329_, _34266_);
  or (_34331_, _34330_, _06216_);
  and (_34332_, _34331_, _09030_);
  and (_34333_, _34332_, _34328_);
  and (_34334_, _34333_, _34324_);
  and (_34335_, _11239_, _07881_);
  or (_34336_, _34335_, _34266_);
  and (_34338_, _34336_, _06524_);
  or (_34339_, _34338_, _34334_);
  and (_34340_, _34339_, _07219_);
  or (_34341_, _34266_, _08128_);
  and (_34342_, _34330_, _06426_);
  and (_34343_, _34342_, _34341_);
  or (_34344_, _34343_, _34340_);
  and (_34345_, _34344_, _07217_);
  and (_34346_, _34272_, _06532_);
  and (_34347_, _34346_, _34341_);
  or (_34349_, _34347_, _06437_);
  or (_34350_, _34349_, _34345_);
  and (_34351_, _15514_, _07881_);
  or (_34352_, _34266_, _07229_);
  or (_34353_, _34352_, _34351_);
  and (_34354_, _34353_, _07231_);
  and (_34355_, _34354_, _34350_);
  nor (_34356_, _11238_, _13557_);
  or (_34357_, _34356_, _34266_);
  and (_34358_, _34357_, _06535_);
  or (_34360_, _34358_, _06559_);
  or (_34361_, _34360_, _34355_);
  or (_34362_, _34268_, _07240_);
  and (_34363_, _34362_, _05933_);
  and (_34364_, _34363_, _34361_);
  and (_34365_, _34296_, _05932_);
  or (_34366_, _34365_, _06566_);
  or (_34367_, _34366_, _34364_);
  and (_34368_, _15695_, _07881_);
  or (_34369_, _34266_, _06570_);
  or (_34371_, _34369_, _34368_);
  and (_34372_, _34371_, _01320_);
  and (_34373_, _34372_, _34367_);
  or (_34374_, _34373_, _34265_);
  and (_43049_, _34374_, _42355_);
  not (_34375_, \oc8051_golden_model_1.SCON [0]);
  nor (_34376_, _01320_, _34375_);
  nand (_34377_, _11254_, _07963_);
  nor (_34378_, _07963_, _34375_);
  nor (_34379_, _34378_, _07217_);
  nand (_34381_, _34379_, _34377_);
  and (_34382_, _07963_, _07135_);
  or (_34383_, _34382_, _34378_);
  or (_34384_, _34383_, _06260_);
  nor (_34385_, _08374_, _13664_);
  or (_34386_, _34385_, _34378_);
  and (_34387_, _34386_, _06285_);
  nor (_34388_, _07143_, _34375_);
  and (_34389_, _07963_, \oc8051_golden_model_1.ACC [0]);
  or (_34390_, _34389_, _34378_);
  and (_34392_, _34390_, _07143_);
  or (_34393_, _34392_, _34388_);
  and (_34394_, _34393_, _06286_);
  or (_34395_, _34394_, _06281_);
  or (_34396_, _34395_, _34387_);
  and (_34397_, _14326_, _08612_);
  nor (_34398_, _08612_, _34375_);
  or (_34399_, _34398_, _06282_);
  or (_34400_, _34399_, _34397_);
  and (_34401_, _34400_, _07169_);
  and (_34403_, _34401_, _34396_);
  and (_34404_, _34383_, _06354_);
  or (_34405_, _34404_, _06345_);
  or (_34406_, _34405_, _34403_);
  or (_34407_, _34390_, _06346_);
  and (_34408_, _34407_, _06278_);
  and (_34409_, _34408_, _34406_);
  and (_34410_, _34378_, _06277_);
  or (_34411_, _34410_, _06270_);
  or (_34412_, _34411_, _34409_);
  or (_34414_, _34386_, _06271_);
  and (_34415_, _34414_, _06267_);
  and (_34416_, _34415_, _34412_);
  and (_34417_, _14358_, _08612_);
  or (_34418_, _34417_, _34398_);
  and (_34419_, _34418_, _06266_);
  or (_34420_, _34419_, _06259_);
  or (_34421_, _34420_, _34416_);
  and (_34422_, _34421_, _34384_);
  or (_34423_, _34422_, _09486_);
  and (_34425_, _09384_, _07963_);
  or (_34426_, _34378_, _06258_);
  or (_34427_, _34426_, _34425_);
  and (_34428_, _34427_, _06251_);
  and (_34429_, _34428_, _34423_);
  and (_34430_, _14413_, _07963_);
  or (_34431_, _34430_, _34378_);
  and (_34432_, _34431_, _05972_);
  or (_34433_, _34432_, _34429_);
  or (_34434_, _34433_, _10080_);
  and (_34436_, _14311_, _07963_);
  or (_34437_, _34378_, _09025_);
  or (_34438_, _34437_, _34436_);
  and (_34439_, _07963_, _08929_);
  or (_34440_, _34439_, _34378_);
  or (_34441_, _34440_, _06216_);
  and (_34442_, _34441_, _09030_);
  and (_34443_, _34442_, _34438_);
  and (_34444_, _34443_, _34434_);
  nor (_34445_, _12532_, _13664_);
  or (_34447_, _34445_, _34378_);
  and (_34448_, _34377_, _06524_);
  and (_34449_, _34448_, _34447_);
  or (_34450_, _34449_, _34444_);
  and (_34451_, _34450_, _07219_);
  nand (_34452_, _34440_, _06426_);
  nor (_34453_, _34452_, _34385_);
  or (_34454_, _34453_, _06532_);
  or (_34455_, _34454_, _34451_);
  and (_34456_, _34455_, _34381_);
  or (_34458_, _34456_, _06437_);
  and (_34459_, _14307_, _07963_);
  or (_34460_, _34378_, _07229_);
  or (_34461_, _34460_, _34459_);
  and (_34462_, _34461_, _07231_);
  and (_34463_, _34462_, _34458_);
  and (_34464_, _34447_, _06535_);
  or (_34465_, _34464_, _06559_);
  or (_34466_, _34465_, _34463_);
  or (_34467_, _34386_, _07240_);
  and (_34469_, _34467_, _34466_);
  or (_34470_, _34469_, _05932_);
  or (_34471_, _34378_, _05933_);
  and (_34472_, _34471_, _34470_);
  or (_34473_, _34472_, _06566_);
  or (_34474_, _34386_, _06570_);
  and (_34475_, _34474_, _01320_);
  and (_34476_, _34475_, _34473_);
  or (_34477_, _34476_, _34376_);
  and (_43051_, _34477_, _42355_);
  not (_34479_, \oc8051_golden_model_1.SCON [1]);
  nor (_34480_, _01320_, _34479_);
  nor (_34481_, _07963_, _34479_);
  and (_34482_, _07963_, _09422_);
  or (_34483_, _34482_, _34481_);
  or (_34484_, _34483_, _07169_);
  or (_34485_, _07963_, \oc8051_golden_model_1.SCON [1]);
  and (_34486_, _14520_, _07963_);
  not (_34487_, _34486_);
  and (_34488_, _34487_, _34485_);
  or (_34490_, _34488_, _06286_);
  and (_34491_, _07963_, \oc8051_golden_model_1.ACC [1]);
  or (_34492_, _34491_, _34481_);
  and (_34493_, _34492_, _07143_);
  nor (_34494_, _07143_, _34479_);
  or (_34495_, _34494_, _06285_);
  or (_34496_, _34495_, _34493_);
  and (_34497_, _34496_, _06282_);
  and (_34498_, _34497_, _34490_);
  nor (_34499_, _08612_, _34479_);
  and (_34501_, _14508_, _08612_);
  or (_34502_, _34501_, _34499_);
  and (_34503_, _34502_, _06281_);
  or (_34504_, _34503_, _06354_);
  or (_34505_, _34504_, _34498_);
  and (_34506_, _34505_, _34484_);
  or (_34507_, _34506_, _06345_);
  or (_34508_, _34492_, _06346_);
  and (_34509_, _34508_, _06278_);
  and (_34510_, _34509_, _34507_);
  and (_34512_, _14511_, _08612_);
  or (_34513_, _34512_, _34499_);
  and (_34514_, _34513_, _06277_);
  or (_34515_, _34514_, _06270_);
  or (_34516_, _34515_, _34510_);
  and (_34517_, _34501_, _14507_);
  or (_34518_, _34499_, _06271_);
  or (_34519_, _34518_, _34517_);
  and (_34520_, _34519_, _06267_);
  and (_34521_, _34520_, _34516_);
  or (_34523_, _34499_, _14551_);
  and (_34524_, _34523_, _06266_);
  and (_34525_, _34524_, _34502_);
  or (_34526_, _34525_, _06259_);
  or (_34527_, _34526_, _34521_);
  or (_34528_, _34483_, _06260_);
  and (_34529_, _34528_, _34527_);
  or (_34530_, _34529_, _09486_);
  and (_34531_, _09339_, _07963_);
  or (_34532_, _34481_, _06258_);
  or (_34534_, _34532_, _34531_);
  and (_34535_, _34534_, _06251_);
  and (_34536_, _34535_, _34530_);
  and (_34537_, _14607_, _07963_);
  or (_34538_, _34537_, _34481_);
  and (_34539_, _34538_, _05972_);
  or (_34540_, _34539_, _34536_);
  and (_34541_, _34540_, _06399_);
  or (_34542_, _14505_, _13664_);
  and (_34543_, _34485_, _06398_);
  and (_34545_, _34543_, _34542_);
  nand (_34546_, _07963_, _07031_);
  and (_34547_, _34546_, _06215_);
  and (_34548_, _34547_, _34485_);
  or (_34549_, _34548_, _06524_);
  or (_34550_, _34549_, _34545_);
  or (_34551_, _34550_, _34541_);
  nor (_34552_, _11252_, _13664_);
  or (_34553_, _34552_, _34481_);
  nand (_34554_, _11251_, _07963_);
  and (_34556_, _34554_, _34553_);
  or (_34557_, _34556_, _09030_);
  and (_34558_, _34557_, _07219_);
  and (_34559_, _34558_, _34551_);
  or (_34560_, _14503_, _13664_);
  and (_34561_, _34485_, _06426_);
  and (_34562_, _34561_, _34560_);
  or (_34563_, _34562_, _06532_);
  or (_34564_, _34563_, _34559_);
  nor (_34565_, _34481_, _07217_);
  nand (_34567_, _34565_, _34554_);
  and (_34568_, _34567_, _07229_);
  and (_34569_, _34568_, _34564_);
  or (_34570_, _34546_, _08325_);
  and (_34571_, _34485_, _06437_);
  and (_34572_, _34571_, _34570_);
  or (_34573_, _34572_, _06535_);
  or (_34574_, _34573_, _34569_);
  or (_34575_, _34553_, _07231_);
  and (_34576_, _34575_, _34574_);
  or (_34578_, _34576_, _06559_);
  or (_34579_, _34488_, _07240_);
  and (_34580_, _34579_, _05933_);
  and (_34581_, _34580_, _34578_);
  and (_34582_, _34513_, _05932_);
  or (_34583_, _34582_, _06566_);
  or (_34584_, _34583_, _34581_);
  or (_34585_, _34481_, _06570_);
  or (_34586_, _34585_, _34486_);
  and (_34587_, _34586_, _01320_);
  and (_34589_, _34587_, _34584_);
  or (_34590_, _34589_, _34480_);
  and (_43052_, _34590_, _42355_);
  and (_34591_, _01324_, \oc8051_golden_model_1.SCON [2]);
  and (_34592_, _13664_, \oc8051_golden_model_1.SCON [2]);
  and (_34593_, _07963_, _08662_);
  or (_34594_, _34593_, _34592_);
  or (_34595_, _34594_, _06260_);
  or (_34596_, _34594_, _07169_);
  and (_34597_, _14703_, _07963_);
  or (_34599_, _34597_, _34592_);
  or (_34600_, _34599_, _06286_);
  and (_34601_, _07963_, \oc8051_golden_model_1.ACC [2]);
  or (_34602_, _34601_, _34592_);
  and (_34603_, _34602_, _07143_);
  and (_34604_, _07144_, \oc8051_golden_model_1.SCON [2]);
  or (_34605_, _34604_, _06285_);
  or (_34606_, _34605_, _34603_);
  and (_34607_, _34606_, _06282_);
  and (_34608_, _34607_, _34600_);
  and (_34610_, _13669_, \oc8051_golden_model_1.SCON [2]);
  and (_34611_, _14716_, _08612_);
  or (_34612_, _34611_, _34610_);
  and (_34613_, _34612_, _06281_);
  or (_34614_, _34613_, _06354_);
  or (_34615_, _34614_, _34608_);
  and (_34616_, _34615_, _34596_);
  or (_34617_, _34616_, _06345_);
  or (_34618_, _34602_, _06346_);
  and (_34619_, _34618_, _06278_);
  and (_34621_, _34619_, _34617_);
  and (_34622_, _14699_, _08612_);
  or (_34623_, _34622_, _34610_);
  and (_34624_, _34623_, _06277_);
  or (_34625_, _34624_, _06270_);
  or (_34626_, _34625_, _34621_);
  and (_34627_, _34611_, _14731_);
  or (_34628_, _34610_, _06271_);
  or (_34629_, _34628_, _34627_);
  and (_34630_, _34629_, _06267_);
  and (_34632_, _34630_, _34626_);
  and (_34633_, _14749_, _08612_);
  or (_34634_, _34633_, _34610_);
  and (_34635_, _34634_, _06266_);
  or (_34636_, _34635_, _06259_);
  or (_34637_, _34636_, _34632_);
  and (_34638_, _34637_, _34595_);
  or (_34639_, _34638_, _09486_);
  and (_34640_, _09293_, _07963_);
  or (_34641_, _34592_, _06258_);
  or (_34643_, _34641_, _34640_);
  and (_34644_, _34643_, _06251_);
  and (_34645_, _34644_, _34639_);
  and (_34646_, _14804_, _07963_);
  or (_34647_, _34592_, _34646_);
  and (_34648_, _34647_, _05972_);
  or (_34649_, _34648_, _34645_);
  or (_34650_, _34649_, _10080_);
  and (_34651_, _14697_, _07963_);
  or (_34652_, _34592_, _09025_);
  or (_34654_, _34652_, _34651_);
  and (_34655_, _07963_, _08980_);
  or (_34656_, _34655_, _34592_);
  or (_34657_, _34656_, _06216_);
  and (_34658_, _34657_, _09030_);
  and (_34659_, _34658_, _34654_);
  and (_34660_, _34659_, _34650_);
  and (_34661_, _11250_, _07963_);
  or (_34662_, _34661_, _34592_);
  and (_34663_, _34662_, _06524_);
  or (_34665_, _34663_, _34660_);
  and (_34666_, _34665_, _07219_);
  or (_34667_, _34592_, _08424_);
  and (_34668_, _34656_, _06426_);
  and (_34669_, _34668_, _34667_);
  or (_34670_, _34669_, _34666_);
  and (_34671_, _34670_, _07217_);
  and (_34672_, _34602_, _06532_);
  and (_34673_, _34672_, _34667_);
  or (_34674_, _34673_, _06437_);
  or (_34676_, _34674_, _34671_);
  and (_34677_, _14694_, _07963_);
  or (_34678_, _34592_, _07229_);
  or (_34679_, _34678_, _34677_);
  and (_34680_, _34679_, _07231_);
  and (_34681_, _34680_, _34676_);
  nor (_34682_, _11249_, _13664_);
  or (_34683_, _34682_, _34592_);
  and (_34684_, _34683_, _06535_);
  or (_34685_, _34684_, _06559_);
  or (_34687_, _34685_, _34681_);
  or (_34688_, _34599_, _07240_);
  and (_34689_, _34688_, _05933_);
  and (_34690_, _34689_, _34687_);
  and (_34691_, _34623_, _05932_);
  or (_34692_, _34691_, _06566_);
  or (_34693_, _34692_, _34690_);
  and (_34694_, _14873_, _07963_);
  or (_34695_, _34592_, _06570_);
  or (_34696_, _34695_, _34694_);
  and (_34698_, _34696_, _01320_);
  and (_34699_, _34698_, _34693_);
  or (_34700_, _34699_, _34591_);
  and (_43053_, _34700_, _42355_);
  and (_34701_, _01324_, \oc8051_golden_model_1.SCON [3]);
  and (_34702_, _13664_, \oc8051_golden_model_1.SCON [3]);
  and (_34703_, _07963_, _09421_);
  or (_34704_, _34703_, _34702_);
  or (_34705_, _34704_, _06260_);
  and (_34706_, _14900_, _07963_);
  or (_34708_, _34706_, _34702_);
  or (_34709_, _34708_, _06286_);
  and (_34710_, _07963_, \oc8051_golden_model_1.ACC [3]);
  or (_34711_, _34710_, _34702_);
  and (_34712_, _34711_, _07143_);
  and (_34713_, _07144_, \oc8051_golden_model_1.SCON [3]);
  or (_34714_, _34713_, _06285_);
  or (_34715_, _34714_, _34712_);
  and (_34716_, _34715_, _06282_);
  and (_34717_, _34716_, _34709_);
  and (_34719_, _13669_, \oc8051_golden_model_1.SCON [3]);
  and (_34720_, _14897_, _08612_);
  or (_34721_, _34720_, _34719_);
  and (_34722_, _34721_, _06281_);
  or (_34723_, _34722_, _06354_);
  or (_34724_, _34723_, _34717_);
  or (_34725_, _34704_, _07169_);
  and (_34726_, _34725_, _34724_);
  or (_34727_, _34726_, _06345_);
  or (_34728_, _34711_, _06346_);
  and (_34730_, _34728_, _06278_);
  and (_34731_, _34730_, _34727_);
  and (_34732_, _14895_, _08612_);
  or (_34733_, _34732_, _34719_);
  and (_34734_, _34733_, _06277_);
  or (_34735_, _34734_, _06270_);
  or (_34736_, _34735_, _34731_);
  or (_34737_, _34719_, _14926_);
  and (_34738_, _34737_, _34721_);
  or (_34739_, _34738_, _06271_);
  and (_34741_, _34739_, _06267_);
  and (_34742_, _34741_, _34736_);
  and (_34743_, _14943_, _08612_);
  or (_34744_, _34743_, _34719_);
  and (_34745_, _34744_, _06266_);
  or (_34746_, _34745_, _06259_);
  or (_34747_, _34746_, _34742_);
  and (_34748_, _34747_, _34705_);
  or (_34749_, _34748_, _09486_);
  and (_34750_, _09247_, _07963_);
  or (_34752_, _34702_, _06258_);
  or (_34753_, _34752_, _34750_);
  and (_34754_, _34753_, _06251_);
  and (_34755_, _34754_, _34749_);
  and (_34756_, _14998_, _07963_);
  or (_34757_, _34702_, _34756_);
  and (_34758_, _34757_, _05972_);
  or (_34759_, _34758_, _34755_);
  or (_34760_, _34759_, _10080_);
  and (_34761_, _14893_, _07963_);
  or (_34762_, _34702_, _09025_);
  or (_34763_, _34762_, _34761_);
  and (_34764_, _07963_, _08809_);
  or (_34765_, _34764_, _34702_);
  or (_34766_, _34765_, _06216_);
  and (_34767_, _34766_, _09030_);
  and (_34768_, _34767_, _34763_);
  and (_34769_, _34768_, _34760_);
  and (_34770_, _12529_, _07963_);
  or (_34771_, _34770_, _34702_);
  and (_34773_, _34771_, _06524_);
  or (_34774_, _34773_, _34769_);
  and (_34775_, _34774_, _07219_);
  or (_34776_, _34702_, _08280_);
  and (_34777_, _34765_, _06426_);
  and (_34778_, _34777_, _34776_);
  or (_34779_, _34778_, _34775_);
  and (_34780_, _34779_, _07217_);
  and (_34781_, _34711_, _06532_);
  and (_34782_, _34781_, _34776_);
  or (_34784_, _34782_, _06437_);
  or (_34785_, _34784_, _34780_);
  and (_34786_, _14890_, _07963_);
  or (_34787_, _34702_, _07229_);
  or (_34788_, _34787_, _34786_);
  and (_34789_, _34788_, _07231_);
  and (_34790_, _34789_, _34785_);
  nor (_34791_, _11247_, _13664_);
  or (_34792_, _34791_, _34702_);
  and (_34793_, _34792_, _06535_);
  or (_34795_, _34793_, _06559_);
  or (_34796_, _34795_, _34790_);
  or (_34797_, _34708_, _07240_);
  and (_34798_, _34797_, _05933_);
  and (_34799_, _34798_, _34796_);
  and (_34800_, _34733_, _05932_);
  or (_34801_, _34800_, _06566_);
  or (_34802_, _34801_, _34799_);
  and (_34803_, _15068_, _07963_);
  or (_34804_, _34702_, _06570_);
  or (_34806_, _34804_, _34803_);
  and (_34807_, _34806_, _01320_);
  and (_34808_, _34807_, _34802_);
  or (_34809_, _34808_, _34701_);
  and (_43054_, _34809_, _42355_);
  and (_34810_, _01324_, \oc8051_golden_model_1.SCON [4]);
  and (_34811_, _13664_, \oc8051_golden_model_1.SCON [4]);
  and (_34812_, _09420_, _07963_);
  or (_34813_, _34812_, _34811_);
  or (_34814_, _34813_, _06260_);
  and (_34816_, _13669_, \oc8051_golden_model_1.SCON [4]);
  and (_34817_, _15145_, _08612_);
  or (_34818_, _34817_, _34816_);
  and (_34819_, _34818_, _06277_);
  and (_34820_, _15133_, _07963_);
  or (_34821_, _34820_, _34811_);
  or (_34822_, _34821_, _06286_);
  and (_34823_, _07963_, \oc8051_golden_model_1.ACC [4]);
  or (_34824_, _34823_, _34811_);
  and (_34825_, _34824_, _07143_);
  and (_34827_, _07144_, \oc8051_golden_model_1.SCON [4]);
  or (_34828_, _34827_, _06285_);
  or (_34829_, _34828_, _34825_);
  and (_34830_, _34829_, _06282_);
  and (_34831_, _34830_, _34822_);
  and (_34832_, _15116_, _08612_);
  or (_34833_, _34832_, _34816_);
  and (_34834_, _34833_, _06281_);
  or (_34835_, _34834_, _06354_);
  or (_34836_, _34835_, _34831_);
  or (_34838_, _34813_, _07169_);
  and (_34839_, _34838_, _34836_);
  or (_34840_, _34839_, _06345_);
  or (_34841_, _34824_, _06346_);
  and (_34842_, _34841_, _06278_);
  and (_34843_, _34842_, _34840_);
  or (_34844_, _34843_, _34819_);
  and (_34845_, _34844_, _06271_);
  or (_34846_, _34816_, _15152_);
  and (_34847_, _34846_, _06270_);
  and (_34849_, _34847_, _34833_);
  or (_34850_, _34849_, _34845_);
  and (_34851_, _34850_, _06267_);
  and (_34852_, _15170_, _08612_);
  or (_34853_, _34852_, _34816_);
  and (_34854_, _34853_, _06266_);
  or (_34855_, _34854_, _06259_);
  or (_34856_, _34855_, _34851_);
  and (_34857_, _34856_, _34814_);
  or (_34858_, _34857_, _09486_);
  and (_34860_, _09437_, _07963_);
  or (_34861_, _34811_, _06258_);
  or (_34862_, _34861_, _34860_);
  and (_34863_, _34862_, _06251_);
  and (_34864_, _34863_, _34858_);
  and (_34865_, _15226_, _07963_);
  or (_34866_, _34865_, _34811_);
  and (_34867_, _34866_, _05972_);
  or (_34868_, _34867_, _10080_);
  or (_34869_, _34868_, _34864_);
  and (_34871_, _15114_, _07963_);
  or (_34872_, _34811_, _09025_);
  or (_34873_, _34872_, _34871_);
  and (_34874_, _08919_, _07963_);
  or (_34875_, _34874_, _34811_);
  or (_34876_, _34875_, _06216_);
  and (_34877_, _34876_, _09030_);
  and (_34878_, _34877_, _34873_);
  and (_34879_, _34878_, _34869_);
  and (_34880_, _11245_, _07963_);
  or (_34882_, _34880_, _34811_);
  and (_34883_, _34882_, _06524_);
  or (_34884_, _34883_, _34879_);
  and (_34885_, _34884_, _07219_);
  or (_34886_, _34811_, _08528_);
  and (_34887_, _34875_, _06426_);
  and (_34888_, _34887_, _34886_);
  or (_34889_, _34888_, _34885_);
  and (_34890_, _34889_, _07217_);
  and (_34891_, _34824_, _06532_);
  and (_34893_, _34891_, _34886_);
  or (_34894_, _34893_, _06437_);
  or (_34895_, _34894_, _34890_);
  and (_34896_, _15111_, _07963_);
  or (_34897_, _34811_, _07229_);
  or (_34898_, _34897_, _34896_);
  and (_34899_, _34898_, _07231_);
  and (_34900_, _34899_, _34895_);
  nor (_34901_, _11244_, _13664_);
  or (_34902_, _34901_, _34811_);
  and (_34904_, _34902_, _06535_);
  or (_34905_, _34904_, _06559_);
  or (_34906_, _34905_, _34900_);
  or (_34907_, _34821_, _07240_);
  and (_34908_, _34907_, _05933_);
  and (_34909_, _34908_, _34906_);
  and (_34910_, _34818_, _05932_);
  or (_34911_, _34910_, _06566_);
  or (_34912_, _34911_, _34909_);
  and (_34913_, _15296_, _07963_);
  or (_34915_, _34811_, _06570_);
  or (_34916_, _34915_, _34913_);
  and (_34917_, _34916_, _01320_);
  and (_34918_, _34917_, _34912_);
  or (_34919_, _34918_, _34810_);
  and (_43055_, _34919_, _42355_);
  and (_34920_, _01324_, \oc8051_golden_model_1.SCON [5]);
  and (_34921_, _13664_, \oc8051_golden_model_1.SCON [5]);
  and (_34922_, _15330_, _07963_);
  or (_34923_, _34922_, _34921_);
  or (_34925_, _34923_, _06286_);
  and (_34926_, _07963_, \oc8051_golden_model_1.ACC [5]);
  or (_34927_, _34926_, _34921_);
  and (_34928_, _34927_, _07143_);
  and (_34929_, _07144_, \oc8051_golden_model_1.SCON [5]);
  or (_34930_, _34929_, _06285_);
  or (_34931_, _34930_, _34928_);
  and (_34932_, _34931_, _06282_);
  and (_34933_, _34932_, _34925_);
  and (_34934_, _13669_, \oc8051_golden_model_1.SCON [5]);
  and (_34936_, _15315_, _08612_);
  or (_34937_, _34936_, _34934_);
  and (_34938_, _34937_, _06281_);
  or (_34939_, _34938_, _06354_);
  or (_34940_, _34939_, _34933_);
  and (_34941_, _09419_, _07963_);
  or (_34942_, _34941_, _34921_);
  or (_34943_, _34942_, _07169_);
  and (_34944_, _34943_, _34940_);
  or (_34945_, _34944_, _06345_);
  or (_34947_, _34927_, _06346_);
  and (_34948_, _34947_, _06278_);
  and (_34949_, _34948_, _34945_);
  and (_34950_, _15342_, _08612_);
  or (_34951_, _34950_, _34934_);
  and (_34952_, _34951_, _06277_);
  or (_34953_, _34952_, _06270_);
  or (_34954_, _34953_, _34949_);
  or (_34955_, _34934_, _15349_);
  and (_34956_, _34955_, _34937_);
  or (_34958_, _34956_, _06271_);
  and (_34959_, _34958_, _06267_);
  and (_34960_, _34959_, _34954_);
  or (_34961_, _34934_, _15365_);
  and (_34962_, _34961_, _06266_);
  and (_34963_, _34962_, _34937_);
  or (_34964_, _34963_, _06259_);
  or (_34965_, _34964_, _34960_);
  or (_34966_, _34942_, _06260_);
  and (_34967_, _34966_, _34965_);
  or (_34969_, _34967_, _09486_);
  and (_34970_, _09436_, _07963_);
  or (_34971_, _34921_, _06258_);
  or (_34972_, _34971_, _34970_);
  and (_34973_, _34972_, _06251_);
  and (_34974_, _34973_, _34969_);
  and (_34975_, _15421_, _07963_);
  or (_34976_, _34975_, _34921_);
  and (_34977_, _34976_, _05972_);
  or (_34978_, _34977_, _10080_);
  or (_34980_, _34978_, _34974_);
  and (_34981_, _15313_, _07963_);
  or (_34982_, _34921_, _09025_);
  or (_34983_, _34982_, _34981_);
  and (_34984_, _08913_, _07963_);
  or (_34985_, _34984_, _34921_);
  or (_34986_, _34985_, _06216_);
  and (_34987_, _34986_, _09030_);
  and (_34988_, _34987_, _34983_);
  and (_34989_, _34988_, _34980_);
  and (_34991_, _12536_, _07963_);
  or (_34992_, _34991_, _34921_);
  and (_34993_, _34992_, _06524_);
  or (_34994_, _34993_, _34989_);
  and (_34995_, _34994_, _07219_);
  or (_34996_, _34921_, _08231_);
  and (_34997_, _34985_, _06426_);
  and (_34998_, _34997_, _34996_);
  or (_34999_, _34998_, _34995_);
  and (_35000_, _34999_, _07217_);
  and (_35002_, _34927_, _06532_);
  and (_35003_, _35002_, _34996_);
  or (_35004_, _35003_, _06437_);
  or (_35005_, _35004_, _35000_);
  and (_35006_, _15310_, _07963_);
  or (_35007_, _34921_, _07229_);
  or (_35008_, _35007_, _35006_);
  and (_35009_, _35008_, _07231_);
  and (_35010_, _35009_, _35005_);
  nor (_35011_, _11241_, _13664_);
  or (_35013_, _35011_, _34921_);
  and (_35014_, _35013_, _06535_);
  or (_35015_, _35014_, _06559_);
  or (_35016_, _35015_, _35010_);
  or (_35017_, _34923_, _07240_);
  and (_35018_, _35017_, _05933_);
  and (_35019_, _35018_, _35016_);
  and (_35020_, _34951_, _05932_);
  or (_35021_, _35020_, _06566_);
  or (_35022_, _35021_, _35019_);
  and (_35024_, _15493_, _07963_);
  or (_35025_, _34921_, _06570_);
  or (_35026_, _35025_, _35024_);
  and (_35027_, _35026_, _01320_);
  and (_35028_, _35027_, _35022_);
  or (_35029_, _35028_, _34920_);
  and (_43056_, _35029_, _42355_);
  and (_35030_, _01324_, \oc8051_golden_model_1.SCON [6]);
  and (_35031_, _13664_, \oc8051_golden_model_1.SCON [6]);
  and (_35032_, _15521_, _07963_);
  or (_35034_, _35032_, _35031_);
  or (_35035_, _35034_, _06286_);
  and (_35036_, _07963_, \oc8051_golden_model_1.ACC [6]);
  or (_35037_, _35036_, _35031_);
  and (_35038_, _35037_, _07143_);
  and (_35039_, _07144_, \oc8051_golden_model_1.SCON [6]);
  or (_35040_, _35039_, _06285_);
  or (_35041_, _35040_, _35038_);
  and (_35042_, _35041_, _06282_);
  and (_35043_, _35042_, _35035_);
  and (_35045_, _13669_, \oc8051_golden_model_1.SCON [6]);
  and (_35046_, _15535_, _08612_);
  or (_35047_, _35046_, _35045_);
  and (_35048_, _35047_, _06281_);
  or (_35049_, _35048_, _06354_);
  or (_35050_, _35049_, _35043_);
  and (_35051_, _09418_, _07963_);
  or (_35052_, _35051_, _35031_);
  or (_35053_, _35052_, _07169_);
  and (_35054_, _35053_, _35050_);
  or (_35056_, _35054_, _06345_);
  or (_35057_, _35037_, _06346_);
  and (_35058_, _35057_, _06278_);
  and (_35059_, _35058_, _35056_);
  and (_35060_, _15544_, _08612_);
  or (_35061_, _35060_, _35045_);
  and (_35062_, _35061_, _06277_);
  or (_35063_, _35062_, _06270_);
  or (_35064_, _35063_, _35059_);
  or (_35065_, _35045_, _15551_);
  and (_35067_, _35065_, _35047_);
  or (_35068_, _35067_, _06271_);
  and (_35069_, _35068_, _06267_);
  and (_35070_, _35069_, _35064_);
  and (_35071_, _15568_, _08612_);
  or (_35072_, _35071_, _35045_);
  and (_35073_, _35072_, _06266_);
  or (_35074_, _35073_, _06259_);
  or (_35075_, _35074_, _35070_);
  or (_35076_, _35052_, _06260_);
  and (_35078_, _35076_, _35075_);
  or (_35079_, _35078_, _09486_);
  and (_35080_, _09435_, _07963_);
  or (_35081_, _35031_, _06258_);
  or (_35082_, _35081_, _35080_);
  and (_35083_, _35082_, _06251_);
  and (_35084_, _35083_, _35079_);
  and (_35085_, _15623_, _07963_);
  or (_35086_, _35085_, _35031_);
  and (_35087_, _35086_, _05972_);
  or (_35089_, _35087_, _10080_);
  or (_35090_, _35089_, _35084_);
  and (_35091_, _15517_, _07963_);
  or (_35092_, _35031_, _09025_);
  or (_35093_, _35092_, _35091_);
  and (_35094_, _08845_, _07963_);
  or (_35095_, _35094_, _35031_);
  or (_35096_, _35095_, _06216_);
  and (_35097_, _35096_, _09030_);
  and (_35098_, _35097_, _35093_);
  and (_35100_, _35098_, _35090_);
  and (_35101_, _11239_, _07963_);
  or (_35102_, _35101_, _35031_);
  and (_35103_, _35102_, _06524_);
  or (_35104_, _35103_, _35100_);
  and (_35105_, _35104_, _07219_);
  or (_35106_, _35031_, _08128_);
  and (_35107_, _35095_, _06426_);
  and (_35108_, _35107_, _35106_);
  or (_35109_, _35108_, _35105_);
  and (_35111_, _35109_, _07217_);
  and (_35112_, _35037_, _06532_);
  and (_35113_, _35112_, _35106_);
  or (_35114_, _35113_, _06437_);
  or (_35115_, _35114_, _35111_);
  and (_35116_, _15514_, _07963_);
  or (_35117_, _35031_, _07229_);
  or (_35118_, _35117_, _35116_);
  and (_35119_, _35118_, _07231_);
  and (_35120_, _35119_, _35115_);
  nor (_35122_, _11238_, _13664_);
  or (_35123_, _35122_, _35031_);
  and (_35124_, _35123_, _06535_);
  or (_35125_, _35124_, _06559_);
  or (_35126_, _35125_, _35120_);
  or (_35127_, _35034_, _07240_);
  and (_35128_, _35127_, _05933_);
  and (_35129_, _35128_, _35126_);
  and (_35130_, _35061_, _05932_);
  or (_35131_, _35130_, _06566_);
  or (_35133_, _35131_, _35129_);
  and (_35134_, _15695_, _07963_);
  or (_35135_, _35031_, _06570_);
  or (_35136_, _35135_, _35134_);
  and (_35137_, _35136_, _01320_);
  and (_35138_, _35137_, _35133_);
  or (_35139_, _35138_, _35030_);
  and (_43057_, _35139_, _42355_);
  nor (_35140_, _01320_, _06766_);
  nor (_35141_, _07919_, _06766_);
  and (_35143_, _07919_, \oc8051_golden_model_1.ACC [0]);
  and (_35144_, _35143_, _08374_);
  or (_35145_, _35144_, _35141_);
  or (_35146_, _35145_, _07217_);
  nor (_35147_, _08374_, _13879_);
  or (_35148_, _35147_, _35141_);
  or (_35149_, _35148_, _06286_);
  or (_35150_, _35143_, _35141_);
  and (_35151_, _35150_, _07143_);
  nor (_35152_, _07143_, _06766_);
  or (_35154_, _35152_, _06285_);
  or (_35155_, _35154_, _35151_);
  and (_35156_, _35155_, _07169_);
  nand (_35157_, _35156_, _35149_);
  nand (_35158_, _35157_, _06768_);
  or (_35159_, _35150_, _06346_);
  and (_35160_, _35159_, _06778_);
  and (_35161_, _35160_, _35158_);
  or (_35162_, _06259_, _07185_);
  or (_35163_, _35162_, _35161_);
  and (_35165_, _08256_, _07135_);
  or (_35166_, _35141_, _06260_);
  or (_35167_, _35166_, _35165_);
  and (_35168_, _35167_, _35163_);
  or (_35169_, _35168_, _09486_);
  or (_35170_, _35141_, _06258_);
  and (_35171_, _09384_, _07919_);
  or (_35172_, _35171_, _35170_);
  and (_35173_, _35172_, _35169_);
  or (_35174_, _35173_, _05972_);
  and (_35176_, _14413_, _08256_);
  or (_35177_, _35141_, _06251_);
  or (_35178_, _35177_, _35176_);
  and (_35179_, _35178_, _06216_);
  and (_35180_, _35179_, _35174_);
  and (_35181_, _07919_, _08929_);
  or (_35182_, _35181_, _35141_);
  and (_35183_, _35182_, _06215_);
  or (_35184_, _35183_, _06398_);
  or (_35185_, _35184_, _35180_);
  and (_35187_, _14311_, _07919_);
  or (_35188_, _35187_, _35141_);
  or (_35189_, _35188_, _09025_);
  and (_35190_, _35189_, _09030_);
  and (_35191_, _35190_, _35185_);
  nor (_35192_, _12532_, _13879_);
  or (_35193_, _35192_, _35141_);
  nor (_35194_, _35144_, _09030_);
  and (_35195_, _35194_, _35193_);
  or (_35196_, _35195_, _35191_);
  and (_35198_, _35196_, _07219_);
  nand (_35199_, _35182_, _06426_);
  nor (_35200_, _35199_, _35147_);
  or (_35201_, _35200_, _06532_);
  or (_35202_, _35201_, _35198_);
  and (_35203_, _35202_, _35146_);
  or (_35204_, _35203_, _06437_);
  and (_35205_, _14307_, _07919_);
  or (_35206_, _35205_, _35141_);
  or (_35207_, _35206_, _07229_);
  and (_35209_, _35207_, _07231_);
  and (_35210_, _35209_, _35204_);
  and (_35211_, _35193_, _06535_);
  or (_35212_, _35211_, _19480_);
  or (_35213_, _35212_, _35210_);
  or (_35214_, _35148_, _06651_);
  and (_35215_, _35214_, _01320_);
  and (_35216_, _35215_, _35213_);
  or (_35217_, _35216_, _35140_);
  and (_43059_, _35217_, _42355_);
  nand (_35219_, _08256_, _07031_);
  or (_35220_, _35219_, _08325_);
  or (_35221_, _07919_, \oc8051_golden_model_1.SP [1]);
  and (_35222_, _35221_, _06437_);
  and (_35223_, _35222_, _35220_);
  and (_35224_, _11251_, _08256_);
  nor (_35225_, _07919_, _07271_);
  or (_35226_, _35225_, _07217_);
  or (_35227_, _35226_, _35224_);
  and (_35228_, _14520_, _08256_);
  not (_35230_, _35228_);
  and (_35231_, _35230_, _35221_);
  or (_35232_, _35231_, _06286_);
  nand (_35233_, _07152_, \oc8051_golden_model_1.SP [1]);
  and (_35234_, _07919_, \oc8051_golden_model_1.ACC [1]);
  or (_35235_, _35234_, _35225_);
  and (_35236_, _35235_, _07143_);
  nor (_35237_, _07143_, _07271_);
  or (_35238_, _35237_, _07152_);
  or (_35239_, _35238_, _35236_);
  and (_35241_, _35239_, _35233_);
  or (_35242_, _35241_, _06285_);
  and (_35243_, _35242_, _05949_);
  and (_35244_, _35243_, _35232_);
  nor (_35245_, _05949_, \oc8051_golden_model_1.SP [1]);
  or (_35246_, _35245_, _06354_);
  or (_35247_, _35246_, _35244_);
  nand (_35248_, _07275_, _06354_);
  and (_35249_, _35248_, _35247_);
  or (_35250_, _35249_, _06345_);
  or (_35252_, _35235_, _06346_);
  and (_35253_, _35252_, _06778_);
  and (_35254_, _35253_, _35250_);
  not (_35255_, _07459_);
  or (_35256_, _35255_, _07279_);
  or (_35257_, _35256_, _35254_);
  or (_35258_, _07459_, _07271_);
  and (_35259_, _35258_, _06260_);
  and (_35260_, _35259_, _35257_);
  or (_35261_, _13879_, _09422_);
  and (_35263_, _35221_, _06259_);
  and (_35264_, _35263_, _35261_);
  or (_35265_, _35264_, _09486_);
  or (_35266_, _35265_, _35260_);
  or (_35267_, _35225_, _06258_);
  and (_35268_, _09339_, _07919_);
  or (_35269_, _35268_, _35267_);
  and (_35270_, _35269_, _06251_);
  and (_35271_, _35270_, _35266_);
  and (_35272_, _35221_, _05972_);
  or (_35274_, _14607_, _13879_);
  and (_35275_, _35274_, _35272_);
  or (_35276_, _35275_, _35271_);
  and (_35277_, _35276_, _06216_);
  and (_35278_, _35221_, _06215_);
  and (_35279_, _35278_, _35219_);
  or (_35280_, _35279_, _06004_);
  or (_35281_, _35280_, _35277_);
  and (_35282_, _06004_, \oc8051_golden_model_1.SP [1]);
  nor (_35283_, _35282_, _06398_);
  and (_35285_, _35283_, _35281_);
  or (_35286_, _14505_, _13879_);
  and (_35287_, _35221_, _06398_);
  and (_35288_, _35287_, _35286_);
  or (_35289_, _35288_, _06524_);
  or (_35290_, _35289_, _35285_);
  and (_35291_, _11253_, _07919_);
  or (_35292_, _35291_, _35225_);
  or (_35293_, _35292_, _09030_);
  and (_35294_, _35293_, _07219_);
  and (_35296_, _35294_, _35290_);
  or (_35297_, _14503_, _13879_);
  and (_35298_, _35221_, _06426_);
  and (_35299_, _35298_, _35297_);
  or (_35300_, _35299_, _06532_);
  or (_35301_, _35300_, _35296_);
  and (_35302_, _35301_, _35227_);
  or (_35303_, _35302_, _06013_);
  and (_35304_, _06013_, \oc8051_golden_model_1.SP [1]);
  nor (_35305_, _35304_, _06437_);
  and (_35307_, _35305_, _35303_);
  or (_35308_, _35307_, _35223_);
  and (_35309_, _35308_, _07231_);
  nor (_35310_, _11252_, _13879_);
  or (_35311_, _35310_, _35225_);
  and (_35312_, _35311_, _06535_);
  or (_35313_, _35312_, _06543_);
  nor (_35314_, _35313_, _35309_);
  or (_35315_, _35314_, _07037_);
  nor (_35316_, _06290_, _06011_);
  nand (_35318_, _35316_, _35315_);
  or (_35319_, _35316_, _07271_);
  and (_35320_, _35319_, _07240_);
  and (_35321_, _35320_, _35318_);
  and (_35322_, _35231_, _06559_);
  or (_35323_, _35322_, _07678_);
  or (_35324_, _35323_, _35321_);
  or (_35325_, _07252_, _07271_);
  and (_35326_, _35325_, _06570_);
  and (_35327_, _35326_, _35324_);
  or (_35329_, _35228_, _35225_);
  and (_35330_, _35329_, _06566_);
  or (_35331_, _35330_, _01324_);
  or (_35332_, _35331_, _35327_);
  or (_35333_, _01320_, \oc8051_golden_model_1.SP [1]);
  and (_35334_, _35333_, _42355_);
  and (_43060_, _35334_, _35332_);
  nor (_35335_, _01320_, _08640_);
  nand (_35336_, _15085_, _06004_);
  and (_35337_, _08256_, _08662_);
  nor (_35339_, _07919_, _08640_);
  or (_35340_, _35339_, _06260_);
  or (_35341_, _35340_, _35337_);
  and (_35342_, _14703_, _08256_);
  or (_35343_, _35342_, _35339_);
  or (_35344_, _35343_, _06286_);
  and (_35345_, _07919_, \oc8051_golden_model_1.ACC [2]);
  or (_35346_, _35345_, _35339_);
  or (_35347_, _35346_, _07144_);
  or (_35348_, _07143_, \oc8051_golden_model_1.SP [2]);
  and (_35350_, _35348_, _07858_);
  and (_35351_, _35350_, _35347_);
  and (_35352_, _07854_, _07152_);
  or (_35353_, _35352_, _06285_);
  or (_35354_, _35353_, _35351_);
  and (_35355_, _35354_, _05949_);
  and (_35356_, _35355_, _35344_);
  nor (_35357_, _15085_, _05949_);
  or (_35358_, _35357_, _06354_);
  or (_35359_, _35358_, _35356_);
  nand (_35361_, _08659_, _06354_);
  and (_35362_, _35361_, _35359_);
  or (_35363_, _35362_, _06345_);
  or (_35364_, _35346_, _06346_);
  and (_35365_, _35364_, _06778_);
  and (_35366_, _35365_, _35363_);
  or (_35367_, _07701_, _07458_);
  or (_35368_, _35367_, _35366_);
  nor (_35369_, _07854_, _05946_);
  nor (_35370_, _35369_, _05974_);
  and (_35372_, _35370_, _35368_);
  and (_35373_, _07854_, _05974_);
  or (_35374_, _35373_, _06259_);
  or (_35375_, _35374_, _35372_);
  and (_35376_, _35375_, _35341_);
  or (_35377_, _35376_, _09486_);
  or (_35378_, _35339_, _06258_);
  and (_35379_, _09293_, _07919_);
  or (_35380_, _35379_, _35378_);
  and (_35381_, _35380_, _06251_);
  and (_35383_, _35381_, _35377_);
  and (_35384_, _14804_, _07919_);
  or (_35385_, _35384_, _35339_);
  and (_35386_, _35385_, _05972_);
  or (_35387_, _35386_, _06215_);
  or (_35388_, _35387_, _35383_);
  and (_35389_, _07919_, _08980_);
  or (_35390_, _35389_, _35339_);
  or (_35391_, _35390_, _06216_);
  and (_35392_, _35391_, _35388_);
  or (_35394_, _35392_, _06004_);
  and (_35395_, _35394_, _35336_);
  or (_35396_, _35395_, _06398_);
  and (_35397_, _14697_, _07919_);
  or (_35398_, _35397_, _35339_);
  or (_35399_, _35398_, _09025_);
  and (_35400_, _35399_, _09030_);
  and (_35401_, _35400_, _35396_);
  and (_35402_, _11250_, _07919_);
  or (_35403_, _35402_, _35339_);
  and (_35405_, _35403_, _06524_);
  or (_35406_, _35405_, _35401_);
  and (_35407_, _35406_, _07219_);
  or (_35408_, _35339_, _08424_);
  and (_35409_, _35390_, _06426_);
  and (_35410_, _35409_, _35408_);
  or (_35411_, _35410_, _35407_);
  and (_35412_, _35411_, _12729_);
  and (_35413_, _35346_, _06532_);
  and (_35414_, _35413_, _35408_);
  and (_35416_, _07854_, _06013_);
  or (_35417_, _35416_, _06437_);
  or (_35418_, _35417_, _35414_);
  or (_35419_, _35418_, _35412_);
  and (_35420_, _14694_, _07919_);
  or (_35421_, _35420_, _35339_);
  or (_35422_, _35421_, _07229_);
  and (_35423_, _35422_, _35419_);
  or (_35424_, _35423_, _06535_);
  nor (_35425_, _11249_, _13879_);
  or (_35427_, _35425_, _35339_);
  or (_35428_, _35427_, _07231_);
  and (_35429_, _35428_, _12782_);
  and (_35430_, _35429_, _35424_);
  and (_35431_, _15085_, _06543_);
  or (_35432_, _35431_, _06011_);
  or (_35433_, _35432_, _35430_);
  nand (_35434_, _15085_, _06011_);
  and (_35435_, _35434_, _06291_);
  and (_35436_, _35435_, _35433_);
  and (_35438_, _15085_, _06290_);
  or (_35439_, _35438_, _06559_);
  or (_35440_, _35439_, _35436_);
  or (_35441_, _35343_, _07240_);
  and (_35442_, _35441_, _07252_);
  and (_35443_, _35442_, _35440_);
  nor (_35444_, _15085_, _07252_);
  or (_35445_, _35444_, _06566_);
  or (_35446_, _35445_, _35443_);
  and (_35447_, _14873_, _08256_);
  or (_35449_, _35339_, _06570_);
  or (_35450_, _35449_, _35447_);
  and (_35451_, _35450_, _01320_);
  and (_35452_, _35451_, _35446_);
  or (_35453_, _35452_, _35335_);
  and (_43061_, _35453_, _42355_);
  nor (_35454_, _01320_, _06353_);
  or (_35455_, _07857_, _07252_);
  nand (_35456_, _15089_, _06004_);
  and (_35457_, _08256_, _09421_);
  nor (_35458_, _07919_, _06353_);
  or (_35459_, _35458_, _09486_);
  or (_35460_, _35459_, _35457_);
  and (_35461_, _35460_, _13787_);
  and (_35462_, _14900_, _08256_);
  or (_35463_, _35462_, _35458_);
  or (_35464_, _35463_, _06286_);
  and (_35465_, _07919_, \oc8051_golden_model_1.ACC [3]);
  or (_35466_, _35465_, _35458_);
  or (_35467_, _35466_, _07144_);
  or (_35469_, _07143_, \oc8051_golden_model_1.SP [3]);
  and (_35470_, _35469_, _07858_);
  and (_35471_, _35470_, _35467_);
  and (_35472_, _07857_, _07152_);
  or (_35473_, _35472_, _06285_);
  or (_35474_, _35473_, _35471_);
  and (_35475_, _35474_, _05949_);
  and (_35476_, _35475_, _35464_);
  nor (_35477_, _15089_, _05949_);
  or (_35478_, _35477_, _06354_);
  or (_35480_, _35478_, _35476_);
  nand (_35481_, _08647_, _06354_);
  and (_35482_, _35481_, _35480_);
  or (_35483_, _35482_, _06345_);
  or (_35484_, _35466_, _06346_);
  and (_35485_, _35484_, _06778_);
  and (_35486_, _35485_, _35483_);
  or (_35487_, _07630_, _35255_);
  or (_35488_, _35487_, _35486_);
  or (_35489_, _07857_, _07459_);
  and (_35491_, _35489_, _06260_);
  and (_35492_, _35491_, _35488_);
  or (_35493_, _35492_, _35461_);
  or (_35494_, _35458_, _06258_);
  and (_35495_, _09247_, _07919_);
  or (_35496_, _35495_, _35494_);
  and (_35497_, _35496_, _06251_);
  and (_35498_, _35497_, _35493_);
  and (_35499_, _14998_, _07919_);
  or (_35500_, _35499_, _35458_);
  and (_35502_, _35500_, _05972_);
  or (_35503_, _35502_, _06215_);
  or (_35504_, _35503_, _35498_);
  and (_35505_, _07919_, _08809_);
  or (_35506_, _35505_, _35458_);
  or (_35507_, _35506_, _06216_);
  and (_35508_, _35507_, _35504_);
  or (_35509_, _35508_, _06004_);
  and (_35510_, _35509_, _35456_);
  or (_35511_, _35510_, _06398_);
  and (_35513_, _14893_, _07919_);
  or (_35514_, _35513_, _35458_);
  or (_35515_, _35514_, _09025_);
  and (_35516_, _35515_, _09030_);
  and (_35517_, _35516_, _35511_);
  and (_35518_, _12529_, _07919_);
  or (_35519_, _35518_, _35458_);
  and (_35520_, _35519_, _06524_);
  or (_35521_, _35520_, _35517_);
  and (_35522_, _35521_, _07219_);
  or (_35524_, _35458_, _08280_);
  and (_35525_, _35506_, _06426_);
  and (_35526_, _35525_, _35524_);
  or (_35527_, _35526_, _35522_);
  and (_35528_, _35527_, _12729_);
  and (_35529_, _35466_, _06532_);
  and (_35530_, _35529_, _35524_);
  and (_35531_, _07857_, _06013_);
  or (_35532_, _35531_, _06437_);
  or (_35533_, _35532_, _35530_);
  or (_35535_, _35533_, _35528_);
  and (_35536_, _14890_, _08256_);
  or (_35537_, _35458_, _07229_);
  or (_35538_, _35537_, _35536_);
  and (_35539_, _35538_, _35535_);
  or (_35540_, _35539_, _06535_);
  nor (_35541_, _11247_, _13879_);
  or (_35542_, _35541_, _35458_);
  or (_35543_, _35542_, _07231_);
  and (_35544_, _35543_, _12782_);
  and (_35546_, _35544_, _35540_);
  nor (_35547_, _08644_, _06353_);
  or (_35548_, _35547_, _08645_);
  and (_35549_, _35548_, _06543_);
  or (_35550_, _35549_, _06011_);
  or (_35551_, _35550_, _35546_);
  nand (_35552_, _15089_, _06011_);
  and (_35553_, _35552_, _35551_);
  or (_35554_, _35553_, _06290_);
  or (_35555_, _35548_, _06291_);
  and (_35557_, _35555_, _07240_);
  and (_35558_, _35557_, _35554_);
  and (_35559_, _35463_, _06559_);
  or (_35560_, _35559_, _07678_);
  or (_35561_, _35560_, _35558_);
  and (_35562_, _35561_, _35455_);
  or (_35563_, _35562_, _06566_);
  and (_35564_, _15068_, _08256_);
  or (_35565_, _35458_, _06570_);
  or (_35566_, _35565_, _35564_);
  and (_35568_, _35566_, _01320_);
  and (_35569_, _35568_, _35563_);
  or (_35570_, _35569_, _35454_);
  and (_43063_, _35570_, _42355_);
  nor (_35571_, _07585_, \oc8051_golden_model_1.SP [4]);
  nor (_35572_, _35571_, _13776_);
  or (_35573_, _35572_, _09057_);
  and (_35574_, _09420_, _08256_);
  nor (_35575_, _07919_, _13811_);
  or (_35576_, _35575_, _09486_);
  or (_35578_, _35576_, _35574_);
  and (_35579_, _35578_, _13787_);
  and (_35580_, _15133_, _08256_);
  or (_35581_, _35580_, _35575_);
  or (_35582_, _35581_, _06286_);
  and (_35583_, _07919_, \oc8051_golden_model_1.ACC [4]);
  or (_35584_, _35583_, _35575_);
  or (_35585_, _35584_, _07144_);
  or (_35586_, _07143_, \oc8051_golden_model_1.SP [4]);
  and (_35587_, _35586_, _07858_);
  and (_35589_, _35587_, _35585_);
  and (_35590_, _35572_, _07152_);
  or (_35591_, _35590_, _06285_);
  or (_35592_, _35591_, _35589_);
  and (_35593_, _35592_, _05949_);
  and (_35594_, _35593_, _35582_);
  and (_35595_, _35572_, _07460_);
  or (_35596_, _35595_, _06354_);
  or (_35597_, _35596_, _35594_);
  and (_35598_, _13812_, _06766_);
  nor (_35600_, _08646_, _13811_);
  nor (_35601_, _35600_, _35598_);
  nand (_35602_, _35601_, _06354_);
  and (_35603_, _35602_, _35597_);
  or (_35604_, _35603_, _06345_);
  or (_35605_, _35584_, _06346_);
  and (_35606_, _35605_, _06778_);
  and (_35607_, _35606_, _35604_);
  and (_35608_, _07586_, \oc8051_golden_model_1.SP [4]);
  nor (_35609_, _07586_, \oc8051_golden_model_1.SP [4]);
  nor (_35611_, _35609_, _35608_);
  nand (_35612_, _35611_, _06276_);
  nand (_35613_, _35612_, _07459_);
  or (_35614_, _35613_, _35607_);
  or (_35615_, _35572_, _07459_);
  and (_35616_, _35615_, _06260_);
  and (_35617_, _35616_, _35614_);
  or (_35618_, _35617_, _35579_);
  or (_35619_, _35575_, _06258_);
  and (_35620_, _09437_, _07919_);
  or (_35622_, _35620_, _35619_);
  and (_35623_, _35622_, _06251_);
  and (_35624_, _35623_, _35618_);
  and (_35625_, _15226_, _07919_);
  or (_35626_, _35625_, _35575_);
  and (_35627_, _35626_, _05972_);
  or (_35628_, _35627_, _06215_);
  or (_35629_, _35628_, _35624_);
  and (_35630_, _08919_, _07919_);
  or (_35631_, _35630_, _35575_);
  or (_35633_, _35631_, _06216_);
  and (_35634_, _35633_, _35629_);
  or (_35635_, _35634_, _06004_);
  or (_35636_, _35572_, _13852_);
  and (_35637_, _35636_, _35635_);
  or (_35638_, _35637_, _06398_);
  and (_35639_, _15114_, _07919_);
  or (_35640_, _35639_, _35575_);
  or (_35641_, _35640_, _09025_);
  and (_35642_, _35641_, _09030_);
  and (_35644_, _35642_, _35638_);
  and (_35645_, _11245_, _07919_);
  or (_35646_, _35645_, _35575_);
  and (_35647_, _35646_, _06524_);
  or (_35648_, _35647_, _35644_);
  and (_35649_, _35648_, _07219_);
  or (_35650_, _35575_, _08528_);
  and (_35651_, _35631_, _06426_);
  and (_35652_, _35651_, _35650_);
  or (_35653_, _35652_, _35649_);
  and (_35655_, _35653_, _12729_);
  and (_35656_, _35584_, _06532_);
  and (_35657_, _35656_, _35650_);
  and (_35658_, _35572_, _06013_);
  or (_35659_, _35658_, _06437_);
  or (_35660_, _35659_, _35657_);
  or (_35661_, _35660_, _35655_);
  and (_35662_, _15111_, _07919_);
  or (_35663_, _35662_, _35575_);
  or (_35664_, _35663_, _07229_);
  and (_35666_, _35664_, _35661_);
  or (_35667_, _35666_, _06535_);
  nor (_35668_, _11244_, _13879_);
  or (_35669_, _35668_, _35575_);
  or (_35670_, _35669_, _07231_);
  and (_35671_, _35670_, _12782_);
  and (_35672_, _35671_, _35667_);
  nor (_35673_, _08645_, _13811_);
  or (_35674_, _35673_, _13812_);
  and (_35675_, _35674_, _06543_);
  or (_35677_, _35675_, _06011_);
  or (_35678_, _35677_, _35672_);
  and (_35679_, _35678_, _35573_);
  or (_35680_, _35679_, _06290_);
  or (_35681_, _35674_, _06291_);
  and (_35682_, _35681_, _07240_);
  and (_35683_, _35682_, _35680_);
  and (_35684_, _35581_, _06559_);
  or (_35685_, _35684_, _07678_);
  or (_35686_, _35685_, _35683_);
  or (_35688_, _35572_, _07252_);
  and (_35689_, _35688_, _06570_);
  and (_35690_, _35689_, _35686_);
  and (_35691_, _15296_, _08256_);
  or (_35692_, _35691_, _35575_);
  and (_35693_, _35692_, _06566_);
  or (_35694_, _35693_, _01324_);
  or (_35695_, _35694_, _35690_);
  or (_35696_, _01320_, \oc8051_golden_model_1.SP [4]);
  and (_35697_, _35696_, _42355_);
  and (_43064_, _35697_, _35695_);
  nor (_35699_, _01320_, _13810_);
  nor (_35700_, _13776_, \oc8051_golden_model_1.SP [5]);
  nor (_35701_, _35700_, _13777_);
  or (_35702_, _35701_, _07252_);
  and (_35703_, _09419_, _08256_);
  nor (_35704_, _07919_, _13810_);
  or (_35705_, _35704_, _09486_);
  or (_35706_, _35705_, _35703_);
  and (_35707_, _35706_, _13787_);
  and (_35709_, _15330_, _08256_);
  or (_35710_, _35709_, _35704_);
  or (_35711_, _35710_, _06286_);
  and (_35712_, _07919_, \oc8051_golden_model_1.ACC [5]);
  or (_35713_, _35712_, _35704_);
  or (_35714_, _35713_, _07144_);
  or (_35715_, _07143_, \oc8051_golden_model_1.SP [5]);
  and (_35716_, _35715_, _07858_);
  and (_35717_, _35716_, _35714_);
  and (_35718_, _35701_, _07152_);
  or (_35720_, _35718_, _06285_);
  or (_35721_, _35720_, _35717_);
  and (_35722_, _35721_, _05949_);
  and (_35723_, _35722_, _35711_);
  and (_35724_, _35701_, _07460_);
  or (_35725_, _35724_, _06354_);
  or (_35726_, _35725_, _35723_);
  and (_35727_, _13813_, _06766_);
  nor (_35728_, _35598_, _13810_);
  nor (_35729_, _35728_, _35727_);
  nand (_35731_, _35729_, _06354_);
  and (_35732_, _35731_, _35726_);
  or (_35733_, _35732_, _06345_);
  or (_35734_, _35713_, _06346_);
  and (_35735_, _35734_, _06778_);
  and (_35736_, _35735_, _35733_);
  nor (_35737_, _35608_, \oc8051_golden_model_1.SP [5]);
  nor (_35738_, _35737_, _13825_);
  nand (_35739_, _35738_, _06276_);
  nand (_35740_, _35739_, _07459_);
  or (_35742_, _35740_, _35736_);
  or (_35743_, _35701_, _07459_);
  and (_35744_, _35743_, _06260_);
  and (_35745_, _35744_, _35742_);
  or (_35746_, _35745_, _35707_);
  or (_35747_, _35704_, _06258_);
  and (_35748_, _09436_, _07919_);
  or (_35749_, _35748_, _35747_);
  and (_35750_, _35749_, _06251_);
  and (_35751_, _35750_, _35746_);
  and (_35753_, _15421_, _07919_);
  or (_35754_, _35753_, _35704_);
  and (_35755_, _35754_, _05972_);
  or (_35756_, _35755_, _06215_);
  or (_35757_, _35756_, _35751_);
  and (_35758_, _08913_, _07919_);
  or (_35759_, _35758_, _35704_);
  or (_35760_, _35759_, _06216_);
  and (_35761_, _35760_, _35757_);
  or (_35762_, _35761_, _06004_);
  or (_35764_, _35701_, _13852_);
  and (_35765_, _35764_, _35762_);
  or (_35766_, _35765_, _06398_);
  and (_35767_, _15313_, _07919_);
  or (_35768_, _35767_, _35704_);
  or (_35769_, _35768_, _09025_);
  and (_35770_, _35769_, _09030_);
  and (_35771_, _35770_, _35766_);
  and (_35772_, _12536_, _07919_);
  or (_35773_, _35772_, _35704_);
  and (_35775_, _35773_, _06524_);
  or (_35776_, _35775_, _35771_);
  and (_35777_, _35776_, _07219_);
  or (_35778_, _35704_, _08231_);
  and (_35779_, _35759_, _06426_);
  and (_35780_, _35779_, _35778_);
  or (_35781_, _35780_, _35777_);
  and (_35782_, _35781_, _12729_);
  and (_35783_, _35713_, _06532_);
  and (_35784_, _35783_, _35778_);
  and (_35786_, _35701_, _06013_);
  or (_35787_, _35786_, _06437_);
  or (_35788_, _35787_, _35784_);
  or (_35789_, _35788_, _35782_);
  and (_35790_, _15310_, _07919_);
  or (_35791_, _35790_, _35704_);
  or (_35792_, _35791_, _07229_);
  and (_35793_, _35792_, _35789_);
  or (_35794_, _35793_, _06535_);
  nor (_35795_, _11241_, _13879_);
  or (_35797_, _35795_, _35704_);
  or (_35798_, _35797_, _07231_);
  and (_35799_, _35798_, _12782_);
  and (_35800_, _35799_, _35794_);
  nor (_35801_, _13812_, _13810_);
  or (_35802_, _35801_, _13813_);
  and (_35803_, _35802_, _06543_);
  or (_35804_, _35803_, _06011_);
  or (_35805_, _35804_, _35800_);
  or (_35806_, _35701_, _09057_);
  and (_35808_, _35806_, _35805_);
  or (_35809_, _35808_, _06290_);
  or (_35810_, _35802_, _06291_);
  and (_35811_, _35810_, _07240_);
  and (_35812_, _35811_, _35809_);
  and (_35813_, _35710_, _06559_);
  or (_35814_, _35813_, _07678_);
  or (_35815_, _35814_, _35812_);
  and (_35816_, _35815_, _35702_);
  or (_35817_, _35816_, _06566_);
  and (_35819_, _15493_, _08256_);
  or (_35820_, _35704_, _06570_);
  or (_35821_, _35820_, _35819_);
  and (_35822_, _35821_, _01320_);
  and (_35823_, _35822_, _35817_);
  or (_35824_, _35823_, _35699_);
  and (_43065_, _35824_, _42355_);
  nor (_35825_, _01320_, _13809_);
  nor (_35826_, _07919_, _13809_);
  and (_35827_, _15521_, _08256_);
  or (_35829_, _35827_, _35826_);
  or (_35830_, _35829_, _06286_);
  and (_35831_, _07919_, \oc8051_golden_model_1.ACC [6]);
  or (_35832_, _35831_, _35826_);
  or (_35833_, _35832_, _07144_);
  or (_35834_, _07143_, \oc8051_golden_model_1.SP [6]);
  and (_35835_, _35834_, _07858_);
  and (_35836_, _35835_, _35833_);
  nor (_35837_, _13777_, \oc8051_golden_model_1.SP [6]);
  nor (_35838_, _35837_, _13778_);
  and (_35840_, _35838_, _07152_);
  or (_35841_, _35840_, _06285_);
  or (_35842_, _35841_, _35836_);
  and (_35843_, _35842_, _05949_);
  and (_35844_, _35843_, _35830_);
  and (_35845_, _35838_, _07460_);
  or (_35846_, _35845_, _06354_);
  or (_35847_, _35846_, _35844_);
  nor (_35848_, _35727_, _13809_);
  nor (_35849_, _35848_, _13815_);
  nand (_35851_, _35849_, _06354_);
  and (_35852_, _35851_, _35847_);
  or (_35853_, _35852_, _06345_);
  or (_35854_, _35832_, _06346_);
  and (_35855_, _35854_, _06778_);
  and (_35856_, _35855_, _35853_);
  nor (_35857_, _13825_, \oc8051_golden_model_1.SP [6]);
  nor (_35858_, _35857_, _13826_);
  and (_35859_, _35858_, _06276_);
  or (_35860_, _35859_, _35856_);
  and (_35862_, _35860_, _07459_);
  and (_35863_, _35838_, _35255_);
  or (_35864_, _35863_, _06259_);
  or (_35865_, _35864_, _35862_);
  and (_35866_, _09418_, _08256_);
  or (_35867_, _35826_, _06260_);
  or (_35868_, _35867_, _35866_);
  and (_35869_, _35868_, _35865_);
  or (_35870_, _35869_, _09486_);
  and (_35871_, _09435_, _07919_);
  or (_35873_, _35826_, _06258_);
  or (_35874_, _35873_, _35871_);
  and (_35875_, _35874_, _06251_);
  and (_35876_, _35875_, _35870_);
  and (_35877_, _15623_, _08256_);
  or (_35878_, _35877_, _35826_);
  and (_35879_, _35878_, _05972_);
  or (_35880_, _35879_, _06215_);
  or (_35881_, _35880_, _35876_);
  and (_35882_, _08845_, _07919_);
  or (_35884_, _35882_, _35826_);
  or (_35885_, _35884_, _06216_);
  and (_35886_, _35885_, _35881_);
  or (_35887_, _35886_, _06004_);
  or (_35888_, _35838_, _13852_);
  and (_35889_, _35888_, _35887_);
  or (_35890_, _35889_, _06398_);
  and (_35891_, _15517_, _07919_);
  or (_35892_, _35891_, _35826_);
  or (_35893_, _35892_, _09025_);
  and (_35895_, _35893_, _09030_);
  and (_35896_, _35895_, _35890_);
  and (_35897_, _11239_, _07919_);
  or (_35898_, _35897_, _35826_);
  and (_35899_, _35898_, _06524_);
  or (_35900_, _35899_, _35896_);
  and (_35901_, _35900_, _07219_);
  or (_35902_, _35826_, _08128_);
  and (_35903_, _35884_, _06426_);
  and (_35904_, _35903_, _35902_);
  or (_35906_, _35904_, _35901_);
  and (_35907_, _35906_, _12729_);
  and (_35908_, _35832_, _06532_);
  and (_35909_, _35908_, _35902_);
  and (_35910_, _35838_, _06013_);
  or (_35911_, _35910_, _06437_);
  or (_35912_, _35911_, _35909_);
  or (_35913_, _35912_, _35907_);
  and (_35914_, _15514_, _07919_);
  or (_35915_, _35914_, _35826_);
  or (_35917_, _35915_, _07229_);
  and (_35918_, _35917_, _35913_);
  or (_35919_, _35918_, _06535_);
  nor (_35920_, _11238_, _13879_);
  or (_35921_, _35920_, _35826_);
  or (_35922_, _35921_, _07231_);
  and (_35923_, _35922_, _12782_);
  and (_35924_, _35923_, _35919_);
  nor (_35925_, _13813_, _13809_);
  or (_35926_, _35925_, _13814_);
  and (_35928_, _35926_, _06543_);
  or (_35929_, _35928_, _06011_);
  or (_35930_, _35929_, _35924_);
  or (_35931_, _35838_, _09057_);
  and (_35932_, _35931_, _06291_);
  and (_35933_, _35932_, _35930_);
  and (_35934_, _35926_, _06290_);
  or (_35935_, _35934_, _06559_);
  or (_35936_, _35935_, _35933_);
  or (_35937_, _35829_, _07240_);
  and (_35939_, _35937_, _07252_);
  and (_35940_, _35939_, _35936_);
  and (_35941_, _35838_, _07678_);
  or (_35942_, _35941_, _06566_);
  or (_35943_, _35942_, _35940_);
  and (_35944_, _15695_, _08256_);
  or (_35945_, _35826_, _06570_);
  or (_35946_, _35945_, _35944_);
  and (_35947_, _35946_, _01320_);
  and (_35948_, _35947_, _35943_);
  or (_35950_, _35948_, _35825_);
  and (_43066_, _35950_, _42355_);
  not (_35951_, \oc8051_golden_model_1.SBUF [0]);
  nor (_35952_, _01320_, _35951_);
  nand (_35953_, _11254_, _07894_);
  nor (_35954_, _07894_, _35951_);
  nor (_35955_, _35954_, _07217_);
  nand (_35956_, _35955_, _35953_);
  nor (_35957_, _08374_, _13908_);
  or (_35958_, _35957_, _35954_);
  or (_35960_, _35958_, _06286_);
  and (_35961_, _07894_, \oc8051_golden_model_1.ACC [0]);
  or (_35962_, _35961_, _35954_);
  and (_35963_, _35962_, _07143_);
  nor (_35964_, _07143_, _35951_);
  or (_35965_, _35964_, _06285_);
  or (_35966_, _35965_, _35963_);
  and (_35967_, _35966_, _07169_);
  and (_35968_, _35967_, _35960_);
  and (_35969_, _07894_, _07135_);
  or (_35971_, _35969_, _35954_);
  and (_35972_, _35971_, _06354_);
  or (_35973_, _35972_, _35968_);
  and (_35974_, _35973_, _06346_);
  and (_35975_, _35962_, _06345_);
  or (_35976_, _35975_, _06259_);
  or (_35977_, _35976_, _35974_);
  or (_35978_, _35971_, _06260_);
  and (_35979_, _35978_, _35977_);
  or (_35980_, _35979_, _09486_);
  and (_35982_, _09384_, _07894_);
  or (_35983_, _35954_, _06258_);
  or (_35984_, _35983_, _35982_);
  and (_35985_, _35984_, _35980_);
  or (_35986_, _35985_, _05972_);
  and (_35987_, _14413_, _07894_);
  or (_35988_, _35954_, _06251_);
  or (_35989_, _35988_, _35987_);
  and (_35990_, _35989_, _06216_);
  and (_35991_, _35990_, _35986_);
  and (_35993_, _07894_, _08929_);
  or (_35994_, _35993_, _35954_);
  and (_35995_, _35994_, _06215_);
  or (_35996_, _35995_, _06398_);
  or (_35997_, _35996_, _35991_);
  and (_35998_, _14311_, _07894_);
  or (_35999_, _35998_, _35954_);
  or (_36000_, _35999_, _09025_);
  and (_36001_, _36000_, _09030_);
  and (_36002_, _36001_, _35997_);
  nor (_36004_, _12532_, _13908_);
  or (_36005_, _36004_, _35954_);
  and (_36006_, _35953_, _06524_);
  and (_36007_, _36006_, _36005_);
  or (_36008_, _36007_, _36002_);
  and (_36009_, _36008_, _07219_);
  nand (_36010_, _35994_, _06426_);
  nor (_36011_, _36010_, _35957_);
  or (_36012_, _36011_, _06532_);
  or (_36013_, _36012_, _36009_);
  and (_36015_, _36013_, _35956_);
  or (_36016_, _36015_, _06437_);
  and (_36017_, _14307_, _07894_);
  or (_36018_, _35954_, _07229_);
  or (_36019_, _36018_, _36017_);
  and (_36020_, _36019_, _07231_);
  and (_36021_, _36020_, _36016_);
  and (_36022_, _36005_, _06535_);
  or (_36023_, _36022_, _19480_);
  or (_36024_, _36023_, _36021_);
  or (_36026_, _35958_, _06651_);
  and (_36027_, _36026_, _01320_);
  and (_36028_, _36027_, _36024_);
  or (_36029_, _36028_, _35952_);
  and (_43068_, _36029_, _42355_);
  or (_36030_, _07894_, \oc8051_golden_model_1.SBUF [1]);
  and (_36031_, _14520_, _07894_);
  not (_36032_, _36031_);
  and (_36033_, _36032_, _36030_);
  or (_36034_, _36033_, _06286_);
  and (_36036_, _13908_, \oc8051_golden_model_1.SBUF [1]);
  and (_36037_, _07894_, \oc8051_golden_model_1.ACC [1]);
  or (_36038_, _36037_, _36036_);
  and (_36039_, _36038_, _07143_);
  and (_36040_, _07144_, \oc8051_golden_model_1.SBUF [1]);
  or (_36041_, _36040_, _06285_);
  or (_36042_, _36041_, _36039_);
  and (_36043_, _36042_, _07169_);
  and (_36044_, _36043_, _36034_);
  and (_36045_, _07894_, _09422_);
  or (_36047_, _36045_, _36036_);
  and (_36048_, _36047_, _06354_);
  or (_36049_, _36048_, _36044_);
  and (_36050_, _36049_, _06346_);
  and (_36051_, _36038_, _06345_);
  or (_36052_, _36051_, _06259_);
  or (_36053_, _36052_, _36050_);
  or (_36054_, _36047_, _06260_);
  and (_36055_, _36054_, _36053_);
  or (_36056_, _36055_, _09486_);
  and (_36058_, _09339_, _07894_);
  or (_36059_, _36036_, _06258_);
  or (_36060_, _36059_, _36058_);
  and (_36061_, _36060_, _06251_);
  and (_36062_, _36061_, _36056_);
  or (_36063_, _14607_, _13908_);
  and (_36064_, _36030_, _05972_);
  and (_36065_, _36064_, _36063_);
  or (_36066_, _36065_, _36062_);
  and (_36067_, _36066_, _06399_);
  or (_36069_, _14505_, _13908_);
  and (_36070_, _36030_, _06398_);
  and (_36071_, _36070_, _36069_);
  nand (_36072_, _07894_, _07031_);
  and (_36073_, _36072_, _06215_);
  and (_36074_, _36073_, _36030_);
  or (_36075_, _36074_, _06524_);
  or (_36076_, _36075_, _36071_);
  or (_36077_, _36076_, _36067_);
  nor (_36078_, _11252_, _13908_);
  or (_36080_, _36078_, _36036_);
  nand (_36081_, _11251_, _07894_);
  and (_36082_, _36081_, _36080_);
  or (_36083_, _36082_, _09030_);
  and (_36084_, _36083_, _07219_);
  and (_36085_, _36084_, _36077_);
  or (_36086_, _14503_, _13908_);
  and (_36087_, _36030_, _06426_);
  and (_36088_, _36087_, _36086_);
  or (_36089_, _36088_, _06532_);
  or (_36091_, _36089_, _36085_);
  nor (_36092_, _36036_, _07217_);
  nand (_36093_, _36092_, _36081_);
  and (_36094_, _36093_, _07229_);
  and (_36095_, _36094_, _36091_);
  or (_36096_, _36072_, _08325_);
  and (_36097_, _36096_, _06437_);
  and (_36098_, _36097_, _36030_);
  or (_36099_, _36098_, _06535_);
  or (_36100_, _36099_, _36095_);
  or (_36102_, _36080_, _07231_);
  and (_36103_, _36102_, _36100_);
  or (_36104_, _36103_, _06559_);
  or (_36105_, _36033_, _07240_);
  and (_36106_, _36105_, _06570_);
  and (_36107_, _36106_, _36104_);
  or (_36108_, _36036_, _36031_);
  and (_36109_, _36108_, _06566_);
  or (_36110_, _36109_, _01324_);
  or (_36111_, _36110_, _36107_);
  or (_36113_, _01320_, \oc8051_golden_model_1.SBUF [1]);
  and (_36114_, _36113_, _42355_);
  and (_43069_, _36114_, _36111_);
  and (_36115_, _01324_, \oc8051_golden_model_1.SBUF [2]);
  and (_36116_, _13908_, \oc8051_golden_model_1.SBUF [2]);
  and (_36117_, _09293_, _07894_);
  or (_36118_, _36117_, _36116_);
  and (_36119_, _36118_, _09486_);
  and (_36120_, _14703_, _07894_);
  or (_36121_, _36120_, _36116_);
  or (_36123_, _36121_, _06286_);
  and (_36124_, _07894_, \oc8051_golden_model_1.ACC [2]);
  or (_36125_, _36124_, _36116_);
  and (_36126_, _36125_, _07143_);
  and (_36127_, _07144_, \oc8051_golden_model_1.SBUF [2]);
  or (_36128_, _36127_, _06285_);
  or (_36129_, _36128_, _36126_);
  and (_36130_, _36129_, _07169_);
  and (_36131_, _36130_, _36123_);
  and (_36132_, _07894_, _08662_);
  or (_36134_, _36132_, _36116_);
  and (_36135_, _36134_, _06354_);
  or (_36136_, _36135_, _36131_);
  and (_36137_, _36136_, _06346_);
  and (_36138_, _36125_, _06345_);
  or (_36139_, _36138_, _06259_);
  or (_36140_, _36139_, _36137_);
  or (_36141_, _36134_, _06260_);
  and (_36142_, _36141_, _06258_);
  and (_36143_, _36142_, _36140_);
  or (_36145_, _36143_, _05972_);
  or (_36146_, _36145_, _36119_);
  and (_36147_, _14804_, _07894_);
  or (_36148_, _36116_, _06251_);
  or (_36149_, _36148_, _36147_);
  and (_36150_, _36149_, _06216_);
  and (_36151_, _36150_, _36146_);
  and (_36152_, _07894_, _08980_);
  or (_36153_, _36152_, _36116_);
  and (_36154_, _36153_, _06215_);
  or (_36156_, _36154_, _06398_);
  or (_36157_, _36156_, _36151_);
  and (_36158_, _14697_, _07894_);
  or (_36159_, _36158_, _36116_);
  or (_36160_, _36159_, _09025_);
  and (_36161_, _36160_, _09030_);
  and (_36162_, _36161_, _36157_);
  and (_36163_, _11250_, _07894_);
  or (_36164_, _36163_, _36116_);
  and (_36165_, _36164_, _06524_);
  or (_36167_, _36165_, _36162_);
  and (_36168_, _36167_, _07219_);
  or (_36169_, _36116_, _08424_);
  and (_36170_, _36153_, _06426_);
  and (_36171_, _36170_, _36169_);
  or (_36172_, _36171_, _36168_);
  and (_36173_, _36172_, _07217_);
  and (_36174_, _36125_, _06532_);
  and (_36175_, _36174_, _36169_);
  or (_36176_, _36175_, _06437_);
  or (_36178_, _36176_, _36173_);
  and (_36179_, _14694_, _07894_);
  or (_36180_, _36116_, _07229_);
  or (_36181_, _36180_, _36179_);
  and (_36182_, _36181_, _07231_);
  and (_36183_, _36182_, _36178_);
  nor (_36184_, _11249_, _13908_);
  or (_36185_, _36184_, _36116_);
  and (_36186_, _36185_, _06535_);
  or (_36187_, _36186_, _36183_);
  and (_36189_, _36187_, _07240_);
  and (_36190_, _36121_, _06559_);
  or (_36191_, _36190_, _06566_);
  or (_36192_, _36191_, _36189_);
  and (_36193_, _14873_, _07894_);
  or (_36194_, _36116_, _06570_);
  or (_36195_, _36194_, _36193_);
  and (_36196_, _36195_, _01320_);
  and (_36197_, _36196_, _36192_);
  or (_36198_, _36197_, _36115_);
  and (_43070_, _36198_, _42355_);
  and (_36199_, _13908_, \oc8051_golden_model_1.SBUF [3]);
  and (_36200_, _14900_, _07894_);
  or (_36201_, _36200_, _36199_);
  or (_36202_, _36201_, _06286_);
  and (_36203_, _07894_, \oc8051_golden_model_1.ACC [3]);
  or (_36204_, _36203_, _36199_);
  and (_36205_, _36204_, _07143_);
  and (_36206_, _07144_, \oc8051_golden_model_1.SBUF [3]);
  or (_36207_, _36206_, _06285_);
  or (_36209_, _36207_, _36205_);
  and (_36210_, _36209_, _07169_);
  and (_36211_, _36210_, _36202_);
  and (_36212_, _07894_, _09421_);
  or (_36213_, _36212_, _36199_);
  and (_36214_, _36213_, _06354_);
  or (_36215_, _36214_, _36211_);
  and (_36216_, _36215_, _06346_);
  and (_36217_, _36204_, _06345_);
  or (_36218_, _36217_, _06259_);
  or (_36220_, _36218_, _36216_);
  or (_36221_, _36213_, _06260_);
  and (_36222_, _36221_, _36220_);
  or (_36223_, _36222_, _09486_);
  and (_36224_, _09247_, _07894_);
  or (_36225_, _36199_, _06258_);
  or (_36226_, _36225_, _36224_);
  and (_36227_, _36226_, _06251_);
  and (_36228_, _36227_, _36223_);
  and (_36229_, _14998_, _07894_);
  or (_36231_, _36229_, _36199_);
  and (_36232_, _36231_, _05972_);
  or (_36233_, _36232_, _10080_);
  or (_36234_, _36233_, _36228_);
  and (_36235_, _14893_, _07894_);
  or (_36236_, _36199_, _09025_);
  or (_36237_, _36236_, _36235_);
  and (_36238_, _07894_, _08809_);
  or (_36239_, _36238_, _36199_);
  or (_36240_, _36239_, _06216_);
  and (_36242_, _36240_, _09030_);
  and (_36243_, _36242_, _36237_);
  and (_36244_, _36243_, _36234_);
  and (_36245_, _12529_, _07894_);
  or (_36246_, _36245_, _36199_);
  and (_36247_, _36246_, _06524_);
  or (_36248_, _36247_, _36244_);
  and (_36249_, _36248_, _07219_);
  or (_36250_, _36199_, _08280_);
  and (_36251_, _36239_, _06426_);
  and (_36253_, _36251_, _36250_);
  or (_36254_, _36253_, _36249_);
  and (_36255_, _36254_, _07217_);
  and (_36256_, _36204_, _06532_);
  and (_36257_, _36256_, _36250_);
  or (_36258_, _36257_, _06437_);
  or (_36259_, _36258_, _36255_);
  and (_36260_, _14890_, _07894_);
  or (_36261_, _36199_, _07229_);
  or (_36262_, _36261_, _36260_);
  and (_36264_, _36262_, _07231_);
  and (_36265_, _36264_, _36259_);
  nor (_36266_, _11247_, _13908_);
  or (_36267_, _36266_, _36199_);
  and (_36268_, _36267_, _06535_);
  or (_36269_, _36268_, _06559_);
  or (_36270_, _36269_, _36265_);
  or (_36271_, _36201_, _07240_);
  and (_36272_, _36271_, _06570_);
  and (_36273_, _36272_, _36270_);
  and (_36275_, _15068_, _07894_);
  or (_36276_, _36275_, _36199_);
  and (_36277_, _36276_, _06566_);
  or (_36278_, _36277_, _01324_);
  or (_36279_, _36278_, _36273_);
  or (_36280_, _01320_, \oc8051_golden_model_1.SBUF [3]);
  and (_36281_, _36280_, _42355_);
  and (_43071_, _36281_, _36279_);
  and (_36282_, _13908_, \oc8051_golden_model_1.SBUF [4]);
  and (_36283_, _09420_, _07894_);
  or (_36285_, _36283_, _36282_);
  or (_36286_, _36285_, _06260_);
  and (_36287_, _15133_, _07894_);
  or (_36288_, _36287_, _36282_);
  or (_36289_, _36288_, _06286_);
  and (_36290_, _07894_, \oc8051_golden_model_1.ACC [4]);
  or (_36291_, _36290_, _36282_);
  and (_36292_, _36291_, _07143_);
  and (_36293_, _07144_, \oc8051_golden_model_1.SBUF [4]);
  or (_36294_, _36293_, _06285_);
  or (_36296_, _36294_, _36292_);
  and (_36297_, _36296_, _07169_);
  and (_36298_, _36297_, _36289_);
  and (_36299_, _36285_, _06354_);
  or (_36300_, _36299_, _36298_);
  and (_36301_, _36300_, _06346_);
  and (_36302_, _36291_, _06345_);
  or (_36303_, _36302_, _06259_);
  or (_36304_, _36303_, _36301_);
  and (_36305_, _36304_, _06258_);
  and (_36307_, _36305_, _36286_);
  and (_36308_, _09437_, _07894_);
  or (_36309_, _36308_, _36282_);
  and (_36310_, _36309_, _09486_);
  or (_36311_, _36310_, _05972_);
  or (_36312_, _36311_, _36307_);
  and (_36313_, _15226_, _07894_);
  or (_36314_, _36282_, _06251_);
  or (_36315_, _36314_, _36313_);
  and (_36316_, _36315_, _06216_);
  and (_36318_, _36316_, _36312_);
  and (_36319_, _08919_, _07894_);
  or (_36320_, _36319_, _36282_);
  and (_36321_, _36320_, _06215_);
  or (_36322_, _36321_, _06398_);
  or (_36323_, _36322_, _36318_);
  and (_36324_, _15114_, _07894_);
  or (_36325_, _36324_, _36282_);
  or (_36326_, _36325_, _09025_);
  and (_36327_, _36326_, _09030_);
  and (_36329_, _36327_, _36323_);
  and (_36330_, _11245_, _07894_);
  or (_36331_, _36330_, _36282_);
  and (_36332_, _36331_, _06524_);
  or (_36333_, _36332_, _36329_);
  and (_36334_, _36333_, _07219_);
  or (_36335_, _36282_, _08528_);
  and (_36336_, _36320_, _06426_);
  and (_36337_, _36336_, _36335_);
  or (_36338_, _36337_, _36334_);
  and (_36340_, _36338_, _07217_);
  and (_36341_, _36291_, _06532_);
  and (_36342_, _36341_, _36335_);
  or (_36343_, _36342_, _06437_);
  or (_36344_, _36343_, _36340_);
  and (_36345_, _15111_, _07894_);
  or (_36346_, _36282_, _07229_);
  or (_36347_, _36346_, _36345_);
  and (_36348_, _36347_, _07231_);
  and (_36349_, _36348_, _36344_);
  nor (_36351_, _11244_, _13908_);
  or (_36352_, _36351_, _36282_);
  and (_36353_, _36352_, _06535_);
  or (_36354_, _36353_, _06559_);
  or (_36355_, _36354_, _36349_);
  or (_36356_, _36288_, _07240_);
  and (_36357_, _36356_, _06570_);
  and (_36358_, _36357_, _36355_);
  and (_36359_, _15296_, _07894_);
  or (_36360_, _36359_, _36282_);
  and (_36362_, _36360_, _06566_);
  or (_36363_, _36362_, _01324_);
  or (_36364_, _36363_, _36358_);
  or (_36365_, _01320_, \oc8051_golden_model_1.SBUF [4]);
  and (_36366_, _36365_, _42355_);
  and (_43072_, _36366_, _36364_);
  and (_36367_, _13908_, \oc8051_golden_model_1.SBUF [5]);
  and (_36368_, _15330_, _07894_);
  or (_36369_, _36368_, _36367_);
  or (_36370_, _36369_, _06286_);
  and (_36372_, _07894_, \oc8051_golden_model_1.ACC [5]);
  or (_36373_, _36372_, _36367_);
  and (_36374_, _36373_, _07143_);
  and (_36375_, _07144_, \oc8051_golden_model_1.SBUF [5]);
  or (_36376_, _36375_, _06285_);
  or (_36377_, _36376_, _36374_);
  and (_36378_, _36377_, _07169_);
  and (_36379_, _36378_, _36370_);
  and (_36380_, _09419_, _07894_);
  or (_36381_, _36380_, _36367_);
  and (_36383_, _36381_, _06354_);
  or (_36384_, _36383_, _36379_);
  and (_36385_, _36384_, _06346_);
  and (_36386_, _36373_, _06345_);
  or (_36387_, _36386_, _06259_);
  or (_36388_, _36387_, _36385_);
  or (_36389_, _36381_, _06260_);
  and (_36390_, _36389_, _36388_);
  or (_36391_, _36390_, _09486_);
  and (_36392_, _09436_, _07894_);
  or (_36394_, _36367_, _06258_);
  or (_36395_, _36394_, _36392_);
  and (_36396_, _36395_, _06251_);
  and (_36397_, _36396_, _36391_);
  and (_36398_, _15421_, _07894_);
  or (_36399_, _36398_, _36367_);
  and (_36400_, _36399_, _05972_);
  or (_36401_, _36400_, _10080_);
  or (_36402_, _36401_, _36397_);
  and (_36403_, _15313_, _07894_);
  or (_36405_, _36367_, _09025_);
  or (_36406_, _36405_, _36403_);
  and (_36407_, _08913_, _07894_);
  or (_36408_, _36407_, _36367_);
  or (_36409_, _36408_, _06216_);
  and (_36410_, _36409_, _09030_);
  and (_36411_, _36410_, _36406_);
  and (_36412_, _36411_, _36402_);
  and (_36413_, _12536_, _07894_);
  or (_36414_, _36413_, _36367_);
  and (_36416_, _36414_, _06524_);
  or (_36417_, _36416_, _36412_);
  and (_36418_, _36417_, _07219_);
  or (_36419_, _36367_, _08231_);
  and (_36420_, _36408_, _06426_);
  and (_36421_, _36420_, _36419_);
  or (_36422_, _36421_, _36418_);
  and (_36423_, _36422_, _07217_);
  and (_36424_, _36373_, _06532_);
  and (_36425_, _36424_, _36419_);
  or (_36427_, _36425_, _06437_);
  or (_36428_, _36427_, _36423_);
  and (_36429_, _15310_, _07894_);
  or (_36430_, _36367_, _07229_);
  or (_36431_, _36430_, _36429_);
  and (_36432_, _36431_, _07231_);
  and (_36433_, _36432_, _36428_);
  nor (_36434_, _11241_, _13908_);
  or (_36435_, _36434_, _36367_);
  and (_36436_, _36435_, _06535_);
  or (_36438_, _36436_, _06559_);
  or (_36439_, _36438_, _36433_);
  or (_36440_, _36369_, _07240_);
  and (_36441_, _36440_, _06570_);
  and (_36442_, _36441_, _36439_);
  and (_36443_, _15493_, _07894_);
  or (_36444_, _36443_, _36367_);
  and (_36445_, _36444_, _06566_);
  or (_36446_, _36445_, _01324_);
  or (_36447_, _36446_, _36442_);
  or (_36449_, _01320_, \oc8051_golden_model_1.SBUF [5]);
  and (_36450_, _36449_, _42355_);
  and (_43073_, _36450_, _36447_);
  and (_36451_, _13908_, \oc8051_golden_model_1.SBUF [6]);
  and (_36452_, _15521_, _07894_);
  or (_36453_, _36452_, _36451_);
  or (_36454_, _36453_, _06286_);
  and (_36455_, _07894_, \oc8051_golden_model_1.ACC [6]);
  or (_36456_, _36455_, _36451_);
  and (_36457_, _36456_, _07143_);
  and (_36459_, _07144_, \oc8051_golden_model_1.SBUF [6]);
  or (_36460_, _36459_, _06285_);
  or (_36461_, _36460_, _36457_);
  and (_36462_, _36461_, _07169_);
  and (_36463_, _36462_, _36454_);
  and (_36464_, _09418_, _07894_);
  or (_36465_, _36464_, _36451_);
  and (_36466_, _36465_, _06354_);
  or (_36467_, _36466_, _36463_);
  and (_36468_, _36467_, _06346_);
  and (_36470_, _36456_, _06345_);
  or (_36471_, _36470_, _06259_);
  or (_36472_, _36471_, _36468_);
  or (_36473_, _36465_, _06260_);
  and (_36474_, _36473_, _36472_);
  or (_36475_, _36474_, _09486_);
  and (_36476_, _09435_, _07894_);
  or (_36477_, _36451_, _06258_);
  or (_36478_, _36477_, _36476_);
  and (_36479_, _36478_, _06251_);
  and (_36481_, _36479_, _36475_);
  and (_36482_, _15623_, _07894_);
  or (_36483_, _36482_, _36451_);
  and (_36484_, _36483_, _05972_);
  or (_36485_, _36484_, _10080_);
  or (_36486_, _36485_, _36481_);
  and (_36487_, _15517_, _07894_);
  or (_36488_, _36451_, _09025_);
  or (_36489_, _36488_, _36487_);
  and (_36490_, _08845_, _07894_);
  or (_36492_, _36490_, _36451_);
  or (_36493_, _36492_, _06216_);
  and (_36494_, _36493_, _09030_);
  and (_36495_, _36494_, _36489_);
  and (_36496_, _36495_, _36486_);
  and (_36497_, _11239_, _07894_);
  or (_36498_, _36497_, _36451_);
  and (_36499_, _36498_, _06524_);
  or (_36500_, _36499_, _36496_);
  and (_36501_, _36500_, _07219_);
  or (_36503_, _36451_, _08128_);
  and (_36504_, _36492_, _06426_);
  and (_36505_, _36504_, _36503_);
  or (_36506_, _36505_, _36501_);
  and (_36507_, _36506_, _07217_);
  and (_36508_, _36456_, _06532_);
  and (_36509_, _36508_, _36503_);
  or (_36510_, _36509_, _06437_);
  or (_36511_, _36510_, _36507_);
  and (_36512_, _15514_, _07894_);
  or (_36514_, _36451_, _07229_);
  or (_36515_, _36514_, _36512_);
  and (_36516_, _36515_, _07231_);
  and (_36517_, _36516_, _36511_);
  nor (_36518_, _11238_, _13908_);
  or (_36519_, _36518_, _36451_);
  and (_36520_, _36519_, _06535_);
  or (_36521_, _36520_, _06559_);
  or (_36522_, _36521_, _36517_);
  or (_36523_, _36453_, _07240_);
  and (_36525_, _36523_, _06570_);
  and (_36526_, _36525_, _36522_);
  and (_36527_, _15695_, _07894_);
  or (_36528_, _36527_, _36451_);
  and (_36529_, _36528_, _06566_);
  or (_36530_, _36529_, _01324_);
  or (_36531_, _36530_, _36526_);
  or (_36532_, _01320_, \oc8051_golden_model_1.SBUF [6]);
  and (_36533_, _36532_, _42355_);
  and (_43074_, _36533_, _36531_);
  not (_36535_, \oc8051_golden_model_1.PSW [0]);
  nor (_36536_, _01320_, _36535_);
  nand (_36537_, _11254_, _07926_);
  nor (_36538_, _07926_, _36535_);
  nor (_36539_, _36538_, _07217_);
  nand (_36540_, _36539_, _36537_);
  and (_36541_, _07926_, _07135_);
  or (_36542_, _36541_, _36538_);
  or (_36543_, _36542_, _06260_);
  nor (_36544_, _08374_, _14234_);
  or (_36546_, _36544_, _36538_);
  or (_36547_, _36546_, _06286_);
  and (_36548_, _07926_, \oc8051_golden_model_1.ACC [0]);
  or (_36549_, _36548_, _36538_);
  and (_36550_, _36549_, _07143_);
  nor (_36551_, _07143_, _36535_);
  or (_36552_, _36551_, _06285_);
  or (_36553_, _36552_, _36550_);
  and (_36554_, _36553_, _06282_);
  and (_36555_, _36554_, _36547_);
  nor (_36557_, _08592_, _36535_);
  and (_36558_, _14326_, _08592_);
  or (_36559_, _36558_, _36557_);
  and (_36560_, _36559_, _06281_);
  or (_36561_, _36560_, _36555_);
  and (_36562_, _36561_, _07169_);
  and (_36563_, _36542_, _06354_);
  or (_36564_, _36563_, _06345_);
  or (_36565_, _36564_, _36562_);
  or (_36566_, _36549_, _06346_);
  and (_36568_, _36566_, _06278_);
  and (_36569_, _36568_, _36565_);
  and (_36570_, _36538_, _06277_);
  or (_36571_, _36570_, _06270_);
  or (_36572_, _36571_, _36569_);
  or (_36573_, _36546_, _06271_);
  and (_36574_, _36573_, _06267_);
  and (_36575_, _36574_, _36572_);
  and (_36576_, _14358_, _08592_);
  or (_36577_, _36576_, _36557_);
  and (_36579_, _36577_, _06266_);
  or (_36580_, _36579_, _06259_);
  or (_36581_, _36580_, _36575_);
  and (_36582_, _36581_, _36543_);
  or (_36583_, _36582_, _09486_);
  and (_36584_, _09384_, _07926_);
  or (_36585_, _36538_, _06258_);
  or (_36586_, _36585_, _36584_);
  and (_36587_, _36586_, _06251_);
  and (_36588_, _36587_, _36583_);
  and (_36590_, _14413_, _07926_);
  or (_36591_, _36590_, _36538_);
  and (_36592_, _36591_, _05972_);
  or (_36593_, _36592_, _36588_);
  or (_36594_, _36593_, _10080_);
  and (_36595_, _14311_, _07926_);
  or (_36596_, _36538_, _09025_);
  or (_36597_, _36596_, _36595_);
  and (_36598_, _07926_, _08929_);
  or (_36599_, _36598_, _36538_);
  or (_36601_, _36599_, _06216_);
  and (_36602_, _36601_, _09030_);
  and (_36603_, _36602_, _36597_);
  and (_36604_, _36603_, _36594_);
  nor (_36605_, _12532_, _14234_);
  or (_36606_, _36605_, _36538_);
  and (_36607_, _36537_, _06524_);
  and (_36608_, _36607_, _36606_);
  or (_36609_, _36608_, _36604_);
  and (_36610_, _36609_, _07219_);
  nand (_36612_, _36599_, _06426_);
  nor (_36613_, _36612_, _36544_);
  or (_36614_, _36613_, _06532_);
  or (_36615_, _36614_, _36610_);
  and (_36616_, _36615_, _36540_);
  or (_36617_, _36616_, _06437_);
  and (_36618_, _14307_, _07926_);
  or (_36619_, _36538_, _07229_);
  or (_36620_, _36619_, _36618_);
  and (_36621_, _36620_, _07231_);
  and (_36623_, _36621_, _36617_);
  and (_36624_, _36606_, _06535_);
  or (_36625_, _36624_, _06559_);
  or (_36626_, _36625_, _36623_);
  or (_36627_, _36546_, _07240_);
  and (_36628_, _36627_, _36626_);
  or (_36629_, _36628_, _05932_);
  or (_36630_, _36538_, _05933_);
  and (_36631_, _36630_, _36629_);
  or (_36632_, _36631_, _06566_);
  or (_36634_, _36546_, _06570_);
  and (_36635_, _36634_, _01320_);
  and (_36636_, _36635_, _36632_);
  or (_36637_, _36636_, _36536_);
  and (_43075_, _36637_, _42355_);
  not (_36638_, \oc8051_golden_model_1.PSW [1]);
  nor (_36639_, _01320_, _36638_);
  nor (_36640_, _07926_, _36638_);
  and (_36641_, _07926_, _09422_);
  or (_36642_, _36641_, _36640_);
  or (_36644_, _36642_, _07169_);
  or (_36645_, _07926_, \oc8051_golden_model_1.PSW [1]);
  and (_36646_, _14520_, _07926_);
  not (_36647_, _36646_);
  and (_36648_, _36647_, _36645_);
  or (_36649_, _36648_, _06286_);
  and (_36650_, _07926_, \oc8051_golden_model_1.ACC [1]);
  or (_36651_, _36650_, _36640_);
  and (_36652_, _36651_, _07143_);
  nor (_36653_, _07143_, _36638_);
  or (_36655_, _36653_, _06285_);
  or (_36656_, _36655_, _36652_);
  and (_36657_, _36656_, _06282_);
  and (_36658_, _36657_, _36649_);
  nor (_36659_, _08592_, _36638_);
  and (_36660_, _14508_, _08592_);
  or (_36661_, _36660_, _36659_);
  and (_36662_, _36661_, _06281_);
  or (_36663_, _36662_, _06354_);
  or (_36664_, _36663_, _36658_);
  and (_36666_, _36664_, _36644_);
  or (_36667_, _36666_, _06345_);
  or (_36668_, _36651_, _06346_);
  and (_36669_, _36668_, _06278_);
  and (_36670_, _36669_, _36667_);
  and (_36671_, _14511_, _08592_);
  or (_36672_, _36671_, _36659_);
  and (_36673_, _36672_, _06277_);
  or (_36674_, _36673_, _06270_);
  or (_36675_, _36674_, _36670_);
  and (_36677_, _36660_, _14507_);
  or (_36678_, _36659_, _06271_);
  or (_36679_, _36678_, _36677_);
  and (_36680_, _36679_, _06267_);
  and (_36681_, _36680_, _36675_);
  or (_36682_, _36659_, _14551_);
  and (_36683_, _36682_, _06266_);
  and (_36684_, _36683_, _36661_);
  or (_36685_, _36684_, _06259_);
  or (_36686_, _36685_, _36681_);
  or (_36688_, _36642_, _06260_);
  and (_36689_, _36688_, _36686_);
  or (_36690_, _36689_, _09486_);
  and (_36691_, _09339_, _07926_);
  or (_36692_, _36640_, _06258_);
  or (_36693_, _36692_, _36691_);
  and (_36694_, _36693_, _06251_);
  and (_36695_, _36694_, _36690_);
  and (_36696_, _14607_, _07926_);
  or (_36697_, _36696_, _36640_);
  and (_36699_, _36697_, _05972_);
  or (_36700_, _36699_, _36695_);
  and (_36701_, _36700_, _06399_);
  or (_36702_, _14505_, _14234_);
  and (_36703_, _36645_, _06398_);
  and (_36704_, _36703_, _36702_);
  nand (_36705_, _07926_, _07031_);
  and (_36706_, _36705_, _06215_);
  and (_36707_, _36706_, _36645_);
  or (_36708_, _36707_, _06524_);
  or (_36710_, _36708_, _36704_);
  or (_36711_, _36710_, _36701_);
  nor (_36712_, _11252_, _14234_);
  or (_36713_, _36712_, _36640_);
  nand (_36714_, _11251_, _07926_);
  and (_36715_, _36714_, _36713_);
  or (_36716_, _36715_, _09030_);
  and (_36717_, _36716_, _07219_);
  and (_36718_, _36717_, _36711_);
  or (_36719_, _14503_, _14234_);
  and (_36721_, _36645_, _06426_);
  and (_36722_, _36721_, _36719_);
  or (_36723_, _36722_, _06532_);
  or (_36724_, _36723_, _36718_);
  nor (_36725_, _36640_, _07217_);
  nand (_36726_, _36725_, _36714_);
  and (_36727_, _36726_, _07229_);
  and (_36728_, _36727_, _36724_);
  or (_36729_, _36705_, _08325_);
  and (_36730_, _36645_, _06437_);
  and (_36732_, _36730_, _36729_);
  or (_36733_, _36732_, _06535_);
  or (_36734_, _36733_, _36728_);
  or (_36735_, _36713_, _07231_);
  and (_36736_, _36735_, _36734_);
  or (_36737_, _36736_, _06559_);
  or (_36738_, _36648_, _07240_);
  and (_36739_, _36738_, _05933_);
  and (_36740_, _36739_, _36737_);
  and (_36741_, _36672_, _05932_);
  or (_36743_, _36741_, _06566_);
  or (_36744_, _36743_, _36740_);
  or (_36745_, _36640_, _06570_);
  or (_36746_, _36745_, _36646_);
  and (_36747_, _36746_, _01320_);
  and (_36748_, _36747_, _36744_);
  or (_36749_, _36748_, _36639_);
  and (_43076_, _36749_, _42355_);
  and (_36750_, _01324_, \oc8051_golden_model_1.PSW [2]);
  not (_36751_, _10924_);
  nor (_36753_, _10562_, _36751_);
  nor (_36754_, _10563_, \oc8051_golden_model_1.ACC [7]);
  nor (_36755_, _36754_, _36753_);
  not (_36756_, _36755_);
  nor (_36757_, _36756_, _14244_);
  nor (_36758_, _36757_, _36753_);
  and (_36759_, _36758_, _11078_);
  and (_36760_, _36753_, _11075_);
  or (_36761_, _36760_, _36759_);
  and (_36762_, _36761_, _11026_);
  and (_36764_, _14234_, \oc8051_golden_model_1.PSW [2]);
  and (_36765_, _14804_, _07926_);
  or (_36766_, _36765_, _36764_);
  and (_36767_, _36766_, _05972_);
  and (_36768_, _07926_, _08662_);
  or (_36769_, _36768_, _36764_);
  or (_36770_, _36769_, _06260_);
  and (_36771_, _36769_, _06354_);
  not (_36772_, _08592_);
  and (_36773_, _36772_, \oc8051_golden_model_1.PSW [2]);
  and (_36775_, _14716_, _08592_);
  or (_36776_, _36775_, _36773_);
  or (_36777_, _36776_, _06282_);
  and (_36778_, _14703_, _07926_);
  or (_36779_, _36778_, _36764_);
  and (_36780_, _36779_, _06285_);
  and (_36781_, _07144_, \oc8051_golden_model_1.PSW [2]);
  and (_36782_, _07926_, \oc8051_golden_model_1.ACC [2]);
  or (_36783_, _36782_, _36764_);
  and (_36784_, _36783_, _07143_);
  or (_36786_, _36784_, _36781_);
  and (_36787_, _36786_, _06286_);
  or (_36788_, _36787_, _06281_);
  or (_36789_, _36788_, _36780_);
  and (_36790_, _36789_, _36777_);
  and (_36791_, _36790_, _07169_);
  or (_36792_, _36791_, _36771_);
  or (_36793_, _36792_, _06345_);
  or (_36794_, _36783_, _06346_);
  and (_36795_, _36794_, _06278_);
  and (_36797_, _36795_, _36793_);
  and (_36798_, _14699_, _08592_);
  or (_36799_, _36798_, _36773_);
  and (_36800_, _36799_, _06277_);
  or (_36801_, _36800_, _36797_);
  and (_36802_, _36801_, _06271_);
  or (_36803_, _36773_, _14731_);
  and (_36804_, _36776_, _06270_);
  and (_36805_, _36804_, _36803_);
  or (_36806_, _36805_, _36802_);
  and (_36808_, _36806_, _10059_);
  or (_36809_, _16450_, _10061_);
  or (_36810_, _36809_, _16568_);
  or (_36811_, _36810_, _16677_);
  or (_36812_, _36811_, _16795_);
  or (_36813_, _36812_, _16912_);
  or (_36814_, _36813_, _17028_);
  or (_36815_, _36814_, _17145_);
  and (_36816_, _36815_, _09520_);
  or (_36817_, _36816_, _17293_);
  or (_36819_, _36817_, _36808_);
  or (_36820_, _10728_, _08023_);
  nor (_36821_, _36820_, _08737_);
  and (_36822_, _36820_, _08737_);
  or (_36823_, _36822_, _36821_);
  and (_36824_, _36823_, _14161_);
  nor (_36825_, _36823_, _14161_);
  nor (_36826_, _36825_, _36824_);
  not (_36827_, _36826_);
  nor (_36828_, _36827_, _10793_);
  and (_36830_, _36827_, _10793_);
  or (_36831_, _36830_, _36828_);
  or (_36832_, _36831_, _10724_);
  and (_36833_, _36832_, _36819_);
  and (_36834_, _36833_, _10555_);
  nor (_36835_, _36755_, _10568_);
  nor (_36836_, _14009_, _10564_);
  or (_36837_, _36836_, _36835_);
  or (_36838_, _36837_, _10617_);
  nand (_36839_, _36837_, _10617_);
  and (_36841_, _36839_, _36838_);
  and (_36842_, _36841_, _10727_);
  or (_36843_, _36842_, _36834_);
  and (_36844_, _36843_, _06386_);
  nor (_36845_, _10494_, _14278_);
  nor (_36846_, _10495_, \oc8051_golden_model_1.ACC [7]);
  nor (_36847_, _36846_, _36845_);
  not (_36848_, _36847_);
  or (_36849_, _36848_, _14175_);
  nand (_36850_, _36848_, _14175_);
  and (_36852_, _36850_, _36849_);
  and (_36853_, _36852_, _10552_);
  nor (_36854_, _36852_, _10552_);
  or (_36855_, _36854_, _36853_);
  and (_36856_, _36855_, _06380_);
  or (_36857_, _36856_, _10486_);
  or (_36858_, _36857_, _36844_);
  not (_36859_, _10933_);
  nor (_36860_, _10804_, _36859_);
  not (_36861_, _36860_);
  nor (_36863_, _10804_, _06294_);
  or (_36864_, _36863_, \oc8051_golden_model_1.ACC [7]);
  and (_36865_, _36864_, _36861_);
  nor (_36866_, _36865_, _14185_);
  and (_36867_, _36865_, _14185_);
  nor (_36868_, _36867_, _36866_);
  and (_36869_, _36868_, _10862_);
  nor (_36870_, _36868_, _10862_);
  or (_36871_, _36870_, _36869_);
  or (_36872_, _36871_, _10487_);
  and (_36874_, _36872_, _06267_);
  and (_36875_, _36874_, _36858_);
  and (_36876_, _14749_, _08592_);
  or (_36877_, _36876_, _36773_);
  and (_36878_, _36877_, _06266_);
  or (_36879_, _36878_, _06259_);
  or (_36880_, _36879_, _36875_);
  and (_36881_, _36880_, _36770_);
  or (_36882_, _36881_, _09486_);
  and (_36883_, _09293_, _07926_);
  or (_36885_, _36764_, _06258_);
  or (_36886_, _36885_, _36883_);
  and (_36887_, _36886_, _06251_);
  and (_36888_, _36887_, _36882_);
  or (_36889_, _36888_, _36767_);
  and (_36890_, _36889_, _09481_);
  nor (_36891_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_36892_, _36891_, _10104_);
  nand (_36893_, _36892_, _09480_);
  nand (_36894_, _36893_, _06399_);
  or (_36896_, _36894_, _36890_);
  and (_36897_, _14697_, _07926_);
  or (_36898_, _36764_, _09025_);
  or (_36899_, _36898_, _36897_);
  and (_36900_, _07926_, _08980_);
  or (_36901_, _36900_, _36764_);
  or (_36902_, _36901_, _06216_);
  and (_36903_, _36902_, _09030_);
  and (_36904_, _36903_, _36899_);
  and (_36905_, _36904_, _36896_);
  and (_36907_, _11250_, _07926_);
  or (_36908_, _36907_, _36764_);
  and (_36909_, _36908_, _06524_);
  or (_36910_, _36909_, _36905_);
  and (_36911_, _36910_, _07219_);
  or (_36912_, _36764_, _08424_);
  and (_36913_, _36901_, _06426_);
  and (_36914_, _36913_, _36912_);
  or (_36915_, _36914_, _36911_);
  and (_36916_, _36915_, _07217_);
  and (_36918_, _36783_, _06532_);
  and (_36919_, _36918_, _36912_);
  or (_36920_, _36919_, _06437_);
  or (_36921_, _36920_, _36916_);
  and (_36922_, _14694_, _07926_);
  or (_36923_, _36922_, _36764_);
  or (_36924_, _36923_, _07229_);
  and (_36925_, _36924_, _07231_);
  and (_36926_, _36925_, _36921_);
  nor (_36927_, _11249_, _14234_);
  or (_36929_, _36927_, _36764_);
  and (_36930_, _36929_, _06535_);
  or (_36931_, _36930_, _11024_);
  or (_36932_, _36931_, _36926_);
  nor (_36933_, _36823_, _13992_);
  nor (_36934_, _36933_, _36821_);
  and (_36935_, _36934_, _11051_);
  and (_36936_, _36821_, _11048_);
  or (_36937_, _36936_, _11023_);
  or (_36938_, _36937_, _36935_);
  and (_36939_, _36938_, _17490_);
  and (_36940_, _36939_, _36932_);
  or (_36941_, _36940_, _36762_);
  and (_36942_, _36941_, _17717_);
  and (_36943_, _36761_, _06892_);
  or (_36944_, _36943_, _06522_);
  or (_36945_, _36944_, _36942_);
  nor (_36946_, _36848_, _14249_);
  nor (_36947_, _36946_, _36845_);
  and (_36948_, _36947_, _11107_);
  and (_36950_, _36845_, _11104_);
  or (_36951_, _36950_, _36948_);
  or (_36952_, _36951_, _06523_);
  and (_36953_, _36952_, _11083_);
  and (_36954_, _36953_, _36945_);
  not (_36955_, _36865_);
  or (_36956_, _36955_, _14255_);
  and (_36957_, _36861_, _11135_);
  and (_36958_, _36957_, _36956_);
  and (_36959_, _36860_, _11132_);
  or (_36961_, _36959_, _36958_);
  nand (_36962_, _36961_, _11082_);
  nand (_36963_, _36962_, _11185_);
  or (_36964_, _36963_, _36954_);
  and (_36965_, _11178_, _10903_);
  not (_36966_, _10902_);
  nor (_36967_, _11178_, _36966_);
  or (_36968_, _36967_, _36965_);
  or (_36969_, _36968_, _11185_);
  and (_36970_, _36969_, _11190_);
  and (_36972_, _36970_, _36964_);
  or (_36973_, _11229_, _10923_);
  nand (_36974_, _11229_, _36751_);
  and (_36975_, _36974_, _11191_);
  and (_36976_, _36975_, _36973_);
  or (_36977_, _36976_, _36972_);
  and (_36978_, _36977_, _12978_);
  or (_36979_, _11267_, _09041_);
  and (_36980_, _14280_, _36979_);
  and (_36981_, _11306_, _36859_);
  or (_36983_, _36981_, _14285_);
  nand (_36984_, _36983_, _07240_);
  or (_36985_, _36984_, _36980_);
  or (_36986_, _36985_, _36978_);
  or (_36987_, _36779_, _07240_);
  and (_36988_, _36987_, _05933_);
  and (_36989_, _36988_, _36986_);
  and (_36990_, _36799_, _05932_);
  or (_36991_, _36990_, _06566_);
  or (_36992_, _36991_, _36989_);
  and (_36994_, _14873_, _07926_);
  or (_36995_, _36764_, _06570_);
  or (_36996_, _36995_, _36994_);
  and (_36997_, _36996_, _01320_);
  and (_36998_, _36997_, _36992_);
  or (_36999_, _36998_, _36750_);
  and (_43077_, _36999_, _42355_);
  nor (_37000_, _01320_, _06362_);
  nor (_37001_, _07926_, _06362_);
  and (_37002_, _14900_, _07926_);
  or (_37004_, _37002_, _37001_);
  or (_37005_, _37004_, _06286_);
  and (_37006_, _07926_, \oc8051_golden_model_1.ACC [3]);
  or (_37007_, _37006_, _37001_);
  and (_37008_, _37007_, _07143_);
  nor (_37009_, _07143_, _06362_);
  or (_37010_, _37009_, _06285_);
  or (_37011_, _37010_, _37008_);
  and (_37012_, _37011_, _06282_);
  and (_37013_, _37012_, _37005_);
  nor (_37015_, _08592_, _06362_);
  and (_37016_, _14897_, _08592_);
  or (_37017_, _37016_, _37015_);
  and (_37018_, _37017_, _06281_);
  or (_37019_, _37018_, _06354_);
  or (_37020_, _37019_, _37013_);
  and (_37021_, _07926_, _09421_);
  or (_37022_, _37021_, _37001_);
  or (_37023_, _37022_, _07169_);
  and (_37024_, _37023_, _37020_);
  or (_37026_, _37024_, _06345_);
  or (_37027_, _37007_, _06346_);
  and (_37028_, _37027_, _06278_);
  and (_37029_, _37028_, _37026_);
  and (_37030_, _14895_, _08592_);
  or (_37031_, _37030_, _37015_);
  and (_37032_, _37031_, _06277_);
  or (_37033_, _37032_, _06270_);
  or (_37034_, _37033_, _37029_);
  or (_37035_, _37015_, _14926_);
  and (_37037_, _37035_, _37017_);
  or (_37038_, _37037_, _06271_);
  and (_37039_, _37038_, _06267_);
  and (_37040_, _37039_, _37034_);
  and (_37041_, _14943_, _08592_);
  or (_37042_, _37041_, _37015_);
  and (_37043_, _37042_, _06266_);
  or (_37044_, _37043_, _06259_);
  or (_37045_, _37044_, _37040_);
  or (_37046_, _37022_, _06260_);
  and (_37048_, _37046_, _06258_);
  and (_37049_, _37048_, _37045_);
  and (_37050_, _09247_, _07926_);
  or (_37051_, _37050_, _37001_);
  and (_37052_, _37051_, _09486_);
  or (_37053_, _37052_, _05972_);
  or (_37054_, _37053_, _37049_);
  and (_37055_, _14998_, _07926_);
  or (_37056_, _37001_, _06251_);
  or (_37057_, _37056_, _37055_);
  and (_37059_, _37057_, _06216_);
  and (_37060_, _37059_, _37054_);
  and (_37061_, _07926_, _08809_);
  or (_37062_, _37061_, _37001_);
  and (_37063_, _37062_, _06215_);
  or (_37064_, _37063_, _06398_);
  or (_37065_, _37064_, _37060_);
  and (_37066_, _14893_, _07926_);
  or (_37067_, _37066_, _37001_);
  or (_37068_, _37067_, _09025_);
  and (_37070_, _37068_, _09030_);
  and (_37071_, _37070_, _37065_);
  and (_37072_, _12529_, _07926_);
  or (_37073_, _37072_, _37001_);
  and (_37074_, _37073_, _06524_);
  or (_37075_, _37074_, _37071_);
  and (_37076_, _37075_, _07219_);
  or (_37077_, _37001_, _08280_);
  and (_37078_, _37062_, _06426_);
  and (_37079_, _37078_, _37077_);
  or (_37081_, _37079_, _37076_);
  and (_37082_, _37081_, _07217_);
  and (_37083_, _37007_, _06532_);
  and (_37084_, _37083_, _37077_);
  or (_37085_, _37084_, _06437_);
  or (_37086_, _37085_, _37082_);
  and (_37087_, _14890_, _07926_);
  or (_37088_, _37001_, _07229_);
  or (_37089_, _37088_, _37087_);
  and (_37090_, _37089_, _07231_);
  and (_37092_, _37090_, _37086_);
  nor (_37093_, _11247_, _14234_);
  or (_37094_, _37093_, _37001_);
  and (_37095_, _37094_, _06535_);
  or (_37096_, _37095_, _06559_);
  or (_37097_, _37096_, _37092_);
  or (_37098_, _37004_, _07240_);
  and (_37099_, _37098_, _05933_);
  and (_37100_, _37099_, _37097_);
  and (_37101_, _37031_, _05932_);
  or (_37103_, _37101_, _06566_);
  or (_37104_, _37103_, _37100_);
  and (_37105_, _15068_, _07926_);
  or (_37106_, _37001_, _06570_);
  or (_37107_, _37106_, _37105_);
  and (_37108_, _37107_, _01320_);
  and (_37109_, _37108_, _37104_);
  or (_37110_, _37109_, _37000_);
  and (_43078_, _37110_, _42355_);
  and (_37111_, _01324_, \oc8051_golden_model_1.PSW [4]);
  and (_37113_, _09437_, _07926_);
  and (_37114_, _14234_, \oc8051_golden_model_1.PSW [4]);
  or (_37115_, _37114_, _06258_);
  or (_37116_, _37115_, _37113_);
  and (_37117_, _09420_, _07926_);
  or (_37118_, _37117_, _37114_);
  or (_37119_, _37118_, _06260_);
  and (_37120_, _15133_, _07926_);
  or (_37121_, _37120_, _37114_);
  or (_37122_, _37121_, _06286_);
  and (_37124_, _07926_, \oc8051_golden_model_1.ACC [4]);
  or (_37125_, _37124_, _37114_);
  and (_37126_, _37125_, _07143_);
  and (_37127_, _07144_, \oc8051_golden_model_1.PSW [4]);
  or (_37128_, _37127_, _06285_);
  or (_37129_, _37128_, _37126_);
  and (_37130_, _37129_, _06282_);
  and (_37131_, _37130_, _37122_);
  and (_37132_, _36772_, \oc8051_golden_model_1.PSW [4]);
  and (_37133_, _15116_, _08592_);
  or (_37135_, _37133_, _37132_);
  and (_37136_, _37135_, _06281_);
  or (_37137_, _37136_, _06354_);
  or (_37138_, _37137_, _37131_);
  or (_37139_, _37118_, _07169_);
  and (_37140_, _37139_, _37138_);
  or (_37141_, _37140_, _06345_);
  or (_37142_, _37125_, _06346_);
  and (_37143_, _37142_, _06278_);
  and (_37144_, _37143_, _37141_);
  and (_37146_, _15145_, _08592_);
  or (_37147_, _37146_, _37132_);
  and (_37148_, _37147_, _06277_);
  or (_37149_, _37148_, _06270_);
  or (_37150_, _37149_, _37144_);
  or (_37151_, _37132_, _15152_);
  and (_37152_, _37151_, _37135_);
  or (_37153_, _37152_, _06271_);
  and (_37154_, _37153_, _06267_);
  and (_37155_, _37154_, _37150_);
  and (_37157_, _15170_, _08592_);
  or (_37158_, _37157_, _37132_);
  and (_37159_, _37158_, _06266_);
  or (_37160_, _37159_, _06259_);
  or (_37161_, _37160_, _37155_);
  and (_37162_, _37161_, _37119_);
  or (_37163_, _37162_, _09486_);
  and (_37164_, _37163_, _37116_);
  or (_37165_, _37164_, _05972_);
  and (_37166_, _15226_, _07926_);
  or (_37168_, _37114_, _06251_);
  or (_37169_, _37168_, _37166_);
  and (_37170_, _37169_, _06216_);
  and (_37171_, _37170_, _37165_);
  and (_37172_, _08919_, _07926_);
  or (_37173_, _37172_, _37114_);
  and (_37174_, _37173_, _06215_);
  or (_37175_, _37174_, _06398_);
  or (_37176_, _37175_, _37171_);
  and (_37177_, _15114_, _07926_);
  or (_37179_, _37177_, _37114_);
  or (_37180_, _37179_, _09025_);
  and (_37181_, _37180_, _09030_);
  and (_37182_, _37181_, _37176_);
  and (_37183_, _11245_, _07926_);
  or (_37184_, _37183_, _37114_);
  and (_37185_, _37184_, _06524_);
  or (_37186_, _37185_, _37182_);
  and (_37187_, _37186_, _07219_);
  or (_37188_, _37114_, _08528_);
  and (_37190_, _37173_, _06426_);
  and (_37191_, _37190_, _37188_);
  or (_37192_, _37191_, _37187_);
  and (_37193_, _37192_, _07217_);
  and (_37194_, _37125_, _06532_);
  and (_37195_, _37194_, _37188_);
  or (_37196_, _37195_, _06437_);
  or (_37197_, _37196_, _37193_);
  and (_37198_, _15111_, _07926_);
  or (_37199_, _37114_, _07229_);
  or (_37201_, _37199_, _37198_);
  and (_37202_, _37201_, _07231_);
  and (_37203_, _37202_, _37197_);
  nor (_37204_, _11244_, _14234_);
  or (_37205_, _37204_, _37114_);
  and (_37206_, _37205_, _06535_);
  or (_37207_, _37206_, _06559_);
  or (_37208_, _37207_, _37203_);
  or (_37209_, _37121_, _07240_);
  and (_37210_, _37209_, _05933_);
  and (_37212_, _37210_, _37208_);
  and (_37213_, _37147_, _05932_);
  or (_37214_, _37213_, _06566_);
  or (_37215_, _37214_, _37212_);
  and (_37216_, _15296_, _07926_);
  or (_37217_, _37114_, _06570_);
  or (_37218_, _37217_, _37216_);
  and (_37219_, _37218_, _01320_);
  and (_37220_, _37219_, _37215_);
  or (_37221_, _37220_, _37111_);
  and (_43079_, _37221_, _42355_);
  and (_37223_, _01324_, \oc8051_golden_model_1.PSW [5]);
  and (_37224_, _14234_, \oc8051_golden_model_1.PSW [5]);
  and (_37225_, _15330_, _07926_);
  or (_37226_, _37225_, _37224_);
  or (_37227_, _37226_, _06286_);
  and (_37228_, _07926_, \oc8051_golden_model_1.ACC [5]);
  or (_37229_, _37228_, _37224_);
  and (_37230_, _37229_, _07143_);
  and (_37231_, _07144_, \oc8051_golden_model_1.PSW [5]);
  or (_37233_, _37231_, _06285_);
  or (_37234_, _37233_, _37230_);
  and (_37235_, _37234_, _06282_);
  and (_37236_, _37235_, _37227_);
  and (_37237_, _36772_, \oc8051_golden_model_1.PSW [5]);
  and (_37238_, _15315_, _08592_);
  or (_37239_, _37238_, _37237_);
  and (_37240_, _37239_, _06281_);
  or (_37241_, _37240_, _06354_);
  or (_37242_, _37241_, _37236_);
  and (_37244_, _09419_, _07926_);
  or (_37245_, _37244_, _37224_);
  or (_37246_, _37245_, _07169_);
  and (_37247_, _37246_, _37242_);
  or (_37248_, _37247_, _06345_);
  or (_37249_, _37229_, _06346_);
  and (_37250_, _37249_, _06278_);
  and (_37251_, _37250_, _37248_);
  and (_37252_, _15342_, _08592_);
  or (_37253_, _37252_, _37237_);
  and (_37255_, _37253_, _06277_);
  or (_37256_, _37255_, _06270_);
  or (_37257_, _37256_, _37251_);
  or (_37258_, _37237_, _15349_);
  and (_37259_, _37258_, _37239_);
  or (_37260_, _37259_, _06271_);
  and (_37261_, _37260_, _06267_);
  and (_37262_, _37261_, _37257_);
  or (_37263_, _37237_, _15365_);
  and (_37264_, _37263_, _06266_);
  and (_37266_, _37264_, _37239_);
  or (_37267_, _37266_, _06259_);
  or (_37268_, _37267_, _37262_);
  or (_37269_, _37245_, _06260_);
  and (_37270_, _37269_, _37268_);
  or (_37271_, _37270_, _09486_);
  and (_37272_, _09436_, _07926_);
  or (_37273_, _37224_, _06258_);
  or (_37274_, _37273_, _37272_);
  and (_37275_, _37274_, _06251_);
  and (_37277_, _37275_, _37271_);
  and (_37278_, _15421_, _07926_);
  or (_37279_, _37278_, _37224_);
  and (_37280_, _37279_, _05972_);
  or (_37281_, _37280_, _10080_);
  or (_37282_, _37281_, _37277_);
  and (_37283_, _15313_, _07926_);
  or (_37284_, _37224_, _09025_);
  or (_37285_, _37284_, _37283_);
  and (_37286_, _08913_, _07926_);
  or (_37288_, _37286_, _37224_);
  or (_37289_, _37288_, _06216_);
  and (_37290_, _37289_, _09030_);
  and (_37291_, _37290_, _37285_);
  and (_37292_, _37291_, _37282_);
  and (_37293_, _12536_, _07926_);
  or (_37294_, _37293_, _37224_);
  and (_37295_, _37294_, _06524_);
  or (_37296_, _37295_, _37292_);
  and (_37297_, _37296_, _07219_);
  or (_37299_, _37224_, _08231_);
  and (_37300_, _37288_, _06426_);
  and (_37301_, _37300_, _37299_);
  or (_37302_, _37301_, _37297_);
  and (_37303_, _37302_, _07217_);
  and (_37304_, _37229_, _06532_);
  and (_37305_, _37304_, _37299_);
  or (_37306_, _37305_, _06437_);
  or (_37307_, _37306_, _37303_);
  and (_37308_, _15310_, _07926_);
  or (_37310_, _37224_, _07229_);
  or (_37311_, _37310_, _37308_);
  and (_37312_, _37311_, _07231_);
  and (_37313_, _37312_, _37307_);
  nor (_37314_, _11241_, _14234_);
  or (_37315_, _37314_, _37224_);
  and (_37316_, _37315_, _06535_);
  or (_37317_, _37316_, _06559_);
  or (_37318_, _37317_, _37313_);
  or (_37319_, _37226_, _07240_);
  and (_37321_, _37319_, _05933_);
  and (_37322_, _37321_, _37318_);
  and (_37323_, _37253_, _05932_);
  or (_37324_, _37323_, _06566_);
  or (_37325_, _37324_, _37322_);
  and (_37326_, _15493_, _07926_);
  or (_37327_, _37224_, _06570_);
  or (_37328_, _37327_, _37326_);
  and (_37329_, _37328_, _01320_);
  and (_37330_, _37329_, _37325_);
  or (_37332_, _37330_, _37223_);
  and (_43081_, _37332_, _42355_);
  nor (_37333_, _01320_, _18155_);
  or (_37334_, _11185_, _11171_);
  or (_37335_, _11027_, _10559_);
  or (_37336_, _37335_, _11069_);
  and (_37337_, _06407_, _06010_);
  and (_37338_, _06409_, _06010_);
  or (_37339_, _11042_, _10745_);
  and (_37340_, _37339_, _11017_);
  nor (_37342_, _07926_, _18155_);
  and (_37343_, _09418_, _07926_);
  or (_37344_, _37343_, _37342_);
  or (_37345_, _37344_, _06260_);
  nor (_37346_, _08592_, _18155_);
  and (_37347_, _15535_, _08592_);
  or (_37348_, _37347_, _37346_);
  or (_37349_, _37346_, _15551_);
  and (_37350_, _37349_, _37348_);
  or (_37351_, _37350_, _06271_);
  and (_37353_, _15521_, _07926_);
  or (_37354_, _37353_, _37342_);
  or (_37355_, _37354_, _06286_);
  and (_37356_, _07926_, \oc8051_golden_model_1.ACC [6]);
  or (_37357_, _37356_, _37342_);
  and (_37358_, _37357_, _07143_);
  nor (_37359_, _07143_, _18155_);
  or (_37360_, _37359_, _06285_);
  or (_37361_, _37360_, _37358_);
  and (_37362_, _37361_, _06282_);
  and (_37364_, _37362_, _37355_);
  and (_37365_, _37348_, _06281_);
  or (_37366_, _37365_, _06354_);
  or (_37367_, _37366_, _37364_);
  or (_37368_, _37344_, _07169_);
  and (_37369_, _37368_, _37367_);
  or (_37370_, _37369_, _06345_);
  or (_37371_, _37357_, _06346_);
  and (_37372_, _37371_, _06278_);
  and (_37373_, _37372_, _37370_);
  and (_37375_, _15544_, _08592_);
  or (_37376_, _37375_, _37346_);
  and (_37377_, _37376_, _06277_);
  or (_37378_, _37377_, _06270_);
  or (_37379_, _37378_, _37373_);
  and (_37380_, _37379_, _37351_);
  or (_37381_, _37380_, _17293_);
  or (_37382_, _10745_, _10724_);
  or (_37383_, _37382_, _10783_);
  and (_37384_, _37383_, _37381_);
  or (_37386_, _37384_, _10727_);
  or (_37387_, _10559_, _10555_);
  or (_37388_, _37387_, _10610_);
  and (_37389_, _37388_, _37386_);
  or (_37390_, _37389_, _12600_);
  or (_37391_, _10491_, _06386_);
  or (_37392_, _37391_, _10542_);
  or (_37393_, _10801_, _10487_);
  or (_37394_, _37393_, _10849_);
  and (_37395_, _37394_, _06267_);
  and (_37397_, _37395_, _37392_);
  and (_37398_, _37397_, _37390_);
  and (_37399_, _15568_, _08592_);
  or (_37400_, _37399_, _37346_);
  and (_37401_, _37400_, _06266_);
  or (_37402_, _37401_, _06259_);
  or (_37403_, _37402_, _37398_);
  and (_37404_, _37403_, _37345_);
  or (_37405_, _37404_, _09486_);
  and (_37406_, _09435_, _07926_);
  or (_37408_, _37342_, _06258_);
  or (_37409_, _37408_, _37406_);
  and (_37410_, _37409_, _06251_);
  and (_37411_, _37410_, _37405_);
  and (_37412_, _15623_, _07926_);
  or (_37413_, _37412_, _37342_);
  and (_37414_, _37413_, _05972_);
  or (_37415_, _37414_, _10080_);
  or (_37416_, _37415_, _37411_);
  and (_37417_, _15517_, _07926_);
  or (_37419_, _37342_, _09025_);
  or (_37420_, _37419_, _37417_);
  and (_37421_, _08845_, _07926_);
  or (_37422_, _37421_, _37342_);
  or (_37423_, _37422_, _06216_);
  and (_37424_, _37423_, _09030_);
  and (_37425_, _37424_, _37420_);
  and (_37426_, _37425_, _37416_);
  and (_37427_, _11239_, _07926_);
  or (_37428_, _37427_, _37342_);
  and (_37430_, _37428_, _06524_);
  or (_37431_, _37430_, _37426_);
  and (_37432_, _37431_, _07219_);
  or (_37433_, _37342_, _08128_);
  and (_37434_, _37422_, _06426_);
  and (_37435_, _37434_, _37433_);
  or (_37436_, _37435_, _37432_);
  and (_37437_, _37436_, _07217_);
  and (_37438_, _37357_, _06532_);
  and (_37439_, _37438_, _37433_);
  or (_37441_, _37439_, _06437_);
  or (_37442_, _37441_, _37437_);
  and (_37443_, _15514_, _07926_);
  or (_37444_, _37443_, _37342_);
  or (_37445_, _37444_, _07229_);
  and (_37446_, _37445_, _37442_);
  or (_37447_, _37446_, _06535_);
  nor (_37448_, _11238_, _14234_);
  or (_37449_, _37448_, _37342_);
  or (_37450_, _37449_, _07231_);
  and (_37452_, _37450_, _11018_);
  and (_37453_, _37452_, _37447_);
  nor (_37454_, _37453_, _37340_);
  nor (_37455_, _37454_, _37338_);
  and (_37456_, _37339_, _37338_);
  nor (_37457_, _37456_, _37455_);
  nor (_37458_, _37457_, _37337_);
  and (_37459_, _37339_, _37337_);
  or (_37460_, _37459_, _06887_);
  or (_37461_, _37460_, _37458_);
  or (_37463_, _37339_, _06888_);
  and (_37464_, _37463_, _11020_);
  and (_37465_, _37464_, _37461_);
  and (_37466_, _37339_, _11019_);
  or (_37467_, _37466_, _13990_);
  or (_37468_, _37467_, _37465_);
  and (_37469_, _37468_, _37336_);
  or (_37470_, _37469_, _06522_);
  or (_37471_, _10491_, _06523_);
  or (_37472_, _37471_, _11098_);
  and (_37474_, _37472_, _11083_);
  and (_37475_, _37474_, _37470_);
  or (_37476_, _11126_, _10801_);
  and (_37477_, _37476_, _11082_);
  or (_37478_, _37477_, _11184_);
  or (_37479_, _37478_, _37475_);
  and (_37480_, _37479_, _37334_);
  or (_37481_, _37480_, _11191_);
  or (_37482_, _11223_, _11190_);
  and (_37483_, _37482_, _06293_);
  and (_37485_, _37483_, _37481_);
  and (_37486_, _11261_, _06292_);
  or (_37487_, _37486_, _10474_);
  or (_37488_, _37487_, _37485_);
  or (_37489_, _11300_, _10475_);
  and (_37490_, _37489_, _37488_);
  or (_37491_, _37490_, _06559_);
  or (_37492_, _37354_, _07240_);
  and (_37493_, _37492_, _05933_);
  and (_37494_, _37493_, _37491_);
  and (_37496_, _37376_, _05932_);
  or (_37497_, _37496_, _06566_);
  or (_37498_, _37497_, _37494_);
  and (_37499_, _15695_, _07926_);
  or (_37500_, _37342_, _06570_);
  or (_37501_, _37500_, _37499_);
  and (_37502_, _37501_, _01320_);
  and (_37503_, _37502_, _37498_);
  or (_37504_, _37503_, _37333_);
  and (_43082_, _37504_, _42355_);
  or (_37506_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand (_37507_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_37508_, _37507_, _37506_);
  or (_37509_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nand (_37510_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_37511_, _37510_, _37509_);
  or (_37512_, _37511_, _37508_);
  or (_37513_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_37514_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_37515_, _37514_, _37513_);
  or (_37517_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_37518_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_37519_, _37518_, _37517_);
  or (_37520_, _37519_, _37515_);
  or (_37521_, _37520_, _37512_);
  nor (_37522_, _10198_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_37523_, _10198_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_37524_, _37523_, _37522_);
  nand (_37525_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_37526_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_37528_, _37526_, _37525_);
  or (_37529_, _37528_, _37524_);
  nand (_37530_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_37531_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_37532_, _37531_, _37530_);
  and (_37533_, _08737_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_37534_, _08737_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_37535_, _37534_, _37533_);
  or (_37536_, _37535_, _37532_);
  or (_37537_, _37536_, _37529_);
  or (_37539_, _37537_, _37521_);
  and (_37540_, inst_finished_r, op0_cnst);
  and (property_invalid_acc, _37540_, _37539_);
  and (_37541_, _05766_, op0_cnst);
  or (_00001_, _37541_, rst);
  buf (_00543_, _42358_);
  buf (_05080_, _42355_);
  buf (_05132_, _42355_);
  buf (_05183_, _42355_);
  buf (_05235_, _42355_);
  buf (_05287_, _42355_);
  buf (_05338_, _42355_);
  buf (_05390_, _42355_);
  buf (_05441_, _42355_);
  buf (_05493_, _42355_);
  buf (_05544_, _42355_);
  buf (_05596_, _42355_);
  buf (_05649_, _42355_);
  buf (_05702_, _42355_);
  buf (_05755_, _42355_);
  buf (_05808_, _42355_);
  buf (_05861_, _42355_);
  buf (_38484_, _38382_);
  buf (_38486_, _38384_);
  buf (_38499_, _38382_);
  buf (_38500_, _38384_);
  buf (_38813_, _38403_);
  buf (_38814_, _38404_);
  buf (_38815_, _38406_);
  buf (_38816_, _38407_);
  buf (_38817_, _38408_);
  buf (_38818_, _38409_);
  buf (_38819_, _38410_);
  buf (_38820_, _38412_);
  buf (_38821_, _38413_);
  buf (_38823_, _38414_);
  buf (_38824_, _38415_);
  buf (_38825_, _38416_);
  buf (_38826_, _38418_);
  buf (_38827_, _38419_);
  buf (_38878_, _38403_);
  buf (_38879_, _38404_);
  buf (_38880_, _38406_);
  buf (_38881_, _38407_);
  buf (_38882_, _38408_);
  buf (_38883_, _38409_);
  buf (_38884_, _38410_);
  buf (_38885_, _38412_);
  buf (_38886_, _38413_);
  buf (_38888_, _38414_);
  buf (_38889_, _38415_);
  buf (_38890_, _38416_);
  buf (_38891_, _38418_);
  buf (_38892_, _38419_);
  buf (_39424_, _39196_);
  buf (_39584_, _39196_);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _05084_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _05088_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _05092_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _05096_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _05100_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _05104_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _05108_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _05077_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _05080_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _05136_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _05140_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _05143_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _05147_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _05151_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _05155_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _05159_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _05129_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _05132_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _05600_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _05604_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _05608_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _05612_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _05616_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _05620_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _05624_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _05593_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _05596_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _05653_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _05657_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _05661_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _05665_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _05669_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _05673_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _05677_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _05646_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _05649_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _05706_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _05710_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _05714_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _05718_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _05722_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _05726_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _05730_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _05699_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _05702_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _05759_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _05763_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _05767_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _05771_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _05775_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _05779_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _05783_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _05752_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _05755_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _05812_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _05816_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _05820_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _05824_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _05828_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _05832_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _05836_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _05805_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _05808_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _05865_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _05869_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _05873_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _05877_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _05881_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _05885_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _05889_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _05858_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _05861_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _05187_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _05191_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _05195_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _05199_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _05203_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _05207_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _05211_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _05180_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _05183_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _05239_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _05243_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _05247_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _05251_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _05254_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _05258_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _05262_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _05232_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _05235_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _05290_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _05294_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _05298_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _05302_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _05306_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _05310_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _05314_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _05284_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _05287_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _05342_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _05346_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _05350_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _05354_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _05358_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _05362_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _05365_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _05335_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _05338_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _05394_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _05397_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _05401_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _05405_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _05409_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _05413_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _05417_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _05387_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _05390_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _05445_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _05449_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _05453_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _05457_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _05461_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _05465_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _05469_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _05438_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _05441_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _05497_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _05501_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _05505_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _05508_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _05512_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _05516_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _05520_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _05490_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _05493_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _05548_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _05552_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _05556_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _05560_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _05564_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _05568_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _05572_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _05541_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _05544_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _40533_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _40534_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _40535_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _40537_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _40538_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _40539_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _40540_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _40310_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _40522_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _40523_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _40524_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _40526_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _40527_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _40528_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _40529_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _40530_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _40510_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _40511_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _40512_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _40513_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _40515_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _40516_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _40517_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _40518_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _40498_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _40499_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _40500_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _40501_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _40503_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _40504_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _40505_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _40506_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _40485_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _40487_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _40488_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _40489_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _40490_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _40491_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _40493_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _40494_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _40473_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _40475_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _40476_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _40477_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _40478_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _40479_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _40481_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _40482_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _40461_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _40462_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _40464_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _40465_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _40466_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _40467_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _40468_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _40470_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _40449_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _40450_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _40452_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _40453_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _40454_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _40455_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _40456_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _40458_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _40437_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _40439_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _40440_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _40441_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _40442_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _40443_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _40445_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _40446_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _40424_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _40427_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _40428_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _40429_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _40430_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _40431_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _40433_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _40434_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _40412_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _40413_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _40416_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _40417_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _40418_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _40419_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _40420_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _40422_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _40401_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _40402_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _40404_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _40405_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _40406_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _40407_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _40408_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _40410_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _40388_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _40390_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _40391_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _40392_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _40393_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _40394_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _40396_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _40397_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _40376_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _40377_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _40379_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _40380_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _40381_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _40382_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _40383_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _40385_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _40362_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _40365_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _40366_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _40367_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _40368_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _40369_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _40371_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _40372_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _40350_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _40351_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _40352_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _40353_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _40354_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _40357_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _40358_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _40359_);
  dff (\oc8051_golden_model_1.B [0], _42890_);
  dff (\oc8051_golden_model_1.B [1], _42891_);
  dff (\oc8051_golden_model_1.B [2], _42892_);
  dff (\oc8051_golden_model_1.B [3], _42893_);
  dff (\oc8051_golden_model_1.B [4], _42894_);
  dff (\oc8051_golden_model_1.B [5], _42896_);
  dff (\oc8051_golden_model_1.B [6], _42897_);
  dff (\oc8051_golden_model_1.B [7], _40311_);
  dff (\oc8051_golden_model_1.ACC [0], _42898_);
  dff (\oc8051_golden_model_1.ACC [1], _42900_);
  dff (\oc8051_golden_model_1.ACC [2], _42901_);
  dff (\oc8051_golden_model_1.ACC [3], _42902_);
  dff (\oc8051_golden_model_1.ACC [4], _42903_);
  dff (\oc8051_golden_model_1.ACC [5], _42904_);
  dff (\oc8051_golden_model_1.ACC [6], _42905_);
  dff (\oc8051_golden_model_1.ACC [7], _40312_);
  dff (\oc8051_golden_model_1.PCON [0], _42907_);
  dff (\oc8051_golden_model_1.PCON [1], _42908_);
  dff (\oc8051_golden_model_1.PCON [2], _42909_);
  dff (\oc8051_golden_model_1.PCON [3], _42910_);
  dff (\oc8051_golden_model_1.PCON [4], _42911_);
  dff (\oc8051_golden_model_1.PCON [5], _42912_);
  dff (\oc8051_golden_model_1.PCON [6], _42913_);
  dff (\oc8051_golden_model_1.PCON [7], _40313_);
  dff (\oc8051_golden_model_1.TMOD [0], _42915_);
  dff (\oc8051_golden_model_1.TMOD [1], _42916_);
  dff (\oc8051_golden_model_1.TMOD [2], _42917_);
  dff (\oc8051_golden_model_1.TMOD [3], _42919_);
  dff (\oc8051_golden_model_1.TMOD [4], _42920_);
  dff (\oc8051_golden_model_1.TMOD [5], _42921_);
  dff (\oc8051_golden_model_1.TMOD [6], _42922_);
  dff (\oc8051_golden_model_1.TMOD [7], _40314_);
  dff (\oc8051_golden_model_1.DPL [0], _42924_);
  dff (\oc8051_golden_model_1.DPL [1], _42925_);
  dff (\oc8051_golden_model_1.DPL [2], _42926_);
  dff (\oc8051_golden_model_1.DPL [3], _42927_);
  dff (\oc8051_golden_model_1.DPL [4], _42928_);
  dff (\oc8051_golden_model_1.DPL [5], _42929_);
  dff (\oc8051_golden_model_1.DPL [6], _42930_);
  dff (\oc8051_golden_model_1.DPL [7], _40315_);
  dff (\oc8051_golden_model_1.DPH [0], _42932_);
  dff (\oc8051_golden_model_1.DPH [1], _42933_);
  dff (\oc8051_golden_model_1.DPH [2], _42934_);
  dff (\oc8051_golden_model_1.DPH [3], _42935_);
  dff (\oc8051_golden_model_1.DPH [4], _42936_);
  dff (\oc8051_golden_model_1.DPH [5], _42938_);
  dff (\oc8051_golden_model_1.DPH [6], _42939_);
  dff (\oc8051_golden_model_1.DPH [7], _40318_);
  dff (\oc8051_golden_model_1.TL1 [0], _42940_);
  dff (\oc8051_golden_model_1.TL1 [1], _42942_);
  dff (\oc8051_golden_model_1.TL1 [2], _42943_);
  dff (\oc8051_golden_model_1.TL1 [3], _42944_);
  dff (\oc8051_golden_model_1.TL1 [4], _42945_);
  dff (\oc8051_golden_model_1.TL1 [5], _42946_);
  dff (\oc8051_golden_model_1.TL1 [6], _42947_);
  dff (\oc8051_golden_model_1.TL1 [7], _40319_);
  dff (\oc8051_golden_model_1.TL0 [0], _42949_);
  dff (\oc8051_golden_model_1.TL0 [1], _42950_);
  dff (\oc8051_golden_model_1.TL0 [2], _42951_);
  dff (\oc8051_golden_model_1.TL0 [3], _42952_);
  dff (\oc8051_golden_model_1.TL0 [4], _42953_);
  dff (\oc8051_golden_model_1.TL0 [5], _42954_);
  dff (\oc8051_golden_model_1.TL0 [6], _42955_);
  dff (\oc8051_golden_model_1.TL0 [7], _40320_);
  dff (\oc8051_golden_model_1.TCON [0], _42957_);
  dff (\oc8051_golden_model_1.TCON [1], _42958_);
  dff (\oc8051_golden_model_1.TCON [2], _42959_);
  dff (\oc8051_golden_model_1.TCON [3], _42961_);
  dff (\oc8051_golden_model_1.TCON [4], _42962_);
  dff (\oc8051_golden_model_1.TCON [5], _42963_);
  dff (\oc8051_golden_model_1.TCON [6], _42964_);
  dff (\oc8051_golden_model_1.TCON [7], _40321_);
  dff (\oc8051_golden_model_1.TH1 [0], _42966_);
  dff (\oc8051_golden_model_1.TH1 [1], _42967_);
  dff (\oc8051_golden_model_1.TH1 [2], _42968_);
  dff (\oc8051_golden_model_1.TH1 [3], _42969_);
  dff (\oc8051_golden_model_1.TH1 [4], _42970_);
  dff (\oc8051_golden_model_1.TH1 [5], _42971_);
  dff (\oc8051_golden_model_1.TH1 [6], _42972_);
  dff (\oc8051_golden_model_1.TH1 [7], _40322_);
  dff (\oc8051_golden_model_1.TH0 [0], _42974_);
  dff (\oc8051_golden_model_1.TH0 [1], _42975_);
  dff (\oc8051_golden_model_1.TH0 [2], _42976_);
  dff (\oc8051_golden_model_1.TH0 [3], _42977_);
  dff (\oc8051_golden_model_1.TH0 [4], _42978_);
  dff (\oc8051_golden_model_1.TH0 [5], _42980_);
  dff (\oc8051_golden_model_1.TH0 [6], _42981_);
  dff (\oc8051_golden_model_1.TH0 [7], _40324_);
  dff (\oc8051_golden_model_1.PC [0], _42983_);
  dff (\oc8051_golden_model_1.PC [1], _42984_);
  dff (\oc8051_golden_model_1.PC [2], _42985_);
  dff (\oc8051_golden_model_1.PC [3], _42987_);
  dff (\oc8051_golden_model_1.PC [4], _42988_);
  dff (\oc8051_golden_model_1.PC [5], _42989_);
  dff (\oc8051_golden_model_1.PC [6], _42990_);
  dff (\oc8051_golden_model_1.PC [7], _42991_);
  dff (\oc8051_golden_model_1.PC [8], _42992_);
  dff (\oc8051_golden_model_1.PC [9], _42993_);
  dff (\oc8051_golden_model_1.PC [10], _42994_);
  dff (\oc8051_golden_model_1.PC [11], _42995_);
  dff (\oc8051_golden_model_1.PC [12], _42996_);
  dff (\oc8051_golden_model_1.PC [13], _42998_);
  dff (\oc8051_golden_model_1.PC [14], _42999_);
  dff (\oc8051_golden_model_1.PC [15], _40325_);
  dff (\oc8051_golden_model_1.P2 [0], _43000_);
  dff (\oc8051_golden_model_1.P2 [1], _43002_);
  dff (\oc8051_golden_model_1.P2 [2], _43003_);
  dff (\oc8051_golden_model_1.P2 [3], _43004_);
  dff (\oc8051_golden_model_1.P2 [4], _43005_);
  dff (\oc8051_golden_model_1.P2 [5], _43006_);
  dff (\oc8051_golden_model_1.P2 [6], _43007_);
  dff (\oc8051_golden_model_1.P2 [7], _40326_);
  dff (\oc8051_golden_model_1.P3 [0], _43009_);
  dff (\oc8051_golden_model_1.P3 [1], _43010_);
  dff (\oc8051_golden_model_1.P3 [2], _43011_);
  dff (\oc8051_golden_model_1.P3 [3], _43012_);
  dff (\oc8051_golden_model_1.P3 [4], _43013_);
  dff (\oc8051_golden_model_1.P3 [5], _43014_);
  dff (\oc8051_golden_model_1.P3 [6], _43015_);
  dff (\oc8051_golden_model_1.P3 [7], _40327_);
  dff (\oc8051_golden_model_1.P0 [0], _43017_);
  dff (\oc8051_golden_model_1.P0 [1], _43018_);
  dff (\oc8051_golden_model_1.P0 [2], _43019_);
  dff (\oc8051_golden_model_1.P0 [3], _43021_);
  dff (\oc8051_golden_model_1.P0 [4], _43022_);
  dff (\oc8051_golden_model_1.P0 [5], _43023_);
  dff (\oc8051_golden_model_1.P0 [6], _43024_);
  dff (\oc8051_golden_model_1.P0 [7], _40328_);
  dff (\oc8051_golden_model_1.P1 [0], _43026_);
  dff (\oc8051_golden_model_1.P1 [1], _43027_);
  dff (\oc8051_golden_model_1.P1 [2], _43028_);
  dff (\oc8051_golden_model_1.P1 [3], _43029_);
  dff (\oc8051_golden_model_1.P1 [4], _43030_);
  dff (\oc8051_golden_model_1.P1 [5], _43031_);
  dff (\oc8051_golden_model_1.P1 [6], _43032_);
  dff (\oc8051_golden_model_1.P1 [7], _40330_);
  dff (\oc8051_golden_model_1.IP [0], _43034_);
  dff (\oc8051_golden_model_1.IP [1], _43035_);
  dff (\oc8051_golden_model_1.IP [2], _43036_);
  dff (\oc8051_golden_model_1.IP [3], _43037_);
  dff (\oc8051_golden_model_1.IP [4], _43038_);
  dff (\oc8051_golden_model_1.IP [5], _43040_);
  dff (\oc8051_golden_model_1.IP [6], _43041_);
  dff (\oc8051_golden_model_1.IP [7], _40331_);
  dff (\oc8051_golden_model_1.IE [0], _43042_);
  dff (\oc8051_golden_model_1.IE [1], _43044_);
  dff (\oc8051_golden_model_1.IE [2], _43045_);
  dff (\oc8051_golden_model_1.IE [3], _43046_);
  dff (\oc8051_golden_model_1.IE [4], _43047_);
  dff (\oc8051_golden_model_1.IE [5], _43048_);
  dff (\oc8051_golden_model_1.IE [6], _43049_);
  dff (\oc8051_golden_model_1.IE [7], _40332_);
  dff (\oc8051_golden_model_1.SCON [0], _43051_);
  dff (\oc8051_golden_model_1.SCON [1], _43052_);
  dff (\oc8051_golden_model_1.SCON [2], _43053_);
  dff (\oc8051_golden_model_1.SCON [3], _43054_);
  dff (\oc8051_golden_model_1.SCON [4], _43055_);
  dff (\oc8051_golden_model_1.SCON [5], _43056_);
  dff (\oc8051_golden_model_1.SCON [6], _43057_);
  dff (\oc8051_golden_model_1.SCON [7], _40333_);
  dff (\oc8051_golden_model_1.SP [0], _43059_);
  dff (\oc8051_golden_model_1.SP [1], _43060_);
  dff (\oc8051_golden_model_1.SP [2], _43061_);
  dff (\oc8051_golden_model_1.SP [3], _43063_);
  dff (\oc8051_golden_model_1.SP [4], _43064_);
  dff (\oc8051_golden_model_1.SP [5], _43065_);
  dff (\oc8051_golden_model_1.SP [6], _43066_);
  dff (\oc8051_golden_model_1.SP [7], _40334_);
  dff (\oc8051_golden_model_1.SBUF [0], _43068_);
  dff (\oc8051_golden_model_1.SBUF [1], _43069_);
  dff (\oc8051_golden_model_1.SBUF [2], _43070_);
  dff (\oc8051_golden_model_1.SBUF [3], _43071_);
  dff (\oc8051_golden_model_1.SBUF [4], _43072_);
  dff (\oc8051_golden_model_1.SBUF [5], _43073_);
  dff (\oc8051_golden_model_1.SBUF [6], _43074_);
  dff (\oc8051_golden_model_1.SBUF [7], _40336_);
  dff (\oc8051_golden_model_1.PSW [0], _43075_);
  dff (\oc8051_golden_model_1.PSW [1], _43076_);
  dff (\oc8051_golden_model_1.PSW [2], _43077_);
  dff (\oc8051_golden_model_1.PSW [3], _43078_);
  dff (\oc8051_golden_model_1.PSW [4], _43079_);
  dff (\oc8051_golden_model_1.PSW [5], _43081_);
  dff (\oc8051_golden_model_1.PSW [6], _43082_);
  dff (\oc8051_golden_model_1.PSW [7], _40337_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02839_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02851_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02873_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02897_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02919_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00955_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02931_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00925_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02943_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02957_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02971_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02984_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _02998_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03011_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03023_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00974_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02358_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22126_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02546_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02702_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02884_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03126_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03330_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03531_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03732_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03929_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04027_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04126_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04226_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04325_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04419_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04517_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04616_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24284_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38395_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38397_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38398_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38399_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38400_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38401_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38402_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38381_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38403_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38404_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38406_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38407_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38408_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38409_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38410_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38382_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38412_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38413_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38414_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38415_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38416_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38418_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38419_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38384_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34185_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34188_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09685_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34190_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34192_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09688_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34194_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09691_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34196_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34198_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34200_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09694_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34202_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09697_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _09700_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09759_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09761_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09664_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09764_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09767_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09667_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _09770_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _09670_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _09773_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _09776_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09779_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09782_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09785_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09788_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09791_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _09673_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09676_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34183_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09682_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09794_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09679_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39196_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39294_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39295_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39296_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39297_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39298_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39299_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39300_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39197_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39301_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39302_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39303_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39305_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39306_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39307_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39308_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39198_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39309_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39310_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39311_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39312_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39313_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39314_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39316_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39199_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39317_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39318_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39319_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39320_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39321_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39322_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39323_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39201_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _39324_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _39325_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _39327_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _39328_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _39329_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _39330_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _39331_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _39202_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _39332_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _39333_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _39334_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _39335_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _39336_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _39338_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _39339_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _39203_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _39340_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _39341_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _39342_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _39343_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _39344_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _39345_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _39346_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _39204_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _39347_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _39349_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _39350_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _39351_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _39352_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _39353_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _39354_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _39205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _38766_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _38767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _38768_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _38769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38482_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38555_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38556_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38557_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38558_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38559_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38561_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38562_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38563_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38564_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38565_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38567_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38568_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _38569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _38570_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _38575_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _38576_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _38577_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _38578_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _38579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _38580_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _38581_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _38582_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _38583_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _38584_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _38586_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _38587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _38588_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _38589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _38590_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _38770_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _38771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _38772_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _38773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _38775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _38776_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _38777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _38778_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _38779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _38780_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _38781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _38782_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _38783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _38784_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _38786_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _38787_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _38788_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _38789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _38790_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _38791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _38792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _38793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _38794_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _38795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _38797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _38798_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _38799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _38800_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _38801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _38802_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _38803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38506_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38480_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _38804_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _38806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _38807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _38808_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _38809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _38810_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _38812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38483_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _38813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _38814_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _38815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _38816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _38817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _38818_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _38819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38484_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _38820_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _38821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _38823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _38824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _38825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _38826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _38827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38486_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38487_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38488_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _38828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _38829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _38830_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _38831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _38832_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _38834_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _38835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38489_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _38836_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _38837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _38838_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _38839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _38840_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _38841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _38842_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _38843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _38845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _38846_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _38847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _38848_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _38849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _38850_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _38851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38490_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _38852_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _38853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _38854_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _38855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _38856_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _38857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _38858_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _38859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _38860_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _38861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _38862_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _38863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _38864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _38866_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _38867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38492_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38493_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38495_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38494_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _38868_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _38869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _38870_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _38871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _38872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _38873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _38874_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38497_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _38875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _38877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38498_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _38878_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _38879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _38880_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _38881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _38882_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _38883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _38884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38499_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _38885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _38886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _38888_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _38889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _38890_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _38891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _38892_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38500_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _38501_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _38893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _38894_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _38895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _38896_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _38897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _38899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _38900_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _38503_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38504_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _38901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _38902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _38903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38505_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _38904_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _38905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _38906_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _38907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _38908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _38910_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _38911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _38912_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _38913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _38914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _38915_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _38916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _38917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _38918_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _38919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _38921_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _38922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _38923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _38924_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _38925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _38926_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _38927_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _38928_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _38929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _38930_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _38932_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _38933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _38934_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _38935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _38936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _38937_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38507_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _38938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _38939_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _38940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _38941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _38943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _38944_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _38945_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38508_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38509_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38511_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _38946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _38947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _38948_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _38949_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _38950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _38951_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _38952_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _38954_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _38955_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _38956_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _38957_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _38958_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _38959_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _38960_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _38961_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38512_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38513_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38514_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38515_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _38962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _38963_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _38965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _38966_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _38967_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _38968_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _38969_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _38970_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _38971_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _38972_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _38973_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _38974_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _38976_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _38977_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _38978_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38516_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38517_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39582_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39602_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39603_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39604_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39605_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39606_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39607_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39608_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39583_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39584_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39609_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39610_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _03001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02567_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _39418_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _39502_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _39503_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _39504_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _39420_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _39421_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _39422_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39506_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39507_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39508_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39509_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39510_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39511_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39512_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39423_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19771_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19783_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19807_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17968_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08905_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08938_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13662_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13672_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12682_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13716_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13738_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _42360_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _42358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _42355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _42351_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _42349_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _42347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _42345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _42306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _42304_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _42302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _42300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _42298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00171_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _42296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00175_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00177_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _42293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40047_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40056_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40058_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40060_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40062_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40068_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40070_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31058_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40079_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40081_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31081_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40089_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40091_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40093_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40095_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40099_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31103_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17377_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17399_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09488_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10676_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09509_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40552_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41062_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41067_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41069_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41071_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41073_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _40555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41079_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41081_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41084_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _40558_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _40561_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _40564_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41088_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41096_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _40567_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41101_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41103_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41105_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _40570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _40573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _40576_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01632_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02110_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02112_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02129_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02131_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01653_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01656_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01659_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01227_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01229_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00567_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00546_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01232_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01238_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01240_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01244_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00581_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01260_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01262_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01267_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01285_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01287_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01291_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01299_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01301_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00591_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1071 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1071 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1071 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1071 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1073 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1075 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1075 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1076 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1076 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1077 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1077 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1078 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1078 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1079 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1079 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1080 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1080 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1081 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1118 , \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.n1146 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1147 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1147 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1147 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1147 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1147 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1147 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1148 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1148 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1148 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1148 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1148 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1148 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1149 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1149 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1149 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1149 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1149 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1149 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1149 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1150 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1151 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1152 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1152 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1152 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1153 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1154 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1154 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1155 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1155 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1155 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1155 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1155 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1155 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1181 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1181 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1181 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1181 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1181 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1181 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1181 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1181 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1181 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1181 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1181 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1181 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1181 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1183 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1183 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1183 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1183 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1183 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1183 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1185 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1185 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1185 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1185 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1185 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1185 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1185 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1189 [8], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1190 , \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1191 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1191 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1191 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1191 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1192 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1192 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1192 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1196 [4], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1197 , \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1198 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1198 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1198 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1198 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1198 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1198 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1198 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1198 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1198 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1206 , \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.n1207 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1207 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1207 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1207 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1207 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1212 , \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1217 [4], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1218 , \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1226 , \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.n1227 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1227 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1227 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1227 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1227 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1229 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1229 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1229 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1229 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1229 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1229 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1229 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1229 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1229 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1231 [8], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1232 , \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1233 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1233 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1233 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1233 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1234 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1234 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1234 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1236 [4], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1249 [8], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1257 , \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.n1258 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1258 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1258 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1258 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1258 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1260 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1262 [8], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1276 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1278 [4], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1279 , \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1280 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1280 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1280 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1280 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1280 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1280 [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1282 [8], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1290 , \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1291 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1291 [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1291 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1291 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1291 [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1292 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1292 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1292 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1292 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1292 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1295 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1295 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1295 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1295 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1295 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1295 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1295 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1295 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1295 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1296 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1296 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1296 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1296 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1296 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1296 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1297 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1297 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1297 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1297 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1297 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1297 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1297 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1297 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1298 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1299 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1299 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1299 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1299 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1299 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1299 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1299 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1299 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1300 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1300 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1303 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1305 [8], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1306 , \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1307 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1307 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1309 [4], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1310 , \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.n1318 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1318 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1318 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1318 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1318 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1322 [8], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1323 , \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.n1334 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1334 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1334 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1334 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1334 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1338 [8], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1339 , \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1350 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1350 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1354 [8], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1357 [4], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1358 , \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1365 , \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1520 , \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1521 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1521 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1521 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1521 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1521 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1521 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1521 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1680 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1683 , \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.n1691 , \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.n1692 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1692 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1692 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1692 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1692 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1696 , \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.n1698 , \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1709 , \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.n1711 , \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.n1717 , \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.n1718 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1718 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1718 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1718 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1718 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 , \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.n1724 , \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.n1730 , \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1733 , \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.n1734 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1734 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1734 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1734 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1734 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1734 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1734 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1739 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1739 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1739 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1739 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1739 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1739 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1739 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1739 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1739 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1745 , \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.n1746 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1746 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1746 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1746 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1746 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1746 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1746 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1749 , \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.n1750 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1750 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1750 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1750 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1750 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1750 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1750 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1765 , \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.n1766 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1766 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1766 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1766 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1766 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1766 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1766 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1771 , \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.n1772 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1772 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1772 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1772 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1772 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1772 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1772 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.n1778 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1778 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1778 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1778 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1778 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1778 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1778 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1783 , \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.n1784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1791 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1791 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1791 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1791 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1791 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1791 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1792 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1792 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1792 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1792 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1793 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1793 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1793 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1793 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1793 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1793 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1828 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1828 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1828 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1828 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1828 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1828 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1828 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1828 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1847 , \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.n1848 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1848 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1848 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1848 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1848 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1848 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1848 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1852 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1854 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1854 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1854 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1854 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
