
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pcp1, property_invalid_pcp2, property_invalid_pcp3, property_invalid_sjmp, property_invalid_ljmp, property_invalid_ajmp, property_invalid_jc, property_invalid_jnc);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire [15:0] _28201_;
  wire [7:0] _28202_;
  wire [7:0] _28203_;
  wire [7:0] _28204_;
  wire [7:0] _28205_;
  wire [7:0] _28206_;
  wire [7:0] _28207_;
  wire [7:0] _28208_;
  wire [7:0] _28209_;
  wire [7:0] _28210_;
  wire [7:0] _28211_;
  wire [7:0] _28212_;
  wire [7:0] _28213_;
  wire [7:0] _28214_;
  wire [7:0] _28215_;
  wire [7:0] _28216_;
  wire [7:0] _28217_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_ajmp;
  output property_invalid_jc;
  output property_invalid_jnc;
  output property_invalid_ljmp;
  output property_invalid_pcp1;
  output property_invalid_pcp2;
  output property_invalid_pcp3;
  output property_invalid_sjmp;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [31:0] word_in;
  not (_23914_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_23915_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _23914_);
  and (_23916_, _23915_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23917_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _23914_);
  and (_23918_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _23914_);
  nor (_23919_, _23918_, _23917_);
  and (_23920_, _23919_, _23916_);
  not (_23921_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_23922_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _23921_);
  not (_23923_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_23924_, _23923_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nor (_23925_, _23924_, _23922_);
  nand (_23926_, _23925_, _23920_);
  not (_27355_, rst);
  or (_23927_, _23920_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_23928_, _23927_, _27355_);
  and (_23530_, _23928_, _23926_);
  nor (_23929_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_23930_, _23929_);
  and (_23931_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not (_23932_, _23931_);
  and (_23933_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_23934_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_23935_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_23936_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_23937_, _23936_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_23938_, _23937_, _23935_);
  or (_23939_, _23938_, _23934_);
  not (_23940_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_23941_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_23942_, _23941_, _23935_);
  or (_23943_, _23942_, _23940_);
  and (_23944_, _23943_, _23939_);
  or (_23945_, _23937_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_23946_, _23945_);
  nand (_23947_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_23948_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_23949_, _23948_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_23950_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_23951_, _23950_, _23947_);
  and (_23952_, _23951_, _23944_);
  not (_23953_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_23954_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23953_);
  or (_23955_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  not (_23956_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23957_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23956_);
  and (_23958_, _23957_, _23955_);
  or (_23959_, _23958_, _23954_);
  nand (_23960_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23953_);
  or (_23961_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_23962_, _23961_, _23959_);
  or (_23963_, _23941_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23964_, _23963_, _23962_);
  not (_23965_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_23966_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_23967_, _23966_, _23935_);
  or (_23968_, _23967_, _23965_);
  and (_23969_, _23966_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_23970_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_23971_, _23970_, _23968_);
  and (_23972_, _23971_, _23964_);
  and (_23973_, _23972_, _23952_);
  not (_23974_, _23973_);
  or (_23975_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_23976_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or (_23977_, _23956_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_23978_, _23977_, _23976_);
  or (_23979_, _23978_, _23954_);
  or (_23980_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_23981_, _23980_, _23979_);
  or (_23982_, _23981_, _23975_);
  and (_23983_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_23984_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_23985_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_23986_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_23987_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _23986_);
  nor (_23988_, _23987_, _23985_);
  nor (_23989_, _23988_, _23984_);
  and (_23990_, _23989_, _23982_);
  nand (_23991_, _23990_, _23929_);
  not (_23992_, _23922_);
  or (_23993_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_23994_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23956_);
  and (_23995_, _23994_, _23993_);
  or (_23996_, _23995_, _23954_);
  or (_23997_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_23998_, _23997_, _23996_);
  or (_23999_, _23998_, _23975_);
  nand (_24000_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not (_24001_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_24002_, _23987_, _24001_);
  and (_24003_, _24002_, _24000_);
  and (_24004_, _24003_, _23999_);
  or (_24005_, _24004_, _23992_);
  not (_24006_, _23924_);
  or (_24007_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_24008_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23956_);
  and (_24009_, _24008_, _24007_);
  or (_24010_, _24009_, _23954_);
  or (_24011_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_24012_, _24011_, _24010_);
  or (_24013_, _24012_, _23975_);
  nand (_24014_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not (_24015_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_24016_, _23987_, _24015_);
  and (_24017_, _24016_, _24014_);
  and (_24018_, _24017_, _24013_);
  or (_24019_, _24018_, _24006_);
  and (_24020_, _24019_, _24005_);
  or (_24021_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_24022_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23956_);
  and (_24023_, _24022_, _24021_);
  or (_24024_, _24023_, _23954_);
  or (_24025_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_24026_, _24025_, _24024_);
  or (_24027_, _24026_, _23975_);
  nand (_24028_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not (_24029_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_24030_, _23987_, _24029_);
  and (_24031_, _24030_, _24028_);
  nand (_24032_, _24031_, _24027_);
  or (_24033_, _24032_, _23921_);
  nand (_24034_, _24033_, _23925_);
  nand (_24035_, _24034_, _24020_);
  and (_24036_, _24035_, _23991_);
  and (_24037_, _24036_, _23974_);
  or (_24038_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_24039_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23956_);
  and (_24040_, _24039_, _24038_);
  or (_24041_, _24040_, _23954_);
  or (_24042_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_24043_, _24042_, _24041_);
  or (_24044_, _24043_, _23975_);
  nand (_24045_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_24046_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_24047_, _23987_, _24046_);
  and (_24048_, _24047_, _24045_);
  nand (_24049_, _24048_, _24044_);
  or (_24050_, _24049_, _23930_);
  or (_24051_, _23962_, _23975_);
  nand (_24052_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_24053_, _23987_, _23965_);
  and (_24054_, _24053_, _24052_);
  and (_24055_, _24054_, _24051_);
  or (_24056_, _24055_, _23992_);
  or (_24057_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_24058_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23956_);
  and (_24059_, _24058_, _24057_);
  or (_24060_, _24059_, _23954_);
  or (_24061_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_24062_, _24061_, _24060_);
  or (_24063_, _24062_, _23975_);
  nand (_24064_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_24065_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_24066_, _23987_, _24065_);
  and (_24067_, _24066_, _24064_);
  and (_24068_, _24067_, _24063_);
  or (_24069_, _24068_, _24006_);
  and (_24070_, _24069_, _24056_);
  or (_24071_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_24072_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23956_);
  and (_24073_, _24072_, _24071_);
  or (_24074_, _24073_, _23954_);
  or (_24075_, _23960_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_24076_, _24075_, _24074_);
  or (_24077_, _24076_, _23975_);
  nand (_24078_, _23983_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not (_24079_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_24080_, _23987_, _24079_);
  and (_24081_, _24080_, _24078_);
  nand (_24082_, _24081_, _24077_);
  or (_24083_, _24082_, _23921_);
  nand (_24084_, _24083_, _23925_);
  nand (_24085_, _24084_, _24070_);
  and (_24086_, _24085_, _24050_);
  not (_24087_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_24088_, _23938_, _24087_);
  not (_24089_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_24090_, _23942_, _24089_);
  and (_24091_, _24090_, _24088_);
  nand (_24092_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nand (_24093_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_24094_, _24093_, _24092_);
  and (_24095_, _24094_, _24091_);
  or (_24096_, _24012_, _23963_);
  or (_24097_, _23967_, _24015_);
  nand (_24098_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_24099_, _24098_, _24097_);
  and (_24100_, _24099_, _24096_);
  and (_24101_, _24100_, _24095_);
  not (_24102_, _24101_);
  and (_24103_, _24102_, _24086_);
  and (_24104_, _24103_, _24037_);
  and (_24105_, _23974_, _24086_);
  not (_24106_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_24107_, _23938_, _24106_);
  not (_24108_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_24109_, _23942_, _24108_);
  and (_24110_, _24109_, _24107_);
  nand (_24111_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nand (_24112_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_24113_, _24112_, _24111_);
  and (_24114_, _24113_, _24110_);
  or (_24115_, _23998_, _23963_);
  nand (_24116_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  or (_24117_, _23967_, _24001_);
  and (_24118_, _24117_, _24116_);
  and (_24119_, _24118_, _24115_);
  nand (_24120_, _24119_, _24114_);
  and (_24121_, _24120_, _24036_);
  nand (_24122_, _24121_, _24105_);
  and (_24123_, _24120_, _24086_);
  or (_24124_, _24123_, _24037_);
  and (_24125_, _24124_, _24122_);
  and (_24126_, _24125_, _24104_);
  not (_24127_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_24128_, _23938_, _24127_);
  not (_24129_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_24130_, _23942_, _24129_);
  and (_24131_, _24130_, _24128_);
  nand (_24132_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nand (_24133_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_24134_, _24133_, _24132_);
  and (_24135_, _24134_, _24131_);
  or (_24136_, _23963_, _24043_);
  or (_24137_, _23967_, _24046_);
  nand (_24138_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_24139_, _24138_, _24137_);
  and (_24140_, _24139_, _24136_);
  and (_24141_, _24140_, _24135_);
  or (_24142_, _24141_, _24122_);
  not (_24143_, _24141_);
  and (_24144_, _24143_, _24086_);
  not (_24145_, _24144_);
  nand (_24146_, _24145_, _24122_);
  and (_24147_, _24146_, _24142_);
  nand (_24148_, _24147_, _24121_);
  or (_24149_, _24144_, _24121_);
  and (_24150_, _24149_, _24148_);
  nand (_24151_, _24150_, _24126_);
  not (_24152_, _24151_);
  not (_24153_, _24142_);
  and (_24154_, _24147_, _24121_);
  nand (_24155_, _24035_, _23991_);
  or (_24156_, _24141_, _24155_);
  nand (_24157_, _24085_, _24050_);
  not (_24158_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_24159_, _23942_, _24158_);
  not (_24160_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_24161_, _23938_, _24160_);
  and (_24162_, _24161_, _24159_);
  or (_24163_, _23967_, _23985_);
  nand (_24164_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_24165_, _24164_, _24163_);
  and (_24166_, _24165_, _24162_);
  or (_24167_, _23981_, _23963_);
  nand (_24168_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nand (_24169_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_24170_, _24169_, _24168_);
  and (_24171_, _24170_, _24167_);
  and (_24172_, _24171_, _24166_);
  or (_24173_, _24172_, _24157_);
  or (_24174_, _24173_, _24156_);
  nand (_24175_, _24173_, _24156_);
  and (_24176_, _24175_, _24174_);
  nand (_24177_, _24176_, _24154_);
  or (_24178_, _24176_, _24154_);
  and (_24179_, _24178_, _24177_);
  nand (_24180_, _24179_, _24153_);
  or (_24181_, _24179_, _24153_);
  and (_24182_, _24181_, _24180_);
  nand (_24183_, _24182_, _24152_);
  or (_24184_, _24182_, _24152_);
  nand (_24185_, _24184_, _24183_);
  not (_24186_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_24187_, _23938_, _24186_);
  not (_24188_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_24189_, _23942_, _24188_);
  and (_24190_, _24189_, _24187_);
  nand (_24191_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nand (_24192_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_24193_, _24192_, _24191_);
  and (_24194_, _24193_, _24190_);
  or (_24195_, _24026_, _23963_);
  or (_24196_, _23967_, _24029_);
  nand (_24197_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_24198_, _24197_, _24196_);
  and (_24199_, _24198_, _24195_);
  nand (_24200_, _24199_, _24194_);
  and (_24201_, _24200_, _24036_);
  not (_24202_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_24203_, _23938_, _24202_);
  not (_24204_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_24205_, _23942_, _24204_);
  and (_24206_, _24205_, _24203_);
  nand (_24207_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  or (_24208_, _23967_, _24065_);
  and (_24209_, _24208_, _24207_);
  and (_24210_, _24209_, _24206_);
  or (_24211_, _23963_, _24062_);
  nand (_24212_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand (_24213_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_24214_, _24213_, _24212_);
  and (_24215_, _24214_, _24211_);
  nand (_24216_, _24215_, _24210_);
  and (_24217_, _24216_, _24086_);
  and (_24218_, _24217_, _24201_);
  not (_24219_, _24218_);
  and (_24220_, _24200_, _24086_);
  not (_24221_, _24220_);
  and (_24222_, _24216_, _24036_);
  and (_24223_, _24222_, _24221_);
  nand (_24224_, _24223_, _24103_);
  nand (_24225_, _24224_, _24219_);
  not (_24226_, _24104_);
  and (_24227_, _24102_, _24036_);
  or (_24228_, _24227_, _24105_);
  and (_24229_, _24228_, _24226_);
  and (_24230_, _24229_, _24225_);
  not (_24231_, _24126_);
  or (_24232_, _24125_, _24104_);
  and (_24233_, _24232_, _24231_);
  and (_24234_, _24233_, _24230_);
  or (_24235_, _24150_, _24126_);
  and (_24236_, _24235_, _24151_);
  nand (_24237_, _24236_, _24234_);
  not (_24238_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_24239_, _23938_, _24238_);
  not (_24240_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_24241_, _23942_, _24240_);
  nor (_24242_, _24241_, _24239_);
  and (_24243_, _23946_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_24244_, _23949_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_24245_, _24244_, _24243_);
  and (_24246_, _24245_, _24242_);
  nor (_24247_, _23963_, _24076_);
  nor (_24248_, _23967_, _24079_);
  and (_24249_, _23969_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_24250_, _24249_, _24248_);
  not (_24251_, _24250_);
  nor (_24252_, _24251_, _24247_);
  and (_24253_, _24252_, _24246_);
  not (_24254_, _24253_);
  and (_24255_, _24254_, _24036_);
  and (_24256_, _24255_, _24220_);
  or (_24257_, _24217_, _24201_);
  and (_24258_, _24257_, _24219_);
  and (_24259_, _24258_, _24256_);
  or (_24260_, _24223_, _24103_);
  and (_24261_, _24260_, _24224_);
  nand (_24262_, _24261_, _24259_);
  not (_24263_, _24262_);
  nand (_24264_, _24229_, _24225_);
  or (_24265_, _24229_, _24225_);
  and (_24266_, _24265_, _24264_);
  nand (_24267_, _24266_, _24263_);
  nand (_24268_, _24233_, _24230_);
  or (_24269_, _24233_, _24230_);
  nand (_24270_, _24269_, _24268_);
  or (_24271_, _24270_, _24267_);
  or (_24272_, _24236_, _24234_);
  nand (_24273_, _24272_, _24237_);
  or (_24274_, _24273_, _24271_);
  and (_24275_, _24274_, _24237_);
  or (_24276_, _24275_, _24185_);
  nand (_24277_, _24276_, _24183_);
  not (_24278_, _24172_);
  and (_24279_, _24278_, _24036_);
  and (_24280_, _24279_, _24145_);
  and (_24281_, _24180_, _24177_);
  not (_24282_, _24281_);
  nand (_24283_, _24282_, _24280_);
  or (_24284_, _24282_, _24280_);
  and (_24285_, _24284_, _24283_);
  nand (_24286_, _24285_, _24277_);
  and (_24287_, _24283_, _24174_);
  nand (_24288_, _24287_, _24286_);
  nand (_24289_, _24288_, _23933_);
  or (_24290_, _24288_, _23933_);
  nand (_24291_, _24290_, _24289_);
  and (_24292_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or (_24293_, _24285_, _24277_);
  and (_24294_, _24293_, _24286_);
  nand (_24295_, _24294_, _24292_);
  or (_24296_, _24295_, _24291_);
  nand (_24297_, _24296_, _24289_);
  and (_24298_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_24299_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_24300_, _24299_, _24298_);
  and (_24301_, _24300_, _24297_);
  and (_24302_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand (_24303_, _24275_, _24185_);
  and (_24304_, _24303_, _24276_);
  nand (_24305_, _24304_, _24302_);
  or (_24309_, _24304_, _24302_);
  and (_24310_, _24309_, _24305_);
  and (_24311_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nand (_24312_, _24273_, _24271_);
  and (_24313_, _24312_, _24274_);
  nand (_24314_, _24313_, _24311_);
  or (_24315_, _24313_, _24311_);
  nand (_24316_, _24315_, _24314_);
  and (_24317_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nand (_24318_, _24270_, _24267_);
  and (_24319_, _24318_, _24271_);
  nand (_24326_, _24319_, _24317_);
  or (_24332_, _24319_, _24317_);
  and (_24338_, _24332_, _24326_);
  and (_24344_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or (_24345_, _24266_, _24263_);
  and (_24346_, _24345_, _24267_);
  nand (_24347_, _24346_, _24344_);
  and (_24348_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_24349_, _24261_, _24259_);
  and (_24350_, _24349_, _24262_);
  nand (_24351_, _24350_, _24348_);
  and (_24352_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_24353_, _24258_, _24256_);
  or (_24354_, _24258_, _24256_);
  and (_24355_, _24354_, _24353_);
  and (_24356_, _24355_, _24352_);
  not (_24357_, _24356_);
  or (_24358_, _24350_, _24348_);
  nand (_24359_, _24358_, _24351_);
  or (_24360_, _24359_, _24357_);
  nand (_24361_, _24360_, _24351_);
  or (_24362_, _24346_, _24344_);
  and (_24363_, _24362_, _24347_);
  nand (_24364_, _24363_, _24361_);
  nand (_24365_, _24364_, _24347_);
  nand (_24366_, _24365_, _24338_);
  and (_24367_, _24366_, _24326_);
  or (_24368_, _24367_, _24316_);
  nand (_24369_, _24368_, _24314_);
  nand (_24371_, _24369_, _24310_);
  and (_24373_, _24371_, _24305_);
  and (_24374_, _24290_, _24289_);
  or (_24375_, _24294_, _24292_);
  and (_24376_, _24375_, _24295_);
  and (_24377_, _24376_, _24374_);
  nand (_24378_, _24300_, _24377_);
  nor (_24379_, _24378_, _24373_);
  or (_24380_, _24379_, _24301_);
  and (_24381_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_24382_, _23930_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_24383_, _24382_, _24381_);
  nand (_24384_, _24383_, _24380_);
  nor (_24385_, _24384_, _23932_);
  not (_24386_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or (_24387_, _23929_, _24386_);
  nor (_24388_, _24387_, _24385_);
  and (_24389_, _24385_, _24386_);
  or (_24390_, _24389_, _24388_);
  and (_23899_, _24390_, _27355_);
  nor (_24391_, _23920_, _23923_);
  and (_24392_, _23920_, _23923_);
  or (_24393_, _24392_, _24391_);
  and (_02784_, _24393_, _27355_);
  and (_24394_, _24254_, _24086_);
  and (_02984_, _24394_, _27355_);
  nor (_24395_, _24255_, _24220_);
  nor (_24396_, _24395_, _24256_);
  and (_03157_, _24396_, _27355_);
  nor (_24397_, _24355_, _24352_);
  nor (_24398_, _24397_, _24356_);
  and (_03302_, _24398_, _27355_);
  and (_24399_, _24359_, _24357_);
  not (_24400_, _24399_);
  and (_24401_, _24400_, _24360_);
  and (_03443_, _24401_, _27355_);
  or (_24402_, _24363_, _24361_);
  and (_24403_, _24402_, _24364_);
  and (_03584_, _24403_, _27355_);
  or (_24408_, _24365_, _24338_);
  and (_24413_, _24408_, _24366_);
  and (_03782_, _24413_, _27355_);
  and (_24425_, _24367_, _24316_);
  not (_24432_, _24425_);
  and (_24441_, _24432_, _24368_);
  and (_03985_, _24441_, _27355_);
  or (_24442_, _24369_, _24310_);
  and (_24443_, _24442_, _24371_);
  and (_04190_, _24443_, _27355_);
  not (_24444_, _24376_);
  or (_24445_, _24444_, _24373_);
  not (_24446_, _24445_);
  and (_24447_, _24444_, _24373_);
  nor (_24448_, _24447_, _24446_);
  and (_04293_, _24448_, _27355_);
  and (_24449_, _24445_, _24295_);
  or (_24450_, _24449_, _24291_);
  nand (_24451_, _24449_, _24291_);
  and (_24452_, _24451_, _24450_);
  and (_04397_, _24452_, _27355_);
  nand (_24453_, _24450_, _24289_);
  nand (_24454_, _24453_, _24298_);
  or (_24455_, _24453_, _24298_);
  and (_24456_, _24455_, _24454_);
  and (_04499_, _24456_, _27355_);
  not (_24457_, _24380_);
  not (_24458_, _24299_);
  nand (_24459_, _24458_, _24454_);
  and (_24460_, _24459_, _24457_);
  and (_04604_, _24460_, _27355_);
  and (_24461_, _24381_, _24380_);
  nor (_24462_, _24381_, _24380_);
  nor (_24463_, _24462_, _24461_);
  and (_04707_, _24463_, _27355_);
  or (_24464_, _24382_, _24461_);
  and (_24465_, _24464_, _24384_);
  and (_04810_, _24465_, _27355_);
  and (_24466_, _24384_, _23932_);
  or (_24467_, _24466_, _24385_);
  nor (_04914_, _24467_, rst);
  and (_24468_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _23914_);
  nor (_24469_, _24468_, _23915_);
  not (_24471_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_24482_, _23917_, _24471_);
  and (_24487_, _24482_, _24469_);
  and (_24488_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24489_, _24488_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24496_, _24488_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_24506_, _24496_, _24489_);
  and (_00958_, _24506_, _27355_);
  and (_00985_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _27355_);
  nor (_24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_24508_, _24507_, _24172_);
  nor (_24509_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_24510_, _24509_);
  and (_24511_, _24510_, _24508_);
  not (_24512_, _24511_);
  or (_24513_, _24082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_24514_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24515_, _24067_, _24063_);
  or (_24516_, _24515_, _24514_);
  and (_24517_, _24516_, _24513_);
  or (_24518_, _24517_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24519_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_24520_, _24054_, _24051_);
  or (_24521_, _24520_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24522_, _24049_, _24514_);
  and (_24523_, _24522_, _24521_);
  or (_24524_, _24523_, _24519_);
  and (_24525_, _24524_, _24518_);
  or (_24526_, _24525_, _24512_);
  nand (_24527_, _24507_, _24141_);
  nor (_24528_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_24529_, _24528_);
  and (_24530_, _24529_, _24527_);
  and (_24531_, _24032_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24532_, _24531_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_24533_, _24017_, _24013_);
  or (_24534_, _24533_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24535_, _24003_, _23999_);
  or (_24536_, _24535_, _24514_);
  and (_24537_, _24536_, _24534_);
  or (_24538_, _24537_, _24519_);
  nand (_24539_, _24538_, _24532_);
  nand (_24540_, _24539_, _24530_);
  nand (_24541_, _24524_, _24518_);
  or (_24542_, _24541_, _24511_);
  and (_24543_, _24542_, _24526_);
  not (_24544_, _24543_);
  or (_24545_, _24544_, _24540_);
  and (_24546_, _24545_, _24526_);
  or (_24547_, _24539_, _24530_);
  and (_24548_, _24547_, _24540_);
  and (_24549_, _24548_, _24543_);
  not (_24550_, _24507_);
  or (_24551_, _24550_, _24120_);
  nor (_24552_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_24553_, _24552_);
  nand (_24554_, _24553_, _24551_);
  and (_24555_, _24082_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24556_, _24555_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24557_, _24515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24558_, _24520_, _24514_);
  and (_24559_, _24558_, _24557_);
  or (_24560_, _24559_, _24519_);
  and (_24561_, _24560_, _24556_);
  or (_24562_, _24561_, _24554_);
  or (_24563_, _24032_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24564_, _24533_, _24514_);
  and (_24565_, _24564_, _24563_);
  and (_24566_, _24565_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24567_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_24568_, _24567_);
  nand (_24569_, _24507_, _23973_);
  and (_24570_, _24569_, _24568_);
  not (_24571_, _24570_);
  or (_24572_, _24571_, _24566_);
  and (_24573_, _24553_, _24551_);
  nand (_24574_, _24560_, _24556_);
  or (_24575_, _24574_, _24573_);
  nand (_24576_, _24575_, _24562_);
  or (_24577_, _24576_, _24572_);
  nand (_24578_, _24577_, _24562_);
  nand (_24579_, _24578_, _24549_);
  and (_24580_, _24579_, _24546_);
  and (_24581_, _24517_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24582_, _24581_);
  nand (_24583_, _24507_, _24101_);
  nor (_24584_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_24585_, _24584_);
  and (_24586_, _24585_, _24583_);
  nand (_24587_, _24586_, _24582_);
  or (_24588_, _24586_, _24582_);
  nand (_24589_, _24588_, _24587_);
  nand (_24590_, _24531_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24591_, _24550_, _24216_);
  nor (_24592_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_24593_, _24592_);
  and (_24594_, _24593_, _24591_);
  nand (_24595_, _24594_, _24590_);
  and (_24596_, _24555_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24597_, _24550_, _24200_);
  nor (_24598_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_24599_, _24598_);
  nand (_24600_, _24599_, _24597_);
  and (_24601_, _24600_, _24596_);
  or (_24602_, _24594_, _24590_);
  nand (_24603_, _24602_, _24595_);
  or (_24604_, _24603_, _24601_);
  and (_24605_, _24604_, _24595_);
  or (_24606_, _24605_, _24589_);
  nand (_24607_, _24606_, _24587_);
  not (_24608_, _24566_);
  or (_24609_, _24570_, _24608_);
  and (_24610_, _24609_, _24572_);
  not (_24611_, _24610_);
  nor (_24612_, _24576_, _24611_);
  and (_24613_, _24612_, _24549_);
  nand (_24614_, _24613_, _24607_);
  nand (_24615_, _24614_, _24580_);
  not (_24616_, _24049_);
  and (_24617_, _23990_, _24616_);
  nor (_24618_, _24617_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24619_, _24537_, _24523_);
  or (_24620_, _24535_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24621_, _23990_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_24622_, _24621_, _24620_);
  nor (_24623_, _24622_, _24559_);
  nand (_24624_, _24623_, _24619_);
  and (_24625_, _24624_, _24519_);
  nor (_24626_, _24625_, _24618_);
  nor (_24627_, _24565_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24628_, _24622_, _24519_);
  nor (_24629_, _24628_, _24627_);
  not (_24630_, _24629_);
  and (_24631_, _24630_, _24626_);
  and (_24632_, _24631_, _24615_);
  nor (_24633_, _24632_, _24512_);
  not (_24634_, _24633_);
  not (_24635_, _24548_);
  and (_24636_, _24577_, _24562_);
  nand (_24637_, _24612_, _24607_);
  and (_24638_, _24637_, _24636_);
  or (_24639_, _24638_, _24635_);
  and (_24640_, _24639_, _24540_);
  nand (_24641_, _24640_, _24543_);
  or (_24642_, _24640_, _24543_);
  nand (_24643_, _24642_, _24641_);
  nand (_24644_, _24643_, _24632_);
  and (_24645_, _24644_, _24634_);
  and (_24646_, _24645_, _24629_);
  nor (_24647_, _24645_, _24629_);
  and (_24648_, _24638_, _24635_);
  not (_24649_, _24648_);
  nand (_24650_, _24649_, _24639_);
  nand (_24651_, _24650_, _24632_);
  nor (_24652_, _24632_, _24530_);
  not (_24653_, _24652_);
  and (_24654_, _24653_, _24651_);
  and (_24655_, _24654_, _24541_);
  nor (_24656_, _24655_, _24647_);
  or (_24657_, _24656_, _24646_);
  nor (_24658_, _24647_, _24646_);
  not (_24659_, _24655_);
  or (_24660_, _24654_, _24541_);
  and (_24661_, _24660_, _24659_);
  and (_24662_, _24661_, _24658_);
  not (_24663_, _24632_);
  nand (_24664_, _24610_, _24607_);
  and (_24665_, _24664_, _24572_);
  and (_24666_, _24576_, _24665_);
  nor (_24667_, _24576_, _24665_);
  nor (_24668_, _24667_, _24666_);
  nor (_24669_, _24668_, _24663_);
  nor (_24670_, _24632_, _24573_);
  nor (_24671_, _24670_, _24669_);
  and (_24672_, _24671_, _24539_);
  not (_24673_, _24672_);
  nor (_24674_, _24671_, _24539_);
  nor (_24675_, _24632_, _24571_);
  nor (_24676_, _24610_, _24607_);
  not (_24677_, _24676_);
  and (_24678_, _24677_, _24664_);
  and (_24679_, _24678_, _24632_);
  or (_24680_, _24679_, _24675_);
  and (_24681_, _24680_, _24574_);
  not (_24682_, _24681_);
  and (_24683_, _24605_, _24589_);
  not (_24684_, _24683_);
  and (_24685_, _24684_, _24606_);
  or (_24686_, _24685_, _24663_);
  or (_24687_, _24632_, _24586_);
  and (_24688_, _24687_, _24686_);
  nor (_24689_, _24688_, _24608_);
  or (_24690_, _24632_, _24600_);
  not (_24691_, _24596_);
  and (_24694_, _24600_, _24691_);
  nor (_24705_, _24600_, _24691_);
  nor (_24716_, _24705_, _24694_);
  nand (_24727_, _24632_, _24716_);
  nand (_24734_, _24727_, _24690_);
  nand (_24742_, _24734_, _24590_);
  or (_24753_, _24734_, _24590_);
  nand (_24764_, _24753_, _24742_);
  nor (_24775_, _24507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and (_24786_, _24507_, _24253_);
  nor (_24797_, _24786_, _24775_);
  nor (_24808_, _24797_, _24691_);
  or (_24819_, _24808_, _24764_);
  and (_24830_, _24819_, _24742_);
  or (_24841_, _24632_, _24594_);
  and (_24852_, _24603_, _24601_);
  not (_24863_, _24852_);
  and (_24874_, _24863_, _24604_);
  or (_24885_, _24874_, _24663_);
  and (_24896_, _24885_, _24841_);
  nand (_24906_, _24896_, _24582_);
  or (_24907_, _24896_, _24582_);
  nand (_24908_, _24907_, _24906_);
  or (_24909_, _24908_, _24830_);
  and (_24910_, _24688_, _24608_);
  not (_24911_, _24910_);
  and (_24912_, _24911_, _24906_);
  and (_24913_, _24912_, _24909_);
  nor (_24914_, _24913_, _24689_);
  nor (_24915_, _24680_, _24574_);
  nor (_24916_, _24915_, _24681_);
  nand (_24917_, _24916_, _24914_);
  and (_24918_, _24917_, _24682_);
  or (_24919_, _24918_, _24674_);
  nand (_24920_, _24919_, _24673_);
  nand (_24921_, _24920_, _24662_);
  nand (_24922_, _24921_, _24657_);
  and (_24923_, _24922_, _24626_);
  nor (_24924_, _24923_, _24645_);
  and (_24925_, _24920_, _24661_);
  or (_24926_, _24925_, _24655_);
  or (_24927_, _24926_, _24658_);
  nand (_24928_, _24926_, _24658_);
  and (_24929_, _24928_, _24927_);
  and (_24930_, _24929_, _24923_);
  or (_24931_, _24930_, _24924_);
  and (_01001_, _24931_, _27355_);
  and (_03039_, _24923_, _27355_);
  and (_03049_, _24632_, _27355_);
  and (_03068_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _27355_);
  and (_03084_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _27355_);
  and (_03100_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _27355_);
  or (_24932_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24933_, _24488_, rst);
  and (_03108_, _24933_, _24932_);
  nand (_24934_, _24923_, _24596_);
  and (_24935_, _24934_, _24797_);
  nor (_24936_, _24934_, _24797_);
  or (_24937_, _24936_, _24935_);
  and (_03117_, _24937_, _27355_);
  nand (_24938_, _24922_, _24626_);
  and (_24939_, _24808_, _24764_);
  not (_24940_, _24939_);
  and (_24941_, _24940_, _24819_);
  or (_24942_, _24941_, _24938_);
  or (_24943_, _24923_, _24734_);
  and (_24944_, _24943_, _24942_);
  and (_03125_, _24944_, _27355_);
  not (_24945_, _24909_);
  and (_24946_, _24908_, _24830_);
  nor (_24947_, _24946_, _24945_);
  or (_24948_, _24947_, _24938_);
  or (_24949_, _24923_, _24896_);
  and (_24950_, _24949_, _24948_);
  and (_03132_, _24950_, _27355_);
  or (_24951_, _24910_, _24689_);
  and (_24952_, _24909_, _24906_);
  nor (_24953_, _24952_, _24951_);
  and (_24954_, _24952_, _24951_);
  nor (_24955_, _24954_, _24953_);
  or (_24956_, _24955_, _24938_);
  or (_24957_, _24923_, _24688_);
  and (_24958_, _24957_, _24956_);
  and (_03141_, _24958_, _27355_);
  or (_24959_, _24916_, _24914_);
  and (_24960_, _24959_, _24917_);
  or (_24961_, _24960_, _24938_);
  or (_24962_, _24923_, _24680_);
  and (_24963_, _24962_, _24961_);
  and (_03149_, _24963_, _27355_);
  or (_24964_, _24674_, _24672_);
  nand (_24965_, _24964_, _24918_);
  or (_24966_, _24964_, _24918_);
  and (_24967_, _24966_, _24965_);
  or (_24968_, _24967_, _24938_);
  or (_24969_, _24923_, _24671_);
  and (_24970_, _24969_, _24968_);
  and (_03158_, _24970_, _27355_);
  nor (_24971_, _24920_, _24661_);
  or (_24972_, _24971_, _24925_);
  and (_24973_, _24972_, _24923_);
  nor (_24974_, _24923_, _24654_);
  or (_24975_, _24974_, _24973_);
  nor (_03166_, _24975_, rst);
  not (_24976_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_24977_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _23914_);
  and (_24978_, _24977_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24979_, _24978_, _24976_);
  and (_24980_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24981_, _24980_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24982_, _24980_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24983_, _24982_, _24981_);
  and (_24984_, _24983_, _24979_);
  not (_24985_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_24986_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _23914_);
  and (_24988_, _24986_, _24976_);
  and (_24990_, _24988_, _24985_);
  and (_24992_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24994_, _24992_, _24984_);
  not (_24996_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_24998_, _24977_, _24996_);
  and (_25000_, _24998_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_25002_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_25004_, _24998_, _24976_);
  and (_25006_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or (_25008_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_25010_, _25008_, _23914_);
  nor (_25012_, _25010_, _24977_);
  and (_25014_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_25016_, _25014_, _25006_);
  nor (_25018_, _25016_, _25002_);
  and (_25020_, _25018_, _24994_);
  and (_25022_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_25024_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_25026_, _25024_, _24980_);
  and (_25028_, _25026_, _24979_);
  nor (_25030_, _25028_, _25022_);
  and (_25032_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_25034_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_25036_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_25038_, _25036_, _25034_);
  nor (_25040_, _25038_, _25032_);
  and (_25042_, _25040_, _25030_);
  and (_25043_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_25044_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_25045_, _25044_, _25043_);
  not (_25046_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_25047_, _24979_, _25046_);
  not (_25048_, _25047_);
  and (_25049_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_25050_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_25051_, _25050_, _25049_);
  and (_25052_, _25051_, _25048_);
  and (_25053_, _25052_, _25045_);
  and (_25054_, _25053_, _25042_);
  and (_25055_, _25054_, _25020_);
  and (_25056_, _24981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_25057_, _25056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_25058_, _25057_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_25059_, _25058_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_25060_, _25059_);
  not (_25061_, _24979_);
  nor (_25062_, _25058_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_25063_, _25062_, _25061_);
  and (_25064_, _25063_, _25060_);
  not (_25065_, _25064_);
  and (_25066_, _24978_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_25067_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_25068_, _25067_, _25066_);
  and (_25069_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_25070_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_25071_, _25070_, _25069_);
  and (_25072_, _25071_, _25068_);
  and (_25073_, _25072_, _25065_);
  nor (_25074_, _25057_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_25075_, _25074_);
  nor (_25076_, _25058_, _25061_);
  and (_25077_, _25076_, _25075_);
  not (_25078_, _25077_);
  and (_25079_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_25080_, _25079_, _25066_);
  and (_25081_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_25082_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_25083_, _25082_, _25081_);
  and (_25084_, _25083_, _25080_);
  and (_25085_, _25084_, _25078_);
  nor (_25086_, _25085_, _25073_);
  not (_25087_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_25088_, _25059_, _25087_);
  and (_25089_, _25059_, _25087_);
  nor (_25090_, _25089_, _25088_);
  nor (_25091_, _25090_, _25061_);
  not (_25092_, _25091_);
  and (_25093_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_25094_, _25093_);
  not (_25095_, _25066_);
  and (_25096_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_25097_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_25098_, _25097_, _25096_);
  and (_25099_, _25098_, _25095_);
  and (_25100_, _25099_, _25094_);
  and (_25101_, _25100_, _25092_);
  not (_25102_, _25101_);
  and (_25103_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_25104_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_25105_, _25104_, _25103_);
  not (_25106_, _25056_);
  nor (_25107_, _24981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_25108_, _25107_, _25061_);
  and (_25109_, _25108_, _25106_);
  and (_25110_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_25111_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_25112_, _25111_, _25110_);
  not (_25113_, _25112_);
  nor (_25114_, _25113_, _25109_);
  and (_25115_, _25114_, _25105_);
  not (_25116_, _25115_);
  and (_25117_, _25000_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_25118_, _25117_, _25066_);
  nor (_25119_, _25056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_25120_, _25119_, _25061_);
  nor (_25121_, _25120_, _25057_);
  and (_25122_, _25004_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_25123_, _25122_, _25121_);
  and (_25124_, _25123_, _25118_);
  and (_25125_, _25012_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_25126_, _24990_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_25127_, _25126_, _25125_);
  and (_25128_, _25127_, _25124_);
  nor (_25129_, _25128_, _25116_);
  and (_25130_, _25129_, _25102_);
  and (_25131_, _25130_, _25086_);
  nand (_25132_, _25131_, _25055_);
  and (_25133_, _24931_, _24487_);
  and (_25134_, _24390_, _23920_);
  nor (_25135_, _23973_, _24055_);
  and (_25136_, _23973_, _24055_);
  nor (_25137_, _25136_, _25135_);
  nor (_25138_, _24101_, _24018_);
  and (_25139_, _24101_, _24018_);
  nor (_25140_, _25139_, _25138_);
  and (_25141_, _24216_, _24515_);
  nor (_25142_, _24216_, _24515_);
  nor (_25143_, _25142_, _25141_);
  not (_25144_, _25143_);
  and (_25145_, _24200_, _24032_);
  not (_25146_, _24082_);
  nor (_25147_, _24253_, _25146_);
  nor (_25148_, _24200_, _24032_);
  nor (_25149_, _25148_, _25145_);
  and (_25150_, _25149_, _25147_);
  nor (_25151_, _25150_, _25145_);
  nor (_25152_, _25151_, _25144_);
  nor (_25153_, _25152_, _25141_);
  nor (_25155_, _25153_, _25140_);
  and (_25164_, _25153_, _25140_);
  nor (_25165_, _25164_, _25155_);
  nor (_25166_, _23960_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_25167_, _25166_);
  nor (_25168_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_25169_, _25168_, _23958_);
  and (_25170_, _25169_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_25171_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25172_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25171_);
  nand (_25173_, _25172_, _23995_);
  not (_25174_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_25175_, _25174_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_25176_, _25175_, _24040_);
  and (_25177_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_25178_, _25177_, _23978_);
  and (_25179_, _25178_, _25176_);
  and (_25180_, _25179_, _25173_);
  nand (_25181_, _25180_, _25170_);
  not (_25182_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_25183_, _25168_, _24073_);
  and (_25184_, _25183_, _25182_);
  nand (_25185_, _25177_, _24009_);
  nand (_25186_, _25175_, _24059_);
  nand (_25187_, _25172_, _24023_);
  and (_25188_, _25187_, _25186_);
  and (_25189_, _25188_, _25185_);
  nand (_25190_, _25189_, _25184_);
  nand (_25191_, _25190_, _25181_);
  nand (_25192_, _25191_, _23960_);
  and (_25193_, _25192_, _25167_);
  and (_25194_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_25195_, _25194_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_25196_, _25195_);
  and (_25197_, _25196_, _25193_);
  and (_25198_, _25196_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_25199_, _25198_, _25197_);
  and (_25200_, _24253_, _25146_);
  nor (_25201_, _25200_, _25147_);
  not (_25202_, _25201_);
  nor (_25203_, _25202_, _25199_);
  and (_25204_, _25203_, _25149_);
  and (_25205_, _25151_, _25144_);
  nor (_25206_, _25205_, _25152_);
  and (_25207_, _25206_, _25204_);
  not (_25208_, _25207_);
  nor (_25209_, _25208_, _25165_);
  nor (_25210_, _25153_, _25139_);
  or (_25211_, _25210_, _25138_);
  or (_25212_, _25211_, _25209_);
  and (_25213_, _25212_, _25137_);
  and (_25214_, _24120_, _24535_);
  nor (_25215_, _24120_, _24535_);
  nor (_25216_, _25215_, _25214_);
  and (_25217_, _25216_, _25135_);
  nor (_25218_, _25216_, _25135_);
  nor (_25219_, _25218_, _25217_);
  and (_25220_, _25219_, _25213_);
  nor (_25221_, _24141_, _24616_);
  and (_25222_, _24141_, _24616_);
  nor (_25223_, _25222_, _25221_);
  not (_25224_, _25223_);
  nor (_25225_, _25217_, _25214_);
  nor (_25226_, _25225_, _25224_);
  and (_25227_, _25225_, _25224_);
  nor (_25228_, _25227_, _25226_);
  and (_25229_, _25228_, _25220_);
  nor (_25230_, _25226_, _25221_);
  not (_25231_, _25230_);
  nor (_25232_, _25231_, _25229_);
  nor (_25233_, _24172_, _23990_);
  and (_25234_, _24172_, _23990_);
  nor (_25235_, _25234_, _25233_);
  not (_25236_, _25235_);
  nor (_25237_, _25236_, _25232_);
  not (_25238_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_25239_, _24468_, _25238_);
  and (_25240_, _25239_, _23919_);
  nand (_25241_, _25236_, _25232_);
  nand (_25242_, _25241_, _25240_);
  nor (_25243_, _25242_, _25237_);
  not (_25244_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_25245_, _23915_, _25244_);
  and (_25246_, _25245_, _23919_);
  not (_25247_, _25246_);
  nor (_25248_, _24141_, _24049_);
  and (_25249_, _24120_, _24004_);
  and (_25250_, _23973_, _24520_);
  nor (_25251_, _25250_, _25216_);
  nor (_25252_, _25251_, _25249_);
  nor (_25253_, _25252_, _25223_);
  nor (_25254_, _25253_, _25248_);
  and (_25255_, _25252_, _25223_);
  nor (_25256_, _25255_, _25253_);
  not (_25257_, _25256_);
  and (_25258_, _25250_, _25216_);
  nor (_25259_, _25258_, _25251_);
  not (_25260_, _25259_);
  not (_25266_, _25137_);
  not (_25277_, _25140_);
  and (_25288_, _24253_, _24082_);
  nor (_25299_, _25288_, _25149_);
  not (_25310_, _24032_);
  and (_25321_, _24200_, _25310_);
  nor (_25323_, _25321_, _25299_);
  nor (_25324_, _25323_, _25143_);
  and (_25325_, _24216_, _24068_);
  nor (_25326_, _25325_, _25324_);
  nor (_25327_, _25326_, _25277_);
  and (_25328_, _25326_, _25277_);
  nor (_25329_, _25328_, _25327_);
  and (_25330_, _25323_, _25143_);
  nor (_25331_, _25330_, _25324_);
  not (_25332_, _25331_);
  and (_25333_, _25288_, _25149_);
  nor (_25334_, _25333_, _25299_);
  not (_25335_, _25334_);
  nor (_25336_, _25201_, _25199_);
  and (_25337_, _25336_, _25335_);
  and (_25338_, _25337_, _25332_);
  and (_25339_, _25338_, _25329_);
  or (_25340_, _24101_, _24533_);
  and (_25341_, _24101_, _24533_);
  or (_25342_, _25326_, _25341_);
  and (_25343_, _25342_, _25340_);
  or (_25344_, _25343_, _25339_);
  and (_25345_, _25344_, _25266_);
  and (_25346_, _25345_, _25260_);
  and (_25347_, _25346_, _25257_);
  nor (_25348_, _25347_, _25254_);
  nor (_25349_, _25348_, _25235_);
  and (_25350_, _25348_, _25235_);
  nor (_25351_, _25350_, _25349_);
  nor (_25352_, _25351_, _25247_);
  and (_25353_, _23918_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_25354_, _25353_, _25245_);
  not (_25355_, _24200_);
  nor (_25356_, _24253_, _25355_);
  and (_25357_, _25356_, _24216_);
  and (_25358_, _25357_, _24102_);
  and (_25359_, _25358_, _23974_);
  and (_25360_, _25359_, _24120_);
  and (_25361_, _25360_, _24143_);
  and (_25362_, _25361_, _25199_);
  not (_25363_, _25199_);
  not (_25364_, _24120_);
  and (_25365_, _24141_, _25364_);
  nor (_25366_, _24216_, _24200_);
  and (_25367_, _25366_, _24253_);
  and (_25368_, _25367_, _24101_);
  and (_25369_, _25368_, _23973_);
  and (_25370_, _25369_, _25365_);
  and (_25371_, _25370_, _25363_);
  nor (_25372_, _25371_, _25362_);
  and (_25373_, _25372_, _24172_);
  nor (_25374_, _25372_, _24172_);
  nor (_25375_, _25374_, _25373_);
  and (_25376_, _25375_, _25354_);
  not (_25377_, _23990_);
  nor (_25378_, _25199_, _25377_);
  not (_25379_, _25378_);
  and (_25380_, _25199_, _24172_);
  and (_25381_, _25353_, _23916_);
  not (_25382_, _25381_);
  nor (_25383_, _25382_, _25380_);
  and (_25384_, _25383_, _25379_);
  nor (_25385_, _25384_, _25376_);
  not (_25386_, _25365_);
  and (_25390_, _25239_, _24482_);
  nor (_25394_, _25366_, _24101_);
  and (_25395_, _25394_, _25390_);
  and (_25396_, _25395_, _23974_);
  nor (_25397_, _25396_, _25386_);
  nor (_25398_, _25365_, _24172_);
  nor (_25399_, _25398_, _25395_);
  and (_25400_, _25399_, _25199_);
  nor (_25401_, _25400_, _25397_);
  nand (_25402_, _25401_, _24278_);
  or (_25403_, _25401_, _24278_);
  and (_25404_, _25403_, _25390_);
  and (_25405_, _25404_, _25402_);
  and (_25406_, _25353_, _25239_);
  and (_25407_, _25406_, _25363_);
  not (_25408_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_25409_, _23918_, _25408_);
  and (_25410_, _25409_, _25239_);
  not (_25411_, _25410_);
  nor (_25412_, _25411_, _25234_);
  and (_25413_, _25409_, _24469_);
  and (_25414_, _25413_, _25235_);
  nor (_25415_, _25414_, _25412_);
  and (_25416_, _24482_, _23916_);
  and (_25417_, _25416_, _25233_);
  and (_25418_, _25245_, _24482_);
  and (_25419_, _25418_, _24172_);
  nor (_25420_, _25419_, _25417_);
  and (_25421_, _25353_, _24469_);
  and (_25422_, _25421_, _24254_);
  and (_25423_, _24469_, _23919_);
  not (_25424_, _25423_);
  nor (_25425_, _25424_, _24172_);
  and (_25426_, _25409_, _23915_);
  not (_25427_, _25426_);
  nor (_25428_, _25427_, _24141_);
  or (_25429_, _25428_, _25425_);
  nor (_25430_, _25429_, _25422_);
  and (_25431_, _25430_, _25420_);
  nand (_25432_, _25431_, _25415_);
  or (_25433_, _25432_, _25407_);
  nor (_25434_, _25433_, _25405_);
  nand (_25435_, _25434_, _25385_);
  or (_25437_, _25435_, _25352_);
  or (_25438_, _25437_, _25243_);
  or (_25440_, _25438_, _25134_);
  or (_25441_, _25440_, _25133_);
  or (_25443_, _25441_, _25132_);
  not (_25444_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_25446_, \oc8051_top_1.oc8051_decoder1.wr , _23914_);
  not (_25447_, _25446_);
  nor (_25449_, _25447_, _24988_);
  and (_25450_, _25449_, _25444_);
  not (_25452_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_25453_, _25132_, _25452_);
  and (_25455_, _25453_, _25450_);
  and (_25456_, _25455_, _25443_);
  nor (_25458_, _25449_, _25452_);
  not (_25459_, _25240_);
  nor (_25461_, _25237_, _25233_);
  nor (_25462_, _25461_, _25459_);
  not (_25464_, _25462_);
  and (_25465_, _24172_, _25377_);
  nor (_25466_, _25465_, _25349_);
  nor (_25467_, _25466_, _25247_);
  and (_25468_, _25397_, _25199_);
  nor (_25469_, _25468_, _25380_);
  not (_25470_, _25390_);
  not (_25471_, _25397_);
  nor (_25472_, _25199_, _24172_);
  and (_25473_, _25472_, _25471_);
  nor (_25474_, _25473_, _25470_);
  and (_25475_, _25474_, _25469_);
  and (_25476_, _25195_, _25193_);
  and (_25477_, _25409_, _25245_);
  and (_25478_, _25416_, _25193_);
  nor (_25479_, _25478_, _25477_);
  nor (_25480_, _25479_, _25476_);
  nor (_25481_, _25199_, _25193_);
  and (_25482_, _25481_, _25421_);
  and (_25483_, _25418_, _25199_);
  or (_25484_, _25483_, _25482_);
  nor (_25491_, _25198_, _25193_);
  not (_25496_, _25413_);
  nor (_25497_, _25496_, _25197_);
  nor (_25498_, _25497_, _25410_);
  nor (_25499_, _25498_, _25491_);
  nor (_25500_, _25424_, _25199_);
  and (_25501_, _25409_, _23916_);
  not (_25502_, _25501_);
  nor (_25503_, _25502_, _24172_);
  and (_25504_, _25406_, _24254_);
  or (_25505_, _25504_, _25395_);
  or (_25506_, _25505_, _25503_);
  or (_25507_, _25506_, _25500_);
  or (_25508_, _25507_, _25499_);
  or (_25509_, _25508_, _25484_);
  or (_25510_, _25509_, _25480_);
  nor (_25511_, _25510_, _25475_);
  not (_25512_, _25511_);
  nor (_25513_, _25512_, _25467_);
  and (_25514_, _25513_, _25464_);
  not (_25515_, _25020_);
  nor (_25516_, _25053_, _25042_);
  and (_25517_, _25516_, _25515_);
  and (_25518_, _25517_, _25131_);
  nand (_25519_, _25518_, _25514_);
  or (_25520_, _25518_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_25521_, _25449_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_25522_, _25521_, _25520_);
  and (_25523_, _25522_, _25519_);
  or (_25524_, _25523_, _25458_);
  or (_25525_, _25524_, _25456_);
  and (_06524_, _25525_, _27355_);
  nand (_25526_, _24937_, _24487_);
  and (_25527_, _24448_, _23920_);
  and (_25528_, _25202_, _25199_);
  nor (_25529_, _25528_, _25203_);
  not (_25530_, _25529_);
  nor (_25531_, _25246_, _25240_);
  nor (_25532_, _25531_, _25530_);
  nor (_25533_, _25502_, _25199_);
  not (_25534_, _25533_);
  and (_25535_, _25413_, _25201_);
  not (_25536_, _25535_);
  nor (_25537_, _25411_, _25200_);
  not (_25538_, _25537_);
  and (_25539_, _25416_, _25147_);
  and (_25540_, _25418_, _24253_);
  nor (_25541_, _25540_, _25539_);
  and (_25542_, _25541_, _25538_);
  and (_25543_, _25542_, _25536_);
  and (_25544_, _25381_, _24082_);
  and (_25545_, _25354_, _24253_);
  nor (_25546_, _25545_, _25544_);
  and (_25547_, _25477_, _24278_);
  not (_25548_, _25547_);
  and (_25549_, _25353_, _25238_);
  and (_25550_, _25549_, _24200_);
  nor (_25551_, _25423_, _25390_);
  nor (_25552_, _25551_, _24253_);
  nor (_25553_, _25552_, _25550_);
  and (_25554_, _25553_, _25548_);
  and (_25555_, _25554_, _25546_);
  and (_25556_, _25555_, _25543_);
  and (_25557_, _25556_, _25534_);
  not (_25558_, _25557_);
  nor (_25559_, _25558_, _25532_);
  not (_25560_, _25559_);
  nor (_25561_, _25560_, _25527_);
  and (_25562_, _25561_, _25526_);
  not (_25563_, _25562_);
  or (_25564_, _25563_, _25132_);
  not (_25565_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_25566_, _25132_, _25565_);
  and (_25570_, _25566_, _25450_);
  and (_25572_, _25570_, _25564_);
  nor (_25573_, _25449_, _25565_);
  not (_25574_, _25514_);
  or (_25575_, _25574_, _25132_);
  and (_25576_, _25566_, _25521_);
  and (_25577_, _25576_, _25575_);
  or (_25578_, _25577_, _25573_);
  or (_25579_, _25578_, _25572_);
  and (_08841_, _25579_, _27355_);
  nand (_25580_, _24944_, _24487_);
  nor (_25581_, _25394_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_25582_, _25581_, _24200_);
  nor (_25583_, _25581_, _24200_);
  nor (_25584_, _25583_, _25582_);
  nor (_25585_, _25584_, _25470_);
  not (_25595_, _25585_);
  nor (_25596_, _25427_, _24253_);
  and (_25597_, _25423_, _24200_);
  and (_25598_, _25549_, _24216_);
  or (_25599_, _25598_, _25597_);
  nor (_25600_, _25599_, _25596_);
  and (_25601_, _25413_, _25149_);
  nor (_25602_, _25411_, _25148_);
  not (_25603_, _25602_);
  and (_25604_, _25416_, _25145_);
  and (_25605_, _25418_, _25355_);
  nor (_25606_, _25605_, _25604_);
  nand (_25607_, _25606_, _25603_);
  nor (_25608_, _25607_, _25601_);
  and (_25609_, _25608_, _25600_);
  and (_25610_, _25609_, _25595_);
  nor (_25611_, _25149_, _25147_);
  or (_25612_, _25611_, _25150_);
  and (_25613_, _25612_, _25203_);
  nor (_25614_, _25612_, _25203_);
  or (_25615_, _25614_, _25613_);
  and (_25616_, _25615_, _25240_);
  nor (_25617_, _25336_, _25335_);
  nor (_25619_, _25617_, _25337_);
  nor (_25620_, _25619_, _25247_);
  nor (_25621_, _25620_, _25616_);
  and (_25623_, _25621_, _25610_);
  nand (_25624_, _24452_, _23920_);
  and (_25626_, _25381_, _24032_);
  not (_25627_, _25626_);
  and (_25628_, _24253_, _25355_);
  nor (_25630_, _25628_, _25356_);
  and (_25631_, _25630_, _25363_);
  or (_25632_, _25630_, _25363_);
  nand (_25633_, _25632_, _25354_);
  or (_25635_, _25633_, _25631_);
  and (_25636_, _25635_, _25627_);
  and (_25637_, _25636_, _25624_);
  and (_25638_, _25637_, _25623_);
  nand (_25639_, _25638_, _25580_);
  or (_25641_, _25639_, _25132_);
  not (_25642_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_25643_, _25132_, _25642_);
  and (_25644_, _25643_, _25450_);
  and (_25645_, _25644_, _25641_);
  nor (_25646_, _25449_, _25642_);
  nand (_25648_, _25131_, _25020_);
  not (_25649_, _25053_);
  and (_25650_, _25649_, _25042_);
  not (_25651_, _25650_);
  nor (_25652_, _25651_, _25648_);
  nand (_25653_, _25652_, _25514_);
  or (_25654_, _25652_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_25656_, _25654_, _25521_);
  and (_25657_, _25656_, _25653_);
  or (_25658_, _25657_, _25646_);
  or (_25659_, _25658_, _25645_);
  and (_08853_, _25659_, _27355_);
  nand (_25660_, _24456_, _23920_);
  nand (_25661_, _24950_, _24487_);
  and (_25662_, _25381_, _24515_);
  not (_25664_, _24216_);
  nand (_25665_, _25356_, _25199_);
  nand (_25666_, _25628_, _25363_);
  and (_25667_, _25666_, _25665_);
  nand (_25668_, _25667_, _25664_);
  or (_25669_, _25667_, _25664_);
  and (_25670_, _25669_, _25668_);
  and (_25671_, _25670_, _25354_);
  nor (_25672_, _25671_, _25662_);
  nor (_25674_, _25337_, _25332_);
  nor (_25675_, _25674_, _25338_);
  nor (_25676_, _25675_, _25247_);
  not (_25677_, _25676_);
  and (_25678_, _25549_, _24102_);
  and (_25679_, _25416_, _25141_);
  and (_25680_, _25418_, _25664_);
  nor (_25681_, _25680_, _25679_);
  nor (_25682_, _25411_, _25142_);
  and (_25684_, _25413_, _25143_);
  nor (_25685_, _25684_, _25682_);
  and (_25686_, _25423_, _24216_);
  and (_25687_, _25426_, _24200_);
  nor (_25688_, _25687_, _25686_);
  and (_25689_, _25688_, _25685_);
  nand (_25690_, _25689_, _25681_);
  nor (_25691_, _25690_, _25678_);
  and (_25692_, _25691_, _25677_);
  nor (_25693_, _25206_, _25204_);
  nor (_25694_, _25693_, _25459_);
  and (_25695_, _25694_, _25208_);
  nor (_25696_, _25583_, _25664_);
  and (_25697_, _25366_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_25698_, _25697_, _25696_);
  nor (_25699_, _25698_, _25470_);
  nor (_25700_, _25699_, _25695_);
  and (_25701_, _25700_, _25692_);
  and (_25702_, _25701_, _25672_);
  and (_25703_, _25702_, _25661_);
  and (_25704_, _25703_, _25660_);
  not (_25705_, _25704_);
  or (_25706_, _25705_, _25132_);
  not (_25707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_25708_, _25132_, _25707_);
  and (_25709_, _25708_, _25450_);
  and (_25710_, _25709_, _25706_);
  nor (_25711_, _25449_, _25707_);
  or (_25712_, _25516_, _25648_);
  and (_25713_, _25712_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_25714_, _25042_);
  and (_25715_, _25020_, _25053_);
  and (_25716_, _25715_, _25714_);
  not (_25717_, _25716_);
  nor (_25718_, _25717_, _25514_);
  nand (_25719_, _25020_, _25042_);
  nor (_25720_, _25719_, _25707_);
  or (_25721_, _25720_, _25718_);
  and (_25722_, _25721_, _25131_);
  or (_25723_, _25722_, _25713_);
  and (_25724_, _25723_, _25521_);
  or (_25725_, _25724_, _25711_);
  or (_25726_, _25725_, _25710_);
  and (_08864_, _25726_, _27355_);
  nand (_25727_, _24460_, _23920_);
  nand (_25728_, _24958_, _24487_);
  and (_25729_, _25381_, _24533_);
  nand (_25730_, _25357_, _25199_);
  nand (_25731_, _25367_, _25363_);
  nand (_25732_, _25731_, _25730_);
  and (_25733_, _25732_, _24102_);
  or (_25734_, _25732_, _24102_);
  nand (_25735_, _25734_, _25354_);
  nor (_25736_, _25735_, _25733_);
  nor (_25737_, _25736_, _25729_);
  not (_25738_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_25739_, _25366_, _25738_);
  nor (_25740_, _25739_, _24102_);
  or (_25741_, _25740_, _25470_);
  nor (_25742_, _25741_, _25394_);
  not (_25743_, _25742_);
  nor (_25744_, _25411_, _25139_);
  and (_25745_, _25413_, _25140_);
  nor (_25746_, _25745_, _25744_);
  and (_25747_, _25416_, _25138_);
  and (_25748_, _25418_, _24101_);
  nor (_25749_, _25748_, _25747_);
  and (_25750_, _25549_, _23974_);
  not (_25751_, _25750_);
  nor (_25752_, _25424_, _24101_);
  and (_25753_, _25426_, _24216_);
  nor (_25754_, _25753_, _25752_);
  and (_25755_, _25754_, _25751_);
  and (_25756_, _25755_, _25749_);
  and (_25757_, _25756_, _25746_);
  and (_25758_, _25757_, _25743_);
  nor (_25759_, _25338_, _25329_);
  nor (_25760_, _25759_, _25339_);
  nor (_25761_, _25760_, _25247_);
  and (_25762_, _25208_, _25165_);
  or (_25763_, _25762_, _25459_);
  nor (_25764_, _25763_, _25209_);
  nor (_25765_, _25764_, _25761_);
  and (_25766_, _25765_, _25758_);
  and (_25767_, _25766_, _25737_);
  and (_25768_, _25767_, _25728_);
  and (_25769_, _25768_, _25727_);
  not (_25770_, _25769_);
  or (_25771_, _25770_, _25132_);
  not (_25772_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_25773_, _25132_, _25772_);
  and (_25774_, _25773_, _25450_);
  and (_25775_, _25774_, _25771_);
  nor (_25776_, _25449_, _25772_);
  and (_25777_, _25648_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_25778_, _25516_, _25020_);
  and (_25779_, _25778_, _25574_);
  or (_25780_, _25516_, _25515_);
  nor (_25781_, _25780_, _25772_);
  or (_25782_, _25781_, _25779_);
  and (_25783_, _25782_, _25131_);
  or (_25784_, _25783_, _25777_);
  and (_25785_, _25784_, _25521_);
  or (_25786_, _25785_, _25776_);
  or (_25787_, _25786_, _25775_);
  and (_08876_, _25787_, _27355_);
  and (_25788_, _24963_, _24487_);
  and (_25789_, _24463_, _23920_);
  nor (_25790_, _25344_, _25137_);
  and (_25791_, _25344_, _25137_);
  nor (_25792_, _25791_, _25790_);
  and (_25793_, _25792_, _25246_);
  or (_25794_, _25212_, _25137_);
  nor (_25795_, _25459_, _25213_);
  and (_25796_, _25795_, _25794_);
  nor (_25797_, _25199_, _24055_);
  and (_25798_, _25199_, _23974_);
  nor (_25799_, _25798_, _25797_);
  nor (_25800_, _25799_, _25382_);
  and (_25801_, _25358_, _25199_);
  and (_25802_, _25368_, _25363_);
  nor (_25803_, _25802_, _25801_);
  and (_25804_, _25803_, _23973_);
  nor (_25805_, _25803_, _23973_);
  nor (_25806_, _25805_, _25804_);
  and (_25807_, _25806_, _25354_);
  nor (_25808_, _25807_, _25800_);
  or (_25809_, _25395_, _23974_);
  nor (_25810_, _25424_, _23973_);
  nor (_25811_, _25396_, _25470_);
  or (_25812_, _25811_, _25810_);
  and (_25813_, _25812_, _25809_);
  and (_25814_, _25413_, _25137_);
  and (_25815_, _25416_, _25135_);
  nor (_25816_, _25411_, _25136_);
  and (_25817_, _25418_, _23973_);
  or (_25818_, _25817_, _25816_);
  or (_25819_, _25818_, _25815_);
  nor (_25820_, _25819_, _25814_);
  and (_25821_, _25549_, _24120_);
  nor (_25822_, _25427_, _24101_);
  nor (_25823_, _25822_, _25821_);
  nand (_25824_, _25823_, _25820_);
  nor (_25825_, _25824_, _25813_);
  nand (_25826_, _25825_, _25808_);
  or (_25827_, _25826_, _25796_);
  or (_25828_, _25827_, _25793_);
  or (_25829_, _25828_, _25789_);
  or (_25830_, _25829_, _25788_);
  or (_25831_, _25830_, _25132_);
  not (_25832_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_25833_, _25132_, _25832_);
  and (_25834_, _25833_, _25450_);
  and (_25835_, _25834_, _25831_);
  nor (_25836_, _25449_, _25832_);
  not (_25837_, _25131_);
  and (_25838_, _25054_, _25515_);
  nor (_25839_, _25054_, _25515_);
  nor (_25840_, _25839_, _25838_);
  or (_25841_, _25840_, _25837_);
  and (_25842_, _25841_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_25843_, _25838_, _25574_);
  and (_25844_, _25839_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_25845_, _25844_, _25843_);
  and (_25846_, _25845_, _25131_);
  or (_25847_, _25846_, _25842_);
  and (_25848_, _25847_, _25521_);
  or (_25849_, _25848_, _25836_);
  or (_25850_, _25849_, _25835_);
  and (_08887_, _25850_, _27355_);
  and (_25851_, _24970_, _24487_);
  and (_25852_, _24465_, _23920_);
  or (_25853_, _25219_, _25213_);
  nor (_25854_, _25459_, _25220_);
  and (_25855_, _25854_, _25853_);
  nor (_25856_, _25345_, _25260_);
  nor (_25857_, _25856_, _25346_);
  nor (_25858_, _25857_, _25247_);
  nor (_25859_, _25199_, _24004_);
  and (_25860_, _25199_, _24120_);
  nor (_25861_, _25860_, _25859_);
  nor (_25862_, _25861_, _25382_);
  and (_25863_, _25359_, _25199_);
  and (_25864_, _25369_, _25363_);
  nor (_25865_, _25864_, _25863_);
  and (_25866_, _25865_, _25364_);
  not (_25867_, _25354_);
  nor (_25868_, _25865_, _25364_);
  or (_25869_, _25868_, _25867_);
  nor (_25870_, _25869_, _25866_);
  nor (_25871_, _25870_, _25862_);
  nor (_25872_, _25396_, _24120_);
  not (_25873_, _25400_);
  and (_25874_, _25873_, _25872_);
  or (_25875_, _25400_, _25396_);
  and (_25876_, _25875_, _24120_);
  or (_25877_, _25876_, _25874_);
  and (_25878_, _25877_, _25390_);
  and (_25879_, _25413_, _25216_);
  nor (_25880_, _25411_, _25215_);
  not (_25881_, _25880_);
  and (_25882_, _25416_, _25214_);
  and (_25883_, _25418_, _25364_);
  nor (_25884_, _25883_, _25882_);
  nand (_25885_, _25884_, _25881_);
  nor (_25886_, _25885_, _25879_);
  and (_25887_, _25549_, _24143_);
  and (_25888_, _25423_, _24120_);
  nor (_25889_, _25427_, _23973_);
  or (_25890_, _25889_, _25888_);
  nor (_25891_, _25890_, _25887_);
  nand (_25892_, _25891_, _25886_);
  nor (_25893_, _25892_, _25878_);
  nand (_25894_, _25893_, _25871_);
  or (_25895_, _25894_, _25858_);
  or (_25896_, _25895_, _25855_);
  or (_25897_, _25896_, _25852_);
  or (_25898_, _25897_, _25851_);
  or (_25899_, _25898_, _25132_);
  not (_25900_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_25901_, _25132_, _25900_);
  and (_25902_, _25901_, _25450_);
  and (_25903_, _25902_, _25899_);
  nor (_25904_, _25449_, _25900_);
  and (_25905_, _25650_, _25515_);
  and (_25906_, _25905_, _25131_);
  nand (_25907_, _25906_, _25514_);
  or (_25908_, _25906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_25909_, _25908_, _25521_);
  and (_25910_, _25909_, _25907_);
  or (_25911_, _25910_, _25904_);
  or (_25912_, _25911_, _25903_);
  and (_08898_, _25912_, _27355_);
  not (_25913_, _24487_);
  or (_25914_, _24975_, _25913_);
  not (_25915_, _23920_);
  or (_25916_, _24467_, _25915_);
  nor (_25917_, _25346_, _25257_);
  nor (_25918_, _25917_, _25347_);
  nor (_25919_, _25918_, _25247_);
  not (_25920_, _25919_);
  nor (_25921_, _25228_, _25220_);
  not (_25922_, _25921_);
  nor (_25923_, _25459_, _25229_);
  and (_25924_, _25923_, _25922_);
  and (_25925_, _25199_, _24143_);
  nor (_25926_, _25199_, _24616_);
  or (_25927_, _25926_, _25925_);
  and (_25928_, _25927_, _25381_);
  or (_25929_, _25199_, _25364_);
  or (_25930_, _25864_, _25360_);
  and (_25931_, _25930_, _25929_);
  nor (_25932_, _25931_, _24143_);
  and (_25933_, _25931_, _24143_);
  or (_25934_, _25933_, _25867_);
  nor (_25935_, _25934_, _25932_);
  nor (_25936_, _25935_, _25928_);
  nor (_25937_, _25874_, _24141_);
  and (_25938_, _25874_, _24141_);
  nor (_25939_, _25938_, _25937_);
  nor (_25940_, _25939_, _25470_);
  nor (_25941_, _25424_, _24141_);
  not (_25942_, _25941_);
  and (_25943_, _25549_, _24278_);
  and (_25944_, _25426_, _24120_);
  nor (_25945_, _25944_, _25943_);
  and (_25946_, _25945_, _25942_);
  and (_25947_, _25413_, _25223_);
  nor (_25948_, _25411_, _25222_);
  not (_25949_, _25948_);
  and (_25950_, _25416_, _25221_);
  and (_25951_, _25418_, _24141_);
  nor (_25952_, _25951_, _25950_);
  nand (_25953_, _25952_, _25949_);
  nor (_25954_, _25953_, _25947_);
  and (_25955_, _25954_, _25946_);
  not (_25956_, _25955_);
  nor (_25957_, _25956_, _25940_);
  and (_25958_, _25957_, _25936_);
  not (_25959_, _25958_);
  nor (_25960_, _25959_, _25924_);
  and (_25961_, _25960_, _25920_);
  and (_25962_, _25961_, _25916_);
  and (_25963_, _25962_, _25914_);
  not (_25964_, _25963_);
  or (_25965_, _25964_, _25132_);
  not (_25966_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_25967_, _25132_, _25966_);
  and (_25968_, _25967_, _25450_);
  and (_25969_, _25968_, _25965_);
  nor (_25970_, _25449_, _25966_);
  nor (_25971_, _25020_, _25042_);
  and (_25972_, _25971_, _25053_);
  and (_25973_, _25972_, _25131_);
  nand (_25974_, _25973_, _25514_);
  or (_25975_, _25973_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_25976_, _25975_, _25521_);
  and (_25977_, _25976_, _25974_);
  or (_25978_, _25977_, _25970_);
  or (_25979_, _25978_, _25969_);
  and (_08909_, _25979_, _27355_);
  and (_25980_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_25981_, _25980_);
  nor (_25982_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_25983_, _25982_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_25984_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_25985_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_25986_, _25985_, _25984_);
  and (_25987_, _25982_, _23914_);
  and (_25988_, _25987_, _25986_);
  and (_25989_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_25990_, _25989_);
  not (_25991_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_25992_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_25993_, _25992_);
  not (_25994_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand (_25995_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_25996_, _25995_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or (_25997_, _25996_, _25994_);
  not (_25998_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not (_25999_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_26000_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_26001_, _26000_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_26002_, _26001_, _25999_);
  or (_26003_, _26002_, _25998_);
  and (_26004_, _26003_, _25997_);
  or (_26005_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_26006_, _26005_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_26007_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  not (_26008_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_26009_, _26005_, _25999_);
  or (_26010_, _26009_, _26008_);
  and (_26011_, _26010_, _26007_);
  nor (_26012_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_26013_, _26012_, _25999_);
  nand (_26014_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_26015_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not (_26016_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_26017_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26016_);
  nand (_26018_, _26017_, _25999_);
  or (_26019_, _26018_, _26015_);
  and (_26020_, _26019_, _26014_);
  and (_26021_, _26020_, _26011_);
  nand (_26022_, _26021_, _26004_);
  nand (_26023_, _26022_, _25993_);
  nand (_26024_, _26023_, _25991_);
  nor (_26025_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _25991_);
  nor (_26026_, _26025_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_26027_, _26026_, _26024_);
  and (_26028_, _26027_, _25990_);
  nand (_26029_, _26028_, _25988_);
  not (_26030_, _25986_);
  nor (_26031_, _25987_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_26032_, _26031_, _26030_);
  and (_26033_, _26032_, _26029_);
  not (_26034_, _26033_);
  not (_26035_, _25988_);
  and (_26036_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_26037_, _26036_);
  not (_26038_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_26039_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand (_26041_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  not (_26043_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_26045_, _26018_, _26043_);
  and (_26047_, _26045_, _26041_);
  nand (_26049_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not (_26051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_26053_, _26009_, _26051_);
  and (_26055_, _26053_, _26049_);
  not (_26057_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_26059_, _25996_, _26057_);
  not (_26061_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_26063_, _26002_, _26061_);
  and (_26065_, _26063_, _26059_);
  and (_26067_, _26065_, _26055_);
  nand (_26069_, _26067_, _26047_);
  nand (_26071_, _26069_, _25993_);
  nor (_26073_, _26071_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_26075_, _26073_, _26039_);
  nand (_26077_, _26075_, _26038_);
  nand (_26079_, _26077_, _26037_);
  or (_26081_, _26079_, _26035_);
  nor (_26083_, _25987_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_26085_, _26083_, _26030_);
  nand (_26087_, _26085_, _26081_);
  and (_26089_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_26091_, _26089_);
  not (_26093_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_26095_, _26002_, _26093_);
  not (_26097_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_26099_, _26018_, _26097_);
  and (_26101_, _26099_, _26095_);
  nand (_26103_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  not (_26105_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_26107_, _26009_, _26105_);
  and (_26109_, _26107_, _26103_);
  nand (_26110_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  not (_26111_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_26112_, _25996_, _26111_);
  and (_26113_, _26112_, _26110_);
  and (_26114_, _26113_, _26109_);
  and (_26115_, _26114_, _26101_);
  or (_26116_, _26115_, _25992_);
  nand (_26117_, _26116_, _25991_);
  nor (_26118_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _25991_);
  nor (_26119_, _26118_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_26120_, _26119_, _26117_);
  and (_26121_, _26120_, _26091_);
  nand (_26122_, _26121_, _25988_);
  nor (_26123_, _25987_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_26124_, _26123_, _26030_);
  and (_26125_, _26124_, _26122_);
  not (_26126_, _26125_);
  not (_26127_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_26128_, _26009_, _26127_);
  not (_26129_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_26130_, _25996_, _26129_);
  and (_26131_, _26130_, _26128_);
  not (_26132_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_26133_, _26018_, _26132_);
  and (_26134_, _26133_, _26131_);
  not (_26135_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_26136_, _26002_, _26135_);
  and (_26137_, _26136_, _25993_);
  nand (_26138_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_26139_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_26140_, _26139_, _26138_);
  and (_26141_, _26140_, _26137_);
  nand (_26142_, _26141_, _26134_);
  nor (_26143_, _26142_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_26144_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _25991_);
  or (_26145_, _26144_, _26143_);
  nand (_26146_, _26145_, _26038_);
  nor (_26147_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _26038_);
  not (_26148_, _26147_);
  and (_26149_, _26148_, _26146_);
  or (_26150_, _26149_, _26035_);
  nor (_26151_, _25987_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_26152_, _26151_, _26030_);
  and (_26153_, _26152_, _26150_);
  and (_26154_, _26153_, _26126_);
  and (_26155_, _26154_, _26087_);
  and (_26156_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not (_26157_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_26158_, _26009_, _26157_);
  not (_26159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_26160_, _25996_, _26159_);
  nand (_26161_, _26160_, _26158_);
  nor (_26162_, _26161_, _26156_);
  not (_26163_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_26164_, _26002_, _26163_);
  and (_26165_, _26164_, _25993_);
  nand (_26166_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not (_26167_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_26168_, _26018_, _26167_);
  and (_26169_, _26168_, _26166_);
  and (_26170_, _26169_, _26165_);
  nand (_26171_, _26170_, _26162_);
  or (_26172_, _26171_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_26173_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _25991_);
  nor (_26174_, _26173_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_26175_, _26174_, _26172_);
  and (_26176_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_26177_, _26176_, _26175_);
  or (_26178_, _26177_, _26035_);
  nor (_26179_, _25987_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_26180_, _26179_, _26030_);
  and (_26181_, _26180_, _26178_);
  and (_26182_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not (_26183_, _26182_);
  and (_26184_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nand (_26185_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not (_26186_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_26187_, _26018_, _26186_);
  and (_26188_, _26187_, _26185_);
  nand (_26189_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not (_26190_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or (_26191_, _26009_, _26190_);
  and (_26192_, _26191_, _26189_);
  not (_26193_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_26194_, _25996_, _26193_);
  not (_26195_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_26196_, _26002_, _26195_);
  and (_26197_, _26196_, _26194_);
  and (_26198_, _26197_, _26192_);
  nand (_26199_, _26198_, _26188_);
  nand (_26200_, _26199_, _25993_);
  nor (_26201_, _26200_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_26202_, _26201_, _26184_);
  nand (_26203_, _26202_, _26038_);
  nand (_26204_, _26203_, _26183_);
  or (_26205_, _26204_, _26035_);
  nor (_26206_, _25987_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_26207_, _26206_, _26030_);
  nand (_26208_, _26207_, _26205_);
  not (_26209_, _26208_);
  and (_26210_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_26211_, _26210_);
  not (_26212_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_26213_, _25996_, _26212_);
  not (_26214_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_26215_, _26002_, _26214_);
  and (_26216_, _26215_, _26213_);
  nand (_26217_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not (_26218_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or (_26219_, _26009_, _26218_);
  and (_26220_, _26219_, _26217_);
  nand (_26221_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_26222_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_26223_, _26018_, _26222_);
  and (_26224_, _26223_, _26221_);
  and (_26225_, _26224_, _26220_);
  nand (_26226_, _26225_, _26216_);
  and (_26227_, _26226_, _25993_);
  or (_26228_, _26227_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_26229_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _25991_);
  nor (_26230_, _26229_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_26231_, _26230_, _26228_);
  nand (_26232_, _26231_, _26211_);
  or (_26233_, _26232_, _26035_);
  nor (_26234_, _25987_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_26235_, _26234_, _26030_);
  and (_26236_, _26235_, _26233_);
  and (_26237_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_26238_, _26237_);
  and (_26239_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_26240_, _25992_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand (_26241_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  not (_26242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_26243_, _26002_, _26242_);
  and (_26244_, _26243_, _26241_);
  not (_26245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_26246_, _25996_, _26245_);
  not (_26247_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_26248_, _26018_, _26247_);
  and (_26249_, _26248_, _26246_);
  nand (_26250_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  not (_26251_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_26252_, _26009_, _26251_);
  and (_26253_, _26252_, _26250_);
  and (_26254_, _26253_, _26249_);
  and (_26255_, _26254_, _26244_);
  nor (_26256_, _26255_, _26240_);
  or (_26257_, _26256_, _26239_);
  nand (_26258_, _26257_, _26038_);
  nand (_26259_, _26258_, _26238_);
  or (_26260_, _26259_, _26035_);
  nor (_26261_, _25987_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_26262_, _26261_, _26030_);
  nand (_26263_, _26262_, _26260_);
  and (_26264_, _26263_, _26236_);
  and (_26265_, _26264_, _26209_);
  and (_26266_, _26265_, _26181_);
  and (_26267_, _26266_, _26155_);
  and (_26268_, _26267_, _26034_);
  not (_26269_, _26181_);
  nor (_26270_, _26263_, _26236_);
  and (_26271_, _26270_, _26209_);
  and (_26272_, _26271_, _26269_);
  and (_26273_, _26155_, _26034_);
  and (_26274_, _26273_, _26272_);
  or (_26275_, _26274_, _26268_);
  not (_26276_, _26275_);
  and (_26277_, _26125_, _26087_);
  not (_26278_, _26153_);
  and (_26279_, _26278_, _26033_);
  and (_26280_, _26279_, _26277_);
  and (_26281_, _26270_, _26208_);
  and (_26282_, _26281_, _26269_);
  and (_26283_, _26282_, _26280_);
  and (_26284_, _26126_, _26087_);
  nor (_26285_, _26153_, _26033_);
  and (_26286_, _26285_, _26284_);
  and (_26287_, _26286_, _26265_);
  or (_26288_, _26287_, _26283_);
  and (_26289_, _26271_, _26181_);
  and (_26290_, _26289_, _26280_);
  nand (_26291_, _26235_, _26233_);
  and (_26292_, _26263_, _26291_);
  and (_26293_, _26292_, _26208_);
  and (_26294_, _26293_, _26181_);
  and (_26295_, _26294_, _26280_);
  nor (_26296_, _26295_, _26290_);
  nor (_26297_, _26263_, _26291_);
  and (_26298_, _26297_, _26208_);
  and (_26299_, _26298_, _26181_);
  and (_26300_, _26299_, _26273_);
  and (_26301_, _26282_, _26155_);
  nor (_26302_, _26301_, _26300_);
  nand (_26303_, _26302_, _26296_);
  nor (_26304_, _26303_, _26288_);
  and (_26305_, _26304_, _26276_);
  and (_26306_, _26289_, _26155_);
  and (_26307_, _26306_, _26034_);
  and (_26308_, _26265_, _26269_);
  and (_26309_, _26308_, _26273_);
  nor (_26310_, _26309_, _26307_);
  and (_26311_, _26264_, _26208_);
  and (_26312_, _26311_, _26181_);
  and (_26313_, _26312_, _26286_);
  and (_26314_, _26311_, _26269_);
  and (_26315_, _26314_, _26286_);
  and (_26316_, _26294_, _26286_);
  or (_26317_, _26316_, _26315_);
  or (_26318_, _26317_, _26313_);
  not (_26319_, _26318_);
  and (_26320_, _26293_, _26269_);
  nand (_26321_, _26320_, _26280_);
  not (_26322_, _26087_);
  and (_26323_, _26308_, _26322_);
  not (_26324_, _26323_);
  and (_26325_, _26153_, _26125_);
  and (_26326_, _26325_, _26087_);
  and (_26327_, _26326_, _26269_);
  nand (_26328_, _26327_, _26265_);
  and (_26329_, _26328_, _26324_);
  and (_26330_, _26329_, _26321_);
  and (_26331_, _26330_, _26319_);
  and (_26332_, _26331_, _26310_);
  and (_26333_, _26281_, _26181_);
  and (_26334_, _26333_, _26155_);
  and (_26335_, _26292_, _26209_);
  and (_26336_, _26335_, _26269_);
  and (_26337_, _26336_, _26273_);
  nor (_26338_, _26337_, _26334_);
  or (_26339_, _26333_, _26311_);
  and (_26340_, _26339_, _26280_);
  and (_26341_, _26298_, _26269_);
  and (_26342_, _26341_, _26155_);
  and (_26343_, _26286_, _26271_);
  or (_26344_, _26343_, _26342_);
  nor (_26345_, _26344_, _26340_);
  and (_26346_, _26345_, _26338_);
  and (_26347_, _26341_, _26280_);
  and (_26348_, _26280_, _26272_);
  nor (_26349_, _26348_, _26347_);
  and (_26350_, _26297_, _26209_);
  and (_26351_, _26350_, _26269_);
  nand (_26352_, _26351_, _26280_);
  and (_26353_, _26311_, _26273_);
  not (_26354_, _26353_);
  and (_26355_, _26354_, _26352_);
  and (_26356_, _26355_, _26349_);
  and (_26357_, _26336_, _26280_);
  not (_26358_, _26357_);
  and (_26359_, _26335_, _26181_);
  nand (_26360_, _26359_, _26273_);
  and (_26361_, _26360_, _26358_);
  or (_26362_, _26359_, _26266_);
  nand (_26363_, _26362_, _26280_);
  and (_26364_, _26363_, _26361_);
  and (_26365_, _26364_, _26356_);
  and (_26366_, _26365_, _26346_);
  and (_26367_, _26366_, _26332_);
  nand (_26368_, _26367_, _26305_);
  nand (_26369_, _26368_, _25983_);
  not (_26370_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_26371_, _23914_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_26372_, _26371_, _26370_);
  not (_26373_, _26263_);
  and (_26374_, _26373_, _26208_);
  and (_26375_, _26286_, _26374_);
  and (_26376_, _26375_, _26372_);
  and (_26377_, _26153_, _26034_);
  and (_26378_, _26377_, _26284_);
  and (_26379_, _26378_, _26312_);
  and (_26380_, _26378_, _26314_);
  nor (_26381_, _26380_, _26379_);
  and (_26382_, \oc8051_top_1.oc8051_decoder1.state [0], _23914_);
  and (_26383_, _26382_, \oc8051_top_1.oc8051_decoder1.state [1]);
  not (_26384_, _26383_);
  nor (_26385_, _26384_, _26381_);
  nor (_26386_, _26385_, _26376_);
  nand (_26387_, _26386_, _26369_);
  nand (_26388_, _26387_, _23914_);
  and (_26389_, _26388_, _25981_);
  not (_26390_, _26389_);
  and (_26391_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26392_, _26391_);
  not (_26393_, _25983_);
  nand (_26394_, _26289_, _26286_);
  and (_26395_, _26354_, _26394_);
  and (_26396_, _26181_, _26087_);
  and (_26397_, _26396_, _26325_);
  and (_26398_, _26397_, _26265_);
  and (_26399_, _26326_, _26293_);
  nor (_26400_, _26399_, _26398_);
  and (_26401_, _26400_, _26395_);
  and (_26402_, _26397_, _26281_);
  and (_26403_, _26326_, _26311_);
  or (_26404_, _26403_, _26402_);
  and (_26405_, _26326_, _26271_);
  not (_26406_, _26405_);
  nand (_26407_, _26359_, _26326_);
  and (_26408_, _26407_, _26406_);
  not (_26409_, _26408_);
  nor (_26410_, _26409_, _26404_);
  and (_26411_, _26410_, _26401_);
  and (_26412_, _26154_, _26033_);
  and (_26413_, _26412_, _26087_);
  and (_26414_, _26308_, _26413_);
  not (_26415_, _26414_);
  nand (_26416_, _26359_, _26413_);
  nand (_26417_, _26299_, _26413_);
  and (_26418_, _26417_, _26416_);
  and (_26419_, _26418_, _26415_);
  and (_26420_, _26336_, _26326_);
  not (_26421_, _26420_);
  not (_26422_, _26327_);
  nor (_26423_, _26350_, _26281_);
  or (_26424_, _26423_, _26422_);
  nand (_26425_, _26341_, _26326_);
  and (_26426_, _26425_, _26424_);
  and (_26427_, _26426_, _26421_);
  and (_26428_, _26427_, _26419_);
  and (_26429_, _26428_, _26411_);
  or (_26430_, _26429_, _26393_);
  and (_26431_, _26298_, _26286_);
  and (_26432_, _26431_, _26372_);
  nor (_26433_, _26432_, _26385_);
  and (_26434_, _26433_, _26430_);
  or (_26435_, _26434_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_26436_, _26435_, _26392_);
  and (_26437_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_26438_, _26285_, _26277_);
  and (_26439_, _26438_, _26336_);
  and (_26440_, _26438_, _26308_);
  nor (_26441_, _26440_, _26439_);
  and (_26442_, _26441_, _26419_);
  nor (_26443_, _26442_, _26393_);
  not (_26444_, _26443_);
  and (_26445_, _26372_, _26286_);
  and (_26446_, _26445_, _26374_);
  and (_26447_, _26440_, _23914_);
  and (_26448_, _26439_, _23914_);
  nor (_26449_, _26448_, _26447_);
  nor (_26450_, _26449_, _25982_);
  nor (_26451_, _26450_, _26446_);
  and (_26452_, _26451_, _26444_);
  nor (_26453_, _26452_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_26454_, _26453_, _26437_);
  nand (_26455_, _26454_, _27355_);
  nor (_24440_, _26455_, _26436_);
  and (_09474_, _24440_, _26390_);
  and (_26456_, _25450_, _25115_);
  and (_26457_, _25128_, _25085_);
  not (_26458_, _25073_);
  nor (_26459_, _26458_, _25101_);
  and (_26460_, _26459_, _26457_);
  and (_26461_, _26460_, _25650_);
  and (_26462_, _26461_, _25020_);
  and (_26463_, _26462_, _26456_);
  not (_26464_, _26463_);
  and (_26465_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_26466_, _25239_, _24471_);
  nor (_26467_, _26466_, _24487_);
  and (_26468_, _26467_, _25915_);
  and (_26469_, _26468_, _25424_);
  nor (_26470_, _25426_, _25549_);
  and (_26471_, _26470_, _26469_);
  nor (_26472_, _26471_, _24141_);
  not (_26473_, _26472_);
  and (_26474_, _26473_, _25954_);
  and (_26475_, _26474_, _25936_);
  nor (_26476_, _26475_, _26464_);
  nor (_26477_, _26476_, _26465_);
  and (_26478_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_26479_, _26471_, _25364_);
  not (_26480_, _26479_);
  and (_26481_, _26480_, _25886_);
  and (_26482_, _26481_, _25871_);
  nor (_26483_, _26482_, _26464_);
  nor (_26484_, _26483_, _26478_);
  and (_26485_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_26486_, _26471_, _23973_);
  not (_26487_, _26486_);
  and (_26488_, _26487_, _25820_);
  and (_26489_, _26488_, _25808_);
  nor (_26490_, _26489_, _26464_);
  nor (_26491_, _26490_, _26485_);
  and (_26492_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_26493_, _26471_, _24101_);
  not (_26494_, _26493_);
  and (_26495_, _26494_, _25749_);
  and (_26496_, _26495_, _25746_);
  and (_26497_, _26496_, _25737_);
  nor (_26498_, _26497_, _26464_);
  nor (_26499_, _26498_, _26492_);
  and (_26500_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_26501_, _26471_, _25664_);
  not (_26502_, _26501_);
  and (_26503_, _26502_, _25681_);
  and (_26504_, _26503_, _25685_);
  and (_26505_, _26504_, _25672_);
  nor (_26506_, _26505_, _26464_);
  nor (_26507_, _26506_, _26500_);
  and (_26508_, _26464_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_26509_, _26471_, _25355_);
  not (_26510_, _26509_);
  and (_26511_, _26510_, _25608_);
  and (_26512_, _26511_, _25636_);
  nor (_26513_, _26512_, _26464_);
  nor (_26514_, _26513_, _26508_);
  and (_26515_, _26456_, _25020_);
  and (_26516_, _26515_, _26461_);
  nor (_26517_, _26516_, _25046_);
  nor (_26518_, _26471_, _24253_);
  not (_26519_, _26518_);
  and (_26520_, _26519_, _25546_);
  and (_26521_, _26520_, _25543_);
  not (_26522_, _26521_);
  and (_26523_, _26522_, _26516_);
  nor (_26524_, _26523_, _26517_);
  and (_26525_, _26524_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_26526_, _26525_, _26514_);
  and (_26527_, _26526_, _26507_);
  and (_26528_, _26527_, _26499_);
  and (_26529_, _26528_, _26491_);
  and (_26530_, _26529_, _26484_);
  and (_26531_, _26530_, _26477_);
  nor (_26532_, _26516_, _25087_);
  nand (_26533_, _26532_, _26531_);
  or (_26534_, _26532_, _26531_);
  and (_26535_, _26534_, _25061_);
  nand (_26536_, _26535_, _26533_);
  nor (_26537_, _26516_, _25091_);
  and (_26538_, _26537_, _26536_);
  nor (_26539_, _26471_, _24172_);
  not (_26540_, _26539_);
  and (_26541_, _26540_, _25420_);
  and (_26542_, _26541_, _25415_);
  and (_26543_, _26542_, _25385_);
  and (_26544_, _26543_, _26463_);
  nor (_26545_, _26544_, _26538_);
  and (_09496_, _26545_, _27355_);
  not (_26546_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_26547_, _26524_, _26546_);
  nor (_26548_, _26524_, _26546_);
  nor (_26549_, _26548_, _26547_);
  and (_26550_, _26549_, _25061_);
  nor (_26551_, _26550_, _25047_);
  nor (_26552_, _26551_, _26463_);
  nor (_26553_, _26552_, _26523_);
  nand (_10718_, _26553_, _27355_);
  nor (_26554_, _26525_, _26514_);
  nor (_26555_, _26554_, _26526_);
  nor (_26556_, _26555_, _24979_);
  nor (_26557_, _26556_, _25028_);
  nor (_26558_, _26557_, _26463_);
  nor (_26559_, _26558_, _26513_);
  nand (_10729_, _26559_, _27355_);
  nor (_26560_, _26526_, _26507_);
  nor (_26561_, _26560_, _26527_);
  nor (_26562_, _26561_, _24979_);
  nor (_26563_, _26562_, _24984_);
  nor (_26564_, _26563_, _26463_);
  nor (_26565_, _26564_, _26506_);
  nand (_10740_, _26565_, _27355_);
  nor (_26566_, _26527_, _26499_);
  nor (_26567_, _26566_, _26528_);
  nor (_26568_, _26567_, _24979_);
  nor (_26569_, _26568_, _25109_);
  nor (_26570_, _26569_, _26463_);
  nor (_26571_, _26570_, _26498_);
  nor (_10751_, _26571_, rst);
  nor (_26572_, _26528_, _26491_);
  nor (_26573_, _26572_, _26529_);
  nor (_26574_, _26573_, _24979_);
  nor (_26575_, _26574_, _25121_);
  nor (_26576_, _26575_, _26463_);
  nor (_26577_, _26576_, _26490_);
  nor (_10762_, _26577_, rst);
  nor (_26578_, _26529_, _26484_);
  nor (_26579_, _26578_, _26530_);
  nor (_26580_, _26579_, _24979_);
  nor (_26581_, _26580_, _25077_);
  nor (_26582_, _26581_, _26463_);
  nor (_26583_, _26582_, _26483_);
  nor (_10773_, _26583_, rst);
  nor (_26584_, _26530_, _26477_);
  nor (_26585_, _26584_, _26531_);
  nor (_26586_, _26585_, _24979_);
  nor (_26587_, _26586_, _25064_);
  nor (_26588_, _26587_, _26463_);
  nor (_26589_, _26588_, _26476_);
  nor (_10784_, _26589_, rst);
  and (_26590_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _23914_);
  and (_26591_, _26590_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_26592_, _26460_, _25778_);
  nand (_26593_, _26592_, _26456_);
  and (_26594_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_26595_, _25020_, _25115_);
  and (_26596_, _25516_, _26595_);
  and (_26597_, _26596_, _26460_);
  and (_26598_, _26597_, _25449_);
  and (_26599_, _26598_, _25444_);
  and (_26600_, _26599_, _25441_);
  or (_26601_, _26600_, _26594_);
  or (_26602_, _26601_, _26591_);
  not (_26603_, _26591_);
  nor (_26604_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_26605_, _24108_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26606_, _26605_, _26604_);
  nor (_26607_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_26608_, _24089_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26609_, _26608_, _26607_);
  nor (_26610_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_26611_, _24240_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26612_, _26611_, _26610_);
  not (_26613_, _26612_);
  nor (_26614_, _26613_, _25461_);
  nor (_26615_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_26616_, _24188_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26617_, _26616_, _26615_);
  and (_26618_, _26617_, _26614_);
  nor (_26619_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_26620_, _24204_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26621_, _26620_, _26619_);
  and (_26622_, _26621_, _26618_);
  and (_26623_, _26622_, _26609_);
  nor (_26624_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_26625_, _23940_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26626_, _26625_, _26624_);
  and (_26627_, _26626_, _26623_);
  and (_26628_, _26627_, _26606_);
  nor (_26629_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_26630_, _24129_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26631_, _26630_, _26629_);
  and (_26632_, _26631_, _26628_);
  nor (_26633_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_26634_, _24158_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_26635_, _26634_, _26633_);
  or (_26636_, _26635_, _26632_);
  nand (_26637_, _26635_, _26632_);
  and (_26638_, _26637_, _26636_);
  and (_26639_, _26638_, _25240_);
  and (_26640_, _24443_, _23920_);
  and (_26641_, _25361_, _24278_);
  and (_26642_, _26641_, _24082_);
  and (_26643_, _26642_, _24032_);
  and (_26644_, _26643_, _24515_);
  and (_26645_, _26644_, _24533_);
  and (_26646_, _26645_, _24520_);
  or (_26647_, _26646_, _25363_);
  and (_26648_, _25370_, _24172_);
  and (_26649_, _24018_, _24068_);
  nor (_26650_, _24032_, _24082_);
  and (_26651_, _26650_, _26649_);
  and (_26652_, _26651_, _26648_);
  and (_26653_, _24004_, _24055_);
  and (_26654_, _26653_, _26652_);
  nor (_26655_, _26654_, _25199_);
  not (_26656_, _26655_);
  nand (_26657_, _25199_, _24004_);
  and (_26658_, _26657_, _26656_);
  and (_26659_, _26658_, _26647_);
  and (_26660_, _25199_, _24616_);
  nor (_26661_, _26660_, _25926_);
  and (_26662_, _26661_, _26659_);
  or (_26663_, _26662_, _25377_);
  nand (_26664_, _26662_, _25377_);
  and (_26665_, _26664_, _26663_);
  and (_26666_, _26665_, _25354_);
  and (_26667_, _25199_, _25377_);
  or (_26668_, _26667_, _25472_);
  and (_26669_, _26668_, _25381_);
  nor (_26670_, _25502_, _24101_);
  nor (_26671_, _25424_, _23990_);
  and (_26672_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or (_26673_, _26672_, _26671_);
  or (_26674_, _26673_, _26670_);
  or (_26675_, _26674_, _26669_);
  or (_26676_, _26675_, _26666_);
  or (_26677_, _26676_, _26640_);
  or (_26678_, _26677_, _26639_);
  or (_26679_, _26678_, _26603_);
  and (_26680_, _26679_, _27355_);
  and (_12743_, _26680_, _26602_);
  and (_26681_, _26456_, _25716_);
  and (_26682_, _26681_, _26460_);
  nor (_26683_, _26682_, _26591_);
  or (_26684_, _26683_, _25441_);
  not (_26685_, _26683_);
  or (_26686_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_26687_, _26686_, _27355_);
  and (_12764_, _26687_, _26684_);
  nor (_26688_, _26593_, _25562_);
  and (_26689_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_26690_, _26689_, _26591_);
  or (_26691_, _26690_, _26688_);
  and (_26692_, _26613_, _25461_);
  nor (_26693_, _26692_, _26614_);
  and (_26694_, _26693_, _25240_);
  nand (_26695_, _24923_, _24487_);
  nor (_26696_, _25472_, _25380_);
  not (_26697_, _26696_);
  nor (_26698_, _26697_, _25372_);
  nor (_26699_, _26698_, _24082_);
  and (_26700_, _26698_, _24082_);
  nor (_26701_, _26700_, _26699_);
  and (_26702_, _26701_, _25354_);
  and (_26703_, _25423_, _24082_);
  and (_26704_, _24394_, _23920_);
  nor (_26705_, _25502_, _23973_);
  nor (_26706_, _25382_, _24253_);
  or (_26707_, _26706_, _26705_);
  or (_26708_, _26707_, _26704_);
  nor (_26709_, _26708_, _26703_);
  not (_26710_, _26709_);
  nor (_26711_, _26710_, _26702_);
  nand (_26712_, _26711_, _26695_);
  or (_26713_, _26712_, _26694_);
  or (_26714_, _26713_, _26603_);
  and (_26715_, _26714_, _27355_);
  and (_13683_, _26715_, _26691_);
  and (_26716_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_26717_, _26599_, _25639_);
  or (_26718_, _26717_, _26716_);
  or (_26719_, _26718_, _26591_);
  nor (_26720_, _26617_, _26614_);
  not (_26721_, _26720_);
  nor (_26722_, _26618_, _25459_);
  and (_26723_, _26722_, _26721_);
  not (_26724_, _26723_);
  and (_26725_, _24632_, _24487_);
  not (_26726_, _26725_);
  and (_26727_, _25423_, _24032_);
  nor (_26728_, _26642_, _25363_);
  and (_26729_, _26648_, _25146_);
  nor (_26730_, _26729_, _25199_);
  or (_26731_, _26730_, _26728_);
  and (_26732_, _26731_, _25310_);
  not (_26733_, _26732_);
  nor (_26734_, _26731_, _25310_);
  nor (_26735_, _26734_, _25867_);
  and (_26736_, _26735_, _26733_);
  and (_26737_, _24396_, _23920_);
  and (_26738_, _25501_, _24120_);
  and (_26739_, _25381_, _24200_);
  or (_26740_, _26739_, _26738_);
  or (_26741_, _26740_, _26737_);
  or (_26742_, _26741_, _26736_);
  nor (_26743_, _26742_, _26727_);
  and (_26744_, _26743_, _26726_);
  and (_26745_, _26744_, _26724_);
  nand (_26746_, _26745_, _26591_);
  and (_26747_, _26746_, _27355_);
  and (_13694_, _26747_, _26719_);
  nor (_26748_, _26593_, _25704_);
  and (_26749_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_26750_, _26749_, _26591_);
  or (_26751_, _26750_, _26748_);
  nor (_26752_, _26621_, _26618_);
  nor (_26753_, _26752_, _26622_);
  and (_26754_, _26753_, _25240_);
  not (_26755_, _26754_);
  and (_26756_, _26729_, _25310_);
  and (_26757_, _26756_, _25363_);
  and (_26758_, _26643_, _25199_);
  nor (_26759_, _26758_, _26757_);
  and (_26760_, _26759_, _24068_);
  nor (_26761_, _26759_, _24068_);
  nor (_26762_, _26761_, _26760_);
  and (_26763_, _26762_, _25354_);
  and (_26764_, _25381_, _24216_);
  and (_26765_, _25423_, _24515_);
  nor (_26766_, _26765_, _26764_);
  and (_26767_, _24398_, _23920_);
  nor (_26768_, _25502_, _24141_);
  and (_26769_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_26770_, _26769_, _26768_);
  nor (_26771_, _26770_, _26767_);
  and (_26772_, _26771_, _26766_);
  not (_26773_, _26772_);
  nor (_26774_, _26773_, _26763_);
  and (_26775_, _26774_, _26755_);
  nand (_26776_, _26775_, _26591_);
  and (_26777_, _26776_, _27355_);
  and (_13705_, _26777_, _26751_);
  nor (_26778_, _26593_, _25769_);
  and (_26779_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_26780_, _26779_, _26591_);
  or (_26781_, _26780_, _26778_);
  nor (_26782_, _26622_, _26609_);
  not (_26783_, _26782_);
  nor (_26784_, _26623_, _25459_);
  and (_26785_, _26784_, _26783_);
  not (_26786_, _26785_);
  and (_26787_, _24401_, _23920_);
  not (_26788_, _26787_);
  nor (_26789_, _26645_, _25363_);
  nor (_26790_, _26644_, _24533_);
  not (_26791_, _26790_);
  and (_26792_, _26791_, _26789_);
  and (_26793_, _26756_, _24068_);
  nor (_26794_, _26793_, _24018_);
  nor (_26795_, _26794_, _26652_);
  nor (_26796_, _26795_, _25199_);
  nor (_26797_, _26796_, _26792_);
  nor (_26798_, _26797_, _25867_);
  and (_26799_, _25423_, _24533_);
  nor (_26800_, _25382_, _24101_);
  and (_26801_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_26802_, _26801_, _26800_);
  or (_26803_, _26802_, _25503_);
  nor (_26804_, _26803_, _26799_);
  not (_26805_, _26804_);
  nor (_26806_, _26805_, _26798_);
  and (_26807_, _26806_, _26788_);
  and (_26808_, _26807_, _26786_);
  nand (_26809_, _26808_, _26591_);
  and (_26810_, _26809_, _27355_);
  and (_13716_, _26810_, _26781_);
  and (_26811_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_26812_, _26599_, _25830_);
  or (_26813_, _26812_, _26811_);
  or (_26814_, _26813_, _26591_);
  or (_26815_, _26626_, _26623_);
  nor (_26816_, _26627_, _25459_);
  and (_26817_, _26816_, _26815_);
  nor (_26818_, _26652_, _25199_);
  nor (_26819_, _26818_, _26789_);
  or (_26820_, _26819_, _24520_);
  nand (_26821_, _26819_, _24520_);
  and (_26822_, _26821_, _26820_);
  and (_26823_, _26822_, _25354_);
  and (_26824_, _24403_, _23920_);
  or (_26825_, _25199_, _23974_);
  nand (_26826_, _25199_, _24055_);
  and (_26827_, _26826_, _25381_);
  and (_26828_, _26827_, _26825_);
  nor (_26829_, _25502_, _24253_);
  and (_26830_, _25423_, _24520_);
  and (_26831_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_26832_, _26831_, _26830_);
  or (_26833_, _26832_, _26829_);
  or (_26834_, _26833_, _26828_);
  or (_26835_, _26834_, _26824_);
  or (_26836_, _26835_, _26823_);
  or (_26837_, _26836_, _26817_);
  or (_26838_, _26837_, _26603_);
  and (_26839_, _26838_, _27355_);
  and (_13727_, _26839_, _26814_);
  and (_26840_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_26841_, _26599_, _25898_);
  or (_26842_, _26841_, _26840_);
  or (_26843_, _26842_, _26591_);
  or (_26844_, _26627_, _26606_);
  nor (_26845_, _26628_, _25459_);
  and (_26846_, _26845_, _26844_);
  and (_26847_, _24413_, _23920_);
  and (_26848_, _26652_, _24055_);
  nor (_26849_, _26848_, _25199_);
  not (_26850_, _26849_);
  and (_26851_, _26850_, _26647_);
  and (_26852_, _26851_, _24004_);
  nor (_26853_, _26851_, _24004_);
  or (_26854_, _26853_, _26852_);
  and (_26855_, _26854_, _25354_);
  or (_26856_, _25199_, _24120_);
  and (_26857_, _26657_, _25381_);
  and (_26858_, _26857_, _26856_);
  and (_26859_, _25501_, _24200_);
  and (_26860_, _25423_, _24535_);
  and (_26861_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_26862_, _26861_, _26860_);
  or (_26863_, _26862_, _26859_);
  or (_26864_, _26863_, _26858_);
  or (_26865_, _26864_, _26855_);
  or (_26866_, _26865_, _26847_);
  or (_26867_, _26866_, _26846_);
  or (_26868_, _26867_, _26603_);
  and (_26869_, _26868_, _27355_);
  and (_13738_, _26869_, _26843_);
  nor (_26870_, _26593_, _25963_);
  and (_26871_, _26593_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_26872_, _26871_, _26591_);
  or (_26873_, _26872_, _26870_);
  nor (_26874_, _26631_, _26628_);
  nor (_26875_, _26874_, _26632_);
  and (_26876_, _26875_, _25240_);
  not (_26877_, _26876_);
  and (_26878_, _24441_, _23920_);
  nor (_26879_, _26659_, _24616_);
  and (_26880_, _26659_, _24616_);
  nor (_26881_, _26880_, _26879_);
  nor (_26882_, _26881_, _25867_);
  nor (_26883_, _25199_, _24143_);
  not (_26884_, _26883_);
  nor (_26885_, _26660_, _25382_);
  and (_26886_, _26885_, _26884_);
  and (_26887_, _24487_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  and (_26888_, _25501_, _24216_);
  and (_26889_, _25423_, _24049_);
  or (_26890_, _26889_, _26888_);
  nor (_26891_, _26890_, _26887_);
  not (_26892_, _26891_);
  nor (_26893_, _26892_, _26886_);
  not (_26894_, _26893_);
  nor (_26895_, _26894_, _26882_);
  not (_26896_, _26895_);
  nor (_26897_, _26896_, _26878_);
  and (_26898_, _26897_, _26877_);
  nand (_26899_, _26898_, _26591_);
  and (_26900_, _26899_, _27355_);
  and (_13749_, _26900_, _26873_);
  nand (_26901_, _26685_, _25562_);
  or (_26902_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_26903_, _26902_, _27355_);
  and (_13760_, _26903_, _26901_);
  or (_26904_, _26683_, _25639_);
  or (_26905_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_26906_, _26905_, _27355_);
  and (_13771_, _26906_, _26904_);
  nand (_26907_, _26685_, _25704_);
  or (_26908_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_26909_, _26908_, _27355_);
  and (_13782_, _26909_, _26907_);
  nand (_26910_, _26685_, _25769_);
  or (_26911_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_26912_, _26911_, _27355_);
  and (_13793_, _26912_, _26910_);
  or (_26913_, _26683_, _25830_);
  or (_26914_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_26915_, _26914_, _27355_);
  and (_13804_, _26915_, _26913_);
  or (_26916_, _26683_, _25898_);
  or (_26917_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_26918_, _26917_, _27355_);
  and (_13815_, _26918_, _26916_);
  nand (_26919_, _26685_, _25963_);
  or (_26920_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_26921_, _26920_, _27355_);
  and (_13826_, _26921_, _26919_);
  not (_26922_, _25085_);
  nor (_26923_, _26922_, _25073_);
  and (_26924_, _26923_, _25521_);
  and (_26925_, _26924_, _25130_);
  not (_26926_, _25517_);
  nor (_26927_, _26926_, _25514_);
  not (_26928_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_26929_, _25517_, _26928_);
  or (_26930_, _26929_, _26927_);
  and (_26931_, _26930_, _26925_);
  nor (_26932_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_26933_, _26932_);
  nand (_26934_, _26933_, _25514_);
  and (_26935_, _26932_, _26928_);
  nor (_26936_, _26935_, _26925_);
  and (_26937_, _26936_, _26934_);
  nor (_26938_, _25128_, _26922_);
  nor (_26939_, _25073_, _25101_);
  and (_26940_, _26456_, _25055_);
  and (_26941_, _26940_, _26939_);
  and (_26942_, _26941_, _26938_);
  or (_26943_, _26942_, _26937_);
  or (_26944_, _26943_, _26931_);
  nand (_26945_, _26942_, _26543_);
  and (_26946_, _26945_, _27355_);
  and (_15222_, _26946_, _26944_);
  and (_26947_, _25650_, _25020_);
  and (_26948_, _26925_, _26947_);
  nand (_26949_, _26948_, _25514_);
  not (_26950_, _26942_);
  or (_26951_, _26948_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_26952_, _26951_, _26950_);
  and (_26953_, _26952_, _26949_);
  nor (_26954_, _26950_, _26512_);
  or (_26955_, _26954_, _26953_);
  and (_17288_, _26955_, _27355_);
  or (_26956_, _24452_, _24448_);
  or (_26957_, _26956_, _24456_);
  or (_26958_, _26957_, _24460_);
  nor (_26959_, _26958_, _24465_);
  nand (_26960_, _26959_, _24467_);
  and (_26961_, _26960_, _23920_);
  and (_26962_, _25465_, _25348_);
  not (_26963_, _25348_);
  and (_26964_, _25466_, _26963_);
  or (_26965_, _26964_, _26962_);
  and (_26966_, _26965_, _25246_);
  not (_26967_, _25233_);
  nand (_26968_, _25232_, _26967_);
  or (_26969_, _25234_, _25232_);
  and (_26970_, _25240_, _26969_);
  and (_26971_, _26970_, _26968_);
  and (_26972_, _26653_, _24617_);
  and (_26973_, _26651_, _24487_);
  nand (_26974_, _26973_, _26972_);
  nand (_26975_, _26974_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_26976_, _26975_, _26971_);
  or (_26977_, _26976_, _26966_);
  or (_26978_, _26977_, _25789_);
  or (_26979_, _26978_, _25134_);
  or (_26980_, _26979_, _26961_);
  nor (_26981_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_26982_, _26981_, _26925_);
  and (_26983_, _26982_, _26980_);
  and (_26984_, _25717_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_26985_, _26984_, _25718_);
  and (_26986_, _26985_, _26925_);
  or (_26987_, _26986_, _26942_);
  or (_26988_, _26987_, _26983_);
  nand (_26989_, _26942_, _26505_);
  and (_26990_, _26989_, _27355_);
  and (_17297_, _26990_, _26988_);
  and (_26991_, _26925_, _25778_);
  nand (_26992_, _26991_, _25514_);
  or (_26993_, _26991_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_26994_, _26993_, _26950_);
  and (_26995_, _26994_, _26992_);
  nor (_26996_, _26950_, _26497_);
  or (_26997_, _26996_, _26995_);
  and (_17306_, _26997_, _27355_);
  not (_26998_, _26925_);
  or (_26999_, _26998_, _25840_);
  and (_27000_, _26999_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_27001_, _25839_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_27002_, _27001_, _25843_);
  and (_27003_, _27002_, _26925_);
  or (_27004_, _27003_, _27000_);
  and (_27005_, _27004_, _26950_);
  nor (_27006_, _26950_, _26489_);
  or (_27007_, _27006_, _27005_);
  and (_17315_, _27007_, _27355_);
  and (_27008_, _26925_, _25905_);
  nand (_27009_, _27008_, _25514_);
  or (_27010_, _27008_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_27011_, _27010_, _26950_);
  and (_27012_, _27011_, _27009_);
  nor (_27013_, _26950_, _26482_);
  or (_27014_, _27013_, _27012_);
  and (_17324_, _27014_, _27355_);
  and (_27015_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_27016_, _25240_, _25212_);
  and (_27017_, _25344_, _25246_);
  or (_27018_, _27017_, _27016_);
  and (_27019_, _27018_, _27015_);
  nand (_27020_, _27015_, _25424_);
  and (_27021_, _27020_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_27022_, _27021_, _26925_);
  or (_27023_, _27022_, _27019_);
  not (_27024_, _25972_);
  nor (_27025_, _27024_, _25514_);
  or (_27026_, _25972_, _25738_);
  nand (_27027_, _27026_, _26925_);
  or (_27028_, _27027_, _27025_);
  and (_27029_, _27028_, _27023_);
  or (_27030_, _27029_, _26942_);
  nand (_27031_, _26942_, _26475_);
  and (_27032_, _27031_, _27355_);
  and (_17332_, _27032_, _27030_);
  nor (_27033_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_27034_, _27033_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_27035_, _25055_, _25115_);
  and (_27036_, _25128_, _26922_);
  and (_27037_, _27036_, _26939_);
  and (_27038_, _27037_, _27035_);
  and (_27039_, _27038_, _25450_);
  nor (_27040_, _27039_, _27034_);
  not (_27041_, _27040_);
  and (_27042_, _27041_, _25441_);
  not (_27043_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_27044_, _26590_, _27043_);
  and (_27045_, _25128_, _25115_);
  and (_27046_, _27045_, _25086_);
  not (_27047_, _25521_);
  nor (_27048_, _27047_, _25101_);
  and (_27049_, _27048_, _27046_);
  and (_27050_, _27049_, _25517_);
  or (_27051_, _27050_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_27052_, _27044_);
  and (_27053_, _27052_, _27040_);
  nand (_27054_, _27050_, _25514_);
  and (_27055_, _27054_, _27053_);
  and (_27056_, _27055_, _27051_);
  or (_27057_, _27056_, _27044_);
  or (_27058_, _27057_, _27042_);
  or (_27059_, _27052_, _26678_);
  and (_27060_, _27059_, _27058_);
  and (_17824_, _27060_, _27355_);
  or (_27061_, _27040_, _25562_);
  and (_27062_, _27049_, _25055_);
  nor (_27063_, _27062_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not (_27064_, _27063_);
  not (_27065_, _27053_);
  and (_27066_, _27062_, _25514_);
  nor (_27067_, _27066_, _27065_);
  and (_27068_, _27067_, _27064_);
  nor (_27069_, _27068_, _27044_);
  nand (_27070_, _27069_, _27061_);
  or (_27071_, _27052_, _26713_);
  and (_27072_, _27071_, _27070_);
  and (_19498_, _27072_, _27355_);
  nor (_27073_, _27052_, _26745_);
  not (_27074_, _27073_);
  or (_27075_, _27040_, _25639_);
  nor (_27076_, _27049_, _24029_);
  not (_27077_, _27076_);
  not (_27078_, _27049_);
  not (_27079_, _26947_);
  nor (_27080_, _27079_, _25514_);
  nor (_27081_, _26947_, _24029_);
  nor (_27082_, _27081_, _27080_);
  or (_27083_, _27082_, _27078_);
  and (_27084_, _27083_, _27040_);
  and (_27085_, _27084_, _27077_);
  nor (_27086_, _27085_, _27044_);
  nand (_27087_, _27086_, _27075_);
  nand (_27088_, _27087_, _27074_);
  and (_19508_, _27088_, _27355_);
  or (_27089_, _27040_, _25704_);
  and (_27090_, _27049_, _25716_);
  and (_27091_, _27090_, _25514_);
  nor (_27092_, _27090_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_27093_, _27092_, _27065_);
  not (_27094_, _27093_);
  nor (_27095_, _27094_, _27091_);
  nor (_27096_, _27095_, _27044_);
  nand (_27097_, _27096_, _27089_);
  and (_27098_, _27044_, _26775_);
  not (_27099_, _27098_);
  and (_27100_, _27099_, _27097_);
  and (_19518_, _27100_, _27355_);
  or (_27101_, _27040_, _25769_);
  and (_27102_, _27053_, _27078_);
  and (_27103_, _27102_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_27104_, _25778_, _24015_);
  nor (_27105_, _27104_, _25779_);
  and (_27106_, _27049_, _27052_);
  not (_27107_, _27106_);
  nor (_27108_, _27107_, _27105_);
  and (_27109_, _27108_, _27053_);
  nor (_27110_, _27109_, _27103_);
  and (_27111_, _27110_, _27052_);
  nand (_27112_, _27111_, _27101_);
  and (_27113_, _27044_, _26808_);
  not (_27114_, _27113_);
  and (_27115_, _27114_, _27112_);
  and (_19528_, _27115_, _27355_);
  and (_27116_, _27041_, _25830_);
  and (_27117_, _27049_, _25838_);
  or (_27118_, _27117_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_27119_, _27117_, _25514_);
  and (_27120_, _27119_, _27053_);
  and (_27121_, _27120_, _27118_);
  or (_27122_, _27121_, _27044_);
  or (_27123_, _27122_, _27116_);
  or (_27124_, _27052_, _26837_);
  and (_27125_, _27124_, _27123_);
  and (_19539_, _27125_, _27355_);
  and (_27126_, _27041_, _25898_);
  and (_27127_, _27049_, _25905_);
  or (_27128_, _27127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_27129_, _27127_, _25514_);
  and (_27130_, _27129_, _27053_);
  and (_27131_, _27130_, _27128_);
  or (_27132_, _27131_, _27044_);
  or (_27133_, _27132_, _27126_);
  or (_27134_, _27052_, _26867_);
  and (_27135_, _27134_, _27133_);
  and (_19549_, _27135_, _27355_);
  or (_27136_, _27040_, _25963_);
  and (_27137_, _27049_, _25972_);
  nor (_27138_, _27137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_27139_, _27138_);
  and (_27140_, _27137_, _25514_);
  nor (_27141_, _27140_, _27065_);
  and (_27142_, _27141_, _27139_);
  nor (_27143_, _27142_, _27044_);
  and (_27144_, _27143_, _27136_);
  and (_27145_, _27044_, _26898_);
  or (_27146_, _27145_, _27144_);
  nor (_19559_, _27146_, rst);
  and (_27147_, _25085_, _25073_);
  and (_27148_, _27045_, _25102_);
  and (_27149_, _27148_, _27147_);
  and (_27150_, _27149_, _25517_);
  nand (_27151_, _27150_, _25514_);
  or (_27152_, _27150_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_27153_, _27152_, _25521_);
  and (_27154_, _27153_, _27151_);
  and (_27155_, _26460_, _27035_);
  nand (_27156_, _27155_, _26543_);
  or (_27157_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_27158_, _27157_, _25450_);
  and (_27159_, _27158_, _27156_);
  not (_27160_, _25449_);
  and (_27161_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_27162_, _27161_, rst);
  or (_27163_, _27162_, _27159_);
  or (_23900_, _27163_, _27154_);
  and (_27164_, _27147_, _25130_);
  and (_27165_, _27164_, _25517_);
  nand (_27166_, _27165_, _25514_);
  or (_27167_, _27165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_27168_, _27167_, _25521_);
  and (_27169_, _27168_, _27166_);
  and (_27170_, _26938_, _26459_);
  and (_27171_, _27170_, _27035_);
  nand (_27172_, _27171_, _26543_);
  or (_27173_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_27174_, _27173_, _25450_);
  and (_27175_, _27174_, _27172_);
  and (_27176_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_27177_, _27176_, rst);
  or (_27178_, _27177_, _27175_);
  or (_23901_, _27178_, _27169_);
  and (_27179_, _26922_, _25073_);
  and (_27180_, _27179_, _27148_);
  and (_27181_, _27180_, _25517_);
  nand (_27182_, _27181_, _25514_);
  or (_27183_, _27181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_27184_, _27183_, _25521_);
  and (_27185_, _27184_, _27182_);
  and (_27186_, _27036_, _26459_);
  and (_27187_, _27186_, _27035_);
  not (_27188_, _27187_);
  nor (_27189_, _27188_, _26543_);
  and (_27190_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_27191_, _27190_, _27189_);
  and (_27192_, _27191_, _25450_);
  and (_27193_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_27194_, _27193_, rst);
  or (_27195_, _27194_, _27192_);
  or (_23902_, _27195_, _27185_);
  and (_27196_, _27179_, _25130_);
  and (_27197_, _27196_, _25517_);
  nand (_27198_, _27197_, _25514_);
  or (_27199_, _27197_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_27200_, _27199_, _25521_);
  and (_27201_, _27200_, _27198_);
  nor (_27202_, _25128_, _25085_);
  and (_27203_, _26459_, _27202_);
  and (_27204_, _27203_, _27035_);
  not (_27205_, _27204_);
  nor (_27206_, _27205_, _26543_);
  and (_27207_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_27208_, _27207_, _27206_);
  and (_27209_, _27208_, _25450_);
  and (_27210_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_27211_, _27210_, rst);
  or (_27212_, _27211_, _27209_);
  or (_23903_, _27212_, _27201_);
  or (_27213_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_27214_, _27213_, _25521_);
  nand (_27215_, _27155_, _25514_);
  and (_27216_, _27215_, _27214_);
  nand (_27217_, _27155_, _26521_);
  and (_27218_, _27217_, _25450_);
  and (_27219_, _27218_, _27213_);
  not (_27220_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_27221_, _25449_, _27220_);
  or (_27222_, _27221_, rst);
  or (_27223_, _27222_, _27219_);
  or (_24987_, _27223_, _27216_);
  and (_27224_, _25650_, _26595_);
  and (_27225_, _27224_, _26460_);
  nand (_27226_, _27225_, _25514_);
  or (_27227_, _27225_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_27228_, _27227_, _25521_);
  and (_27229_, _27228_, _27226_);
  nand (_27230_, _27155_, _26512_);
  or (_27231_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_27232_, _27231_, _25450_);
  and (_27233_, _27232_, _27230_);
  and (_27234_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_27235_, _27234_, rst);
  or (_27236_, _27235_, _27233_);
  or (_24989_, _27236_, _27229_);
  not (_27237_, _25780_);
  nand (_27238_, _27149_, _27237_);
  and (_27239_, _27238_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not (_27240_, _25719_);
  and (_27241_, _27240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_27242_, _27241_, _25718_);
  and (_27243_, _27242_, _27149_);
  or (_27244_, _27243_, _27239_);
  and (_27245_, _27244_, _25521_);
  nand (_27246_, _27155_, _26505_);
  or (_27247_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_27248_, _27247_, _25450_);
  and (_27249_, _27248_, _27246_);
  and (_27250_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_27251_, _27250_, rst);
  or (_27252_, _27251_, _27249_);
  or (_24991_, _27252_, _27245_);
  nand (_27253_, _27149_, _25020_);
  and (_27254_, _27253_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_27255_, _27237_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_27256_, _27255_, _25779_);
  and (_27257_, _27256_, _27149_);
  or (_27258_, _27257_, _27254_);
  and (_27259_, _27258_, _25521_);
  nand (_27260_, _27155_, _26497_);
  or (_27261_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_27262_, _27261_, _25450_);
  and (_27263_, _27262_, _27260_);
  and (_27264_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_27265_, _27264_, rst);
  or (_27266_, _27265_, _27263_);
  or (_24993_, _27266_, _27259_);
  not (_27267_, _27149_);
  or (_27268_, _27267_, _25840_);
  and (_27269_, _27268_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_27270_, _25839_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_27271_, _27270_, _25843_);
  and (_27272_, _27271_, _27149_);
  or (_27273_, _27272_, _27269_);
  and (_27274_, _27273_, _25521_);
  nand (_27275_, _27155_, _26489_);
  or (_27276_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_27277_, _27276_, _25450_);
  and (_27278_, _27277_, _27275_);
  and (_27279_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_27280_, _27279_, rst);
  or (_27281_, _27280_, _27278_);
  or (_24995_, _27281_, _27274_);
  and (_27282_, _27149_, _25905_);
  nand (_27283_, _27282_, _25514_);
  or (_27284_, _27282_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_27285_, _27284_, _25521_);
  and (_27286_, _27285_, _27283_);
  nand (_27287_, _27155_, _26482_);
  or (_27288_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_27289_, _27288_, _25450_);
  and (_27290_, _27289_, _27287_);
  and (_27291_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_27292_, _27291_, rst);
  or (_27293_, _27292_, _27290_);
  or (_24997_, _27293_, _27286_);
  and (_27295_, _27149_, _25972_);
  nand (_27297_, _27295_, _25514_);
  or (_27299_, _27295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_27300_, _27299_, _25521_);
  and (_27302_, _27300_, _27297_);
  nand (_27304_, _27155_, _26475_);
  or (_27306_, _27155_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_27308_, _27306_, _25450_);
  and (_27309_, _27308_, _27304_);
  and (_27310_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_27311_, _27310_, rst);
  or (_27312_, _27311_, _27309_);
  or (_24999_, _27312_, _27302_);
  and (_27313_, _27164_, _25055_);
  nand (_27314_, _27313_, _25514_);
  or (_27315_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_27316_, _27315_, _25521_);
  and (_27317_, _27316_, _27314_);
  nand (_27318_, _27171_, _26521_);
  and (_27319_, _27318_, _25450_);
  and (_27320_, _27319_, _27315_);
  not (_27321_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_27322_, _25449_, _27321_);
  or (_27323_, _27322_, rst);
  or (_27324_, _27323_, _27320_);
  or (_25001_, _27324_, _27317_);
  and (_27325_, _27164_, _26947_);
  nand (_27326_, _27325_, _25514_);
  or (_27327_, _27325_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_27328_, _27327_, _25521_);
  and (_27329_, _27328_, _27326_);
  nand (_27330_, _27171_, _26512_);
  or (_27331_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_27332_, _27331_, _25450_);
  and (_27333_, _27332_, _27330_);
  and (_27334_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_27335_, _27334_, rst);
  or (_27336_, _27335_, _27333_);
  or (_25003_, _27336_, _27329_);
  and (_27337_, _27164_, _25716_);
  nand (_27338_, _27337_, _25514_);
  or (_27339_, _27337_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_27340_, _27339_, _25521_);
  and (_27342_, _27340_, _27338_);
  nand (_27344_, _27171_, _26505_);
  or (_27346_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_27348_, _27346_, _25450_);
  and (_27350_, _27348_, _27344_);
  and (_27352_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_27354_, _27352_, rst);
  or (_27356_, _27354_, _27350_);
  or (_25005_, _27356_, _27342_);
  and (_27358_, _27164_, _25778_);
  nand (_27360_, _27358_, _25514_);
  or (_27361_, _27358_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_27362_, _27361_, _25521_);
  and (_27363_, _27362_, _27360_);
  nand (_27364_, _27171_, _26497_);
  or (_27365_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_27366_, _27365_, _25450_);
  and (_27367_, _27366_, _27364_);
  and (_27368_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_27369_, _27368_, rst);
  or (_27370_, _27369_, _27367_);
  or (_25007_, _27370_, _27363_);
  and (_27371_, _27164_, _25838_);
  nand (_27372_, _27371_, _25514_);
  or (_27373_, _27371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_27374_, _27373_, _25521_);
  and (_27375_, _27374_, _27372_);
  nand (_27376_, _27171_, _26489_);
  or (_27377_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_27378_, _27377_, _25450_);
  and (_27379_, _27378_, _27376_);
  and (_27380_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_27381_, _27380_, rst);
  or (_27382_, _27381_, _27379_);
  or (_25009_, _27382_, _27375_);
  and (_27383_, _27164_, _25905_);
  nand (_27384_, _27383_, _25514_);
  or (_27385_, _27383_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_27386_, _27385_, _25521_);
  and (_27387_, _27386_, _27384_);
  nand (_27388_, _27171_, _26482_);
  or (_27389_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_27390_, _27389_, _25450_);
  and (_27391_, _27390_, _27388_);
  and (_27392_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_27393_, _27392_, rst);
  or (_27394_, _27393_, _27391_);
  or (_25011_, _27394_, _27387_);
  and (_27395_, _27164_, _25972_);
  nand (_27396_, _27395_, _25514_);
  or (_27397_, _27395_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_27398_, _27397_, _25521_);
  and (_27399_, _27398_, _27396_);
  nand (_27400_, _27171_, _26475_);
  or (_27401_, _27171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_27402_, _27401_, _25450_);
  and (_27403_, _27402_, _27400_);
  and (_27404_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_27405_, _27404_, rst);
  or (_27406_, _27405_, _27403_);
  or (_25013_, _27406_, _27399_);
  and (_27407_, _27180_, _25055_);
  nand (_27408_, _27407_, _25514_);
  or (_27409_, _27187_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_27410_, _27409_, _25521_);
  and (_27411_, _27410_, _27408_);
  nand (_27412_, _27187_, _26521_);
  and (_27413_, _27412_, _25450_);
  and (_27414_, _27413_, _27409_);
  not (_27415_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_27416_, _25449_, _27415_);
  or (_27417_, _27416_, rst);
  or (_27418_, _27417_, _27414_);
  or (_25015_, _27418_, _27411_);
  and (_27419_, _27180_, _26947_);
  nand (_27420_, _27419_, _25514_);
  or (_27421_, _27419_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_27422_, _27421_, _25521_);
  and (_27423_, _27422_, _27420_);
  nor (_27424_, _27188_, _26512_);
  and (_27425_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_27426_, _27425_, _27424_);
  and (_27427_, _27426_, _25450_);
  and (_27428_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_27429_, _27428_, rst);
  or (_27430_, _27429_, _27427_);
  or (_25017_, _27430_, _27423_);
  and (_27431_, _27180_, _25716_);
  nand (_27432_, _27431_, _25514_);
  or (_27433_, _27431_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_27434_, _27433_, _25521_);
  and (_27435_, _27434_, _27432_);
  nor (_27436_, _27188_, _26505_);
  and (_27437_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_27438_, _27437_, _27436_);
  and (_27439_, _27438_, _25450_);
  and (_27440_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_27441_, _27440_, rst);
  or (_27442_, _27441_, _27439_);
  or (_25019_, _27442_, _27435_);
  and (_27443_, _27180_, _25778_);
  nand (_27444_, _27443_, _25514_);
  or (_27445_, _27443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_27446_, _27445_, _25521_);
  and (_27447_, _27446_, _27444_);
  nor (_27448_, _27188_, _26497_);
  and (_27449_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_27450_, _27449_, _27448_);
  and (_27451_, _27450_, _25450_);
  and (_27452_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_27453_, _27452_, rst);
  or (_27454_, _27453_, _27451_);
  or (_25021_, _27454_, _27447_);
  and (_27455_, _27180_, _25838_);
  nand (_27456_, _27455_, _25514_);
  or (_27457_, _27455_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_27458_, _27457_, _25521_);
  and (_27459_, _27458_, _27456_);
  nor (_27460_, _27188_, _26489_);
  and (_27461_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_27462_, _27461_, _27460_);
  and (_27463_, _27462_, _25450_);
  and (_27464_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_27465_, _27464_, rst);
  or (_27466_, _27465_, _27463_);
  or (_25023_, _27466_, _27459_);
  and (_27467_, _27180_, _25905_);
  nand (_27468_, _27467_, _25514_);
  or (_27469_, _27467_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_27470_, _27469_, _25521_);
  and (_27471_, _27470_, _27468_);
  nor (_27472_, _27188_, _26482_);
  and (_27473_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_27474_, _27473_, _27472_);
  and (_27475_, _27474_, _25450_);
  and (_27476_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_27477_, _27476_, rst);
  or (_27478_, _27477_, _27475_);
  or (_25025_, _27478_, _27471_);
  and (_27479_, _27180_, _25972_);
  nand (_27480_, _27479_, _25514_);
  or (_27481_, _27479_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_27482_, _27481_, _25521_);
  and (_27483_, _27482_, _27480_);
  nor (_27484_, _27188_, _26475_);
  and (_27485_, _27188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_27486_, _27485_, _27484_);
  and (_27487_, _27486_, _25450_);
  and (_27488_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_27489_, _27488_, rst);
  or (_27490_, _27489_, _27487_);
  or (_25027_, _27490_, _27483_);
  and (_27491_, _27196_, _25055_);
  nand (_27492_, _27491_, _25514_);
  or (_27493_, _27204_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_27494_, _27493_, _25521_);
  and (_27495_, _27494_, _27492_);
  nand (_27496_, _27204_, _26521_);
  and (_27497_, _27496_, _25450_);
  and (_27498_, _27497_, _27493_);
  not (_27499_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_27500_, _25449_, _27499_);
  or (_27501_, _27500_, rst);
  or (_27502_, _27501_, _27498_);
  or (_25029_, _27502_, _27495_);
  and (_27503_, _27196_, _26947_);
  nand (_27504_, _27503_, _25514_);
  or (_27505_, _27503_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_27506_, _27505_, _25521_);
  and (_27507_, _27506_, _27504_);
  nor (_27508_, _27205_, _26512_);
  and (_27509_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_27510_, _27509_, _27508_);
  and (_27511_, _27510_, _25450_);
  and (_27512_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_27513_, _27512_, rst);
  or (_27514_, _27513_, _27511_);
  or (_25031_, _27514_, _27507_);
  and (_27515_, _27196_, _25716_);
  nand (_27516_, _27515_, _25514_);
  or (_27517_, _27515_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_27518_, _27517_, _25521_);
  and (_27519_, _27518_, _27516_);
  nor (_27520_, _27205_, _26505_);
  and (_27521_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_27522_, _27521_, _27520_);
  and (_27523_, _27522_, _25450_);
  and (_27524_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_27525_, _27524_, rst);
  or (_27526_, _27525_, _27523_);
  or (_25033_, _27526_, _27519_);
  and (_27527_, _27196_, _25778_);
  nand (_27528_, _27527_, _25514_);
  or (_27529_, _27527_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_27530_, _27529_, _25521_);
  and (_27531_, _27530_, _27528_);
  nor (_27532_, _27205_, _26497_);
  and (_27533_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_27534_, _27533_, _27532_);
  and (_27535_, _27534_, _25450_);
  and (_27536_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_27537_, _27536_, rst);
  or (_27538_, _27537_, _27535_);
  or (_25035_, _27538_, _27531_);
  and (_27539_, _27196_, _25838_);
  nand (_27540_, _27539_, _25514_);
  or (_27541_, _27539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_27542_, _27541_, _25521_);
  and (_27543_, _27542_, _27540_);
  nor (_27544_, _27205_, _26489_);
  and (_27545_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_27546_, _27545_, _27544_);
  and (_27547_, _27546_, _25450_);
  and (_27548_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_27549_, _27548_, rst);
  or (_27550_, _27549_, _27547_);
  or (_25037_, _27550_, _27543_);
  and (_27551_, _27196_, _25905_);
  nand (_27552_, _27551_, _25514_);
  or (_27553_, _27551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_27554_, _27553_, _25521_);
  and (_27555_, _27554_, _27552_);
  nor (_27556_, _27205_, _26482_);
  and (_27557_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_27558_, _27557_, _27556_);
  and (_27559_, _27558_, _25450_);
  and (_27560_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_27561_, _27560_, rst);
  or (_27562_, _27561_, _27559_);
  or (_25039_, _27562_, _27555_);
  and (_27563_, _27196_, _25972_);
  nand (_27564_, _27563_, _25514_);
  or (_27565_, _27563_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_27566_, _27565_, _25521_);
  and (_27567_, _27566_, _27564_);
  nor (_27568_, _27205_, _26475_);
  and (_27569_, _27205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_27570_, _27569_, _27568_);
  and (_27571_, _27570_, _25450_);
  and (_27572_, _27160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_27573_, _27572_, rst);
  or (_27574_, _27573_, _27571_);
  or (_25041_, _27574_, _27567_);
  and (_25436_, t0_i, _27355_);
  and (_25439_, t1_i, _27355_);
  not (_27575_, _25450_);
  nor (_27576_, _27575_, _25115_);
  and (_27577_, _27576_, _25778_);
  and (_27578_, _27577_, _26460_);
  nand (_27579_, _27578_, _26543_);
  not (_27580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_27581_, _27580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_27582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_27583_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _27582_);
  nor (_27584_, _27583_, _27581_);
  nor (_27585_, _25020_, _25115_);
  and (_27586_, _27585_, _26461_);
  and (_27587_, _27586_, _25450_);
  nor (_27588_, _27587_, _27584_);
  not (_27589_, _27588_);
  and (_27590_, _27589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_27591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_27592_, t1_i);
  and (_27593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _27592_);
  nor (_27594_, _27593_, _27591_);
  not (_27595_, _27594_);
  not (_27596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_27597_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _27596_);
  nor (_27598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_27599_, _27598_);
  and (_27600_, _27599_, _27597_);
  and (_27601_, _27600_, _27595_);
  and (_27602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_27603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_27604_, _27603_, _27602_);
  and (_27605_, _27604_, _27601_);
  and (_27606_, _27605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_27607_, _27606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_27608_, _27607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_27609_, _27608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_27610_, _27604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_27611_, _27610_, _27601_);
  and (_27612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_27613_, _27612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_27614_, _27613_, _27611_);
  nor (_27615_, _27614_, _27584_);
  and (_27616_, _27615_, _27609_);
  and (_27617_, _27614_, _27581_);
  and (_27618_, _27617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_27619_, _27618_, _27616_);
  nor (_27620_, _27619_, _27587_);
  or (_27621_, _27620_, _27590_);
  or (_27622_, _27621_, _27578_);
  and (_27623_, _27622_, _27355_);
  and (_25442_, _27623_, _27579_);
  and (_27624_, _27578_, _27355_);
  and (_27625_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_27626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_27627_, _27626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_27628_, _27627_, _27611_);
  and (_27629_, _27628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_27630_, _27629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_27631_, _27630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_27632_, _27631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_27633_, _27632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_27634_, _27632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_27635_, _27634_, _27613_);
  not (_27636_, _27583_);
  nor (_27637_, _27613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_27638_, _27637_, _27636_);
  nor (_27639_, _27638_, _27635_);
  and (_27640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_27641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_27642_, _27641_);
  nor (_27643_, _27634_, _27642_);
  or (_27644_, _27643_, _27640_);
  or (_27645_, _27644_, _27639_);
  nand (_27646_, _27645_, _27633_);
  nor (_27647_, _27646_, _27587_);
  not (_27648_, _27587_);
  nor (_27649_, _27648_, _26543_);
  or (_27650_, _27649_, _27647_);
  nor (_27651_, _27578_, rst);
  and (_27652_, _27651_, _27650_);
  or (_25445_, _27652_, _27625_);
  not (_27653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_27654_, _27601_, _27653_);
  or (_27655_, _27654_, _27635_);
  and (_27656_, _27655_, _27583_);
  or (_27657_, _27654_, _27634_);
  and (_27658_, _27657_, _27641_);
  nand (_27659_, _27601_, _27580_);
  and (_27660_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_27661_, _27660_, _27659_);
  or (_27662_, _27661_, _27617_);
  or (_27663_, _27662_, _27658_);
  nor (_27664_, _27663_, _27656_);
  nor (_27665_, _27664_, _27587_);
  and (_25448_, _27665_, _27651_);
  and (_27666_, _27576_, _25716_);
  and (_27667_, _27666_, _26460_);
  not (_27668_, _27667_);
  and (_27669_, _27576_, _25838_);
  and (_27670_, _27669_, _26460_);
  nor (_27671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_27672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_27673_, t0_i);
  and (_27674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _27673_);
  nor (_27675_, _27674_, _27672_);
  not (_27676_, _27675_);
  not (_27677_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_27678_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_27679_, _27678_, _27677_);
  and (_27680_, _27679_, _27676_);
  not (_27681_, _27680_);
  and (_27682_, _27681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_27683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_27684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_27685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_27686_, _27685_, _27684_);
  and (_27687_, _27686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_27688_, _27687_, _27680_);
  and (_27689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_27690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_27691_, _27690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_27692_, _27691_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_27693_, _27692_, _27689_);
  and (_27694_, _27693_, _27688_);
  and (_27695_, _27694_, _27683_);
  or (_27696_, _27695_, _27682_);
  and (_27697_, _27696_, _27671_);
  and (_27698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_27699_, _27698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_27700_, _27699_, _27688_);
  not (_27701_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_27702_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _27701_);
  and (_27703_, _27693_, _27683_);
  and (_27704_, _27703_, _27702_);
  or (_27705_, _27704_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_27706_, _27705_, _27700_);
  not (_27707_, _27671_);
  and (_27708_, _27682_, _27707_);
  or (_27709_, _27708_, _27706_);
  or (_27710_, _27709_, _27697_);
  nand (_27711_, _27710_, _27355_);
  nor (_27712_, _27711_, _27670_);
  and (_25451_, _27712_, _27668_);
  nand (_27713_, _27667_, _26543_);
  not (_27714_, _27670_);
  or (_27715_, _27714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_27716_, _27671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_27717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_27718_, _27717_, _27688_);
  or (_27719_, _27718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_27720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_27721_, _27720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand (_27722_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_27723_, _27722_, _27700_);
  and (_27724_, _27723_, _27707_);
  or (_27725_, _27724_, _27670_);
  and (_27726_, _27725_, _27719_);
  or (_27727_, _27726_, _27716_);
  and (_27728_, _27727_, _27715_);
  or (_27729_, _27728_, _27667_);
  and (_27730_, _27729_, _27355_);
  and (_25454_, _27730_, _27713_);
  nand (_27731_, _27670_, _26543_);
  or (_27732_, _27721_, _27702_);
  not (_27733_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_27734_, _27699_, _27687_);
  and (_27735_, _27680_, _27701_);
  and (_27736_, _27735_, _27734_);
  and (_27737_, _27736_, _27693_);
  and (_27738_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_27739_, _27738_, _27733_);
  and (_27740_, _27738_, _27733_);
  or (_27741_, _27740_, _27739_);
  and (_27742_, _27741_, _27732_);
  and (_27743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_27744_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_27745_, _27744_, _27692_);
  and (_27746_, _27745_, _27689_);
  and (_27747_, _27746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_27748_, _27747_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_27749_, _27744_, _27703_);
  and (_27750_, _27749_, _27748_);
  and (_27751_, _27750_, _27743_);
  and (_27752_, _27694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_27753_, _27752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_27754_, _27695_, _27707_);
  and (_27755_, _27754_, _27753_);
  or (_27756_, _27755_, _27751_);
  or (_27757_, _27756_, _27742_);
  or (_27758_, _27757_, _27670_);
  and (_27759_, _27758_, _27668_);
  and (_27760_, _27759_, _27731_);
  and (_27761_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_27762_, _27761_, _27760_);
  and (_25457_, _27762_, _27355_);
  or (_27763_, _27744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_27764_, _27743_, _27355_);
  and (_27765_, _27764_, _27763_);
  not (_27766_, _27744_);
  or (_27767_, _27766_, _27703_);
  nand (_27768_, _27767_, _27765_);
  nor (_27769_, _27768_, _27670_);
  and (_25460_, _27769_, _27668_);
  and (_27770_, _27576_, _26462_);
  or (_27771_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_27772_, _27771_, _27355_);
  nand (_27773_, _27770_, _26543_);
  and (_25463_, _27773_, _27772_);
  nor (_27774_, _26521_, rst);
  or (_27775_, _27774_, _27651_);
  and (_27776_, _27601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_27777_, _27601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_27778_, _27777_, _27776_);
  and (_27779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_27780_, _27779_, _27587_);
  and (_27781_, _27780_, _27778_);
  and (_27782_, _27613_, _27610_);
  and (_27783_, _27782_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_27784_, _27783_, _27581_);
  nor (_27785_, _27784_, _27587_);
  or (_27786_, _27785_, _27578_);
  not (_27787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_27788_, _27780_, _27787_);
  or (_27789_, _27788_, _27786_);
  or (_27790_, _27789_, _27781_);
  and (_26040_, _27790_, _27775_);
  and (_27791_, _27776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_27792_, _27776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_27793_, _27792_, _27791_);
  nand (_27794_, _27793_, _27780_);
  or (_27795_, _27780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_27796_, _27795_, _27794_);
  and (_27797_, _27608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_27798_, _27797_, _27581_);
  nand (_27799_, _27798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_27800_, _27799_, _27587_);
  or (_27801_, _27800_, _27578_);
  or (_27802_, _27801_, _27796_);
  nand (_27803_, _27578_, _26512_);
  and (_27804_, _27803_, _27355_);
  and (_26042_, _27804_, _27802_);
  not (_27805_, _26505_);
  and (_27806_, _27624_, _27805_);
  nor (_27807_, _27791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_27808_, _27776_, _27602_);
  or (_27809_, _27808_, _27807_);
  nand (_27810_, _27809_, _27780_);
  or (_27811_, _27780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_27812_, _27811_, _27810_);
  nand (_27813_, _27798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_27814_, _27813_, _27587_);
  or (_27815_, _27814_, _27812_);
  and (_27816_, _27815_, _27651_);
  or (_26044_, _27816_, _27806_);
  not (_27817_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_27818_, _27780_, _27817_);
  or (_27819_, _27808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_27820_, _27779_, _27605_);
  and (_27821_, _27820_, _27819_);
  and (_27822_, _27617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_27823_, _27822_, _27821_);
  nor (_27824_, _27823_, _27587_);
  or (_27825_, _27824_, _27818_);
  and (_27826_, _27825_, _27651_);
  not (_27827_, _26497_);
  and (_27828_, _27624_, _27827_);
  or (_26046_, _27828_, _27826_);
  not (_27829_, _26489_);
  and (_27830_, _27624_, _27829_);
  and (_27831_, _27617_, _27648_);
  and (_27832_, _27831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_27833_, _27780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_27834_, _27605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_27835_, _27834_, _27611_);
  nand (_27836_, _27835_, _27780_);
  and (_27837_, _27836_, _27833_);
  or (_27838_, _27837_, _27832_);
  and (_27839_, _27838_, _27651_);
  or (_26048_, _27839_, _27830_);
  not (_27840_, _26482_);
  and (_27841_, _27624_, _27840_);
  and (_27842_, _27589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_27843_, _27611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_27844_, _27611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_27845_, _27844_, _27584_);
  and (_27846_, _27845_, _27843_);
  and (_27847_, _27798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_27848_, _27847_, _27846_);
  nor (_27849_, _27848_, _27587_);
  or (_27850_, _27849_, _27842_);
  and (_27851_, _27850_, _27651_);
  or (_26050_, _27851_, _27841_);
  not (_27852_, _26475_);
  and (_27853_, _27624_, _27852_);
  and (_27854_, _27782_, _27601_);
  and (_27855_, _27581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_27856_, _27855_, _27854_);
  nor (_27857_, _27856_, _27587_);
  or (_27858_, _27588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_27859_, _27844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_27860_, _27859_, _27608_);
  nand (_27861_, _27860_, _27588_);
  and (_27862_, _27861_, _27858_);
  or (_27863_, _27862_, _27857_);
  and (_27864_, _27863_, _27651_);
  or (_26052_, _27864_, _27853_);
  and (_27865_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_27866_, _27641_, _27611_);
  and (_27867_, _27854_, _27583_);
  nor (_27868_, _27867_, _27866_);
  and (_27869_, _27868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_27870_, _27868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_27871_, _27870_, _27869_);
  or (_27872_, _27871_, _27587_);
  nand (_27873_, _27587_, _26521_);
  and (_27874_, _27873_, _27651_);
  and (_27875_, _27874_, _27872_);
  or (_26054_, _27875_, _27865_);
  and (_27876_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_27877_, _27587_, _26512_);
  and (_27878_, _27783_, _27601_);
  nor (_27879_, _27878_, _27636_);
  and (_27880_, _27582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_27881_, _27880_, _27611_);
  nor (_27882_, _27881_, _27583_);
  nor (_27883_, _27882_, _27879_);
  or (_27884_, _27883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_27885_, _27883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_27886_, _27885_, _27884_);
  or (_27887_, _27886_, _27587_);
  and (_27888_, _27887_, _27651_);
  and (_27889_, _27888_, _27877_);
  or (_26056_, _27889_, _27876_);
  and (_27890_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_27891_, _27587_, _26505_);
  and (_27892_, _27626_, _27610_);
  and (_27893_, _27892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_27894_, _27893_, _27601_);
  nor (_27895_, _27894_, _27642_);
  or (_27896_, _27895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand (_27897_, _27628_, _27613_);
  and (_27898_, _27897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or (_27899_, _27898_, _27896_);
  and (_27900_, _27899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_27901_, _27867_, _27626_);
  and (_27902_, _27626_, _27641_);
  and (_27903_, _27902_, _27611_);
  nor (_27904_, _27903_, _27901_);
  nor (_27905_, _27904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_27906_, _27905_, _27900_);
  or (_27907_, _27906_, _27587_);
  and (_27908_, _27907_, _27651_);
  and (_27909_, _27908_, _27891_);
  or (_26058_, _27909_, _27890_);
  and (_27910_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_27911_, _27587_, _26497_);
  and (_27912_, _27783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_27913_, _27912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_27914_, _27913_, _27601_);
  and (_27915_, _27914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_27916_, _27914_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_27917_, _27916_, _27583_);
  nor (_27918_, _27917_, _27915_);
  and (_27919_, _27896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_27920_, _27894_, _27641_);
  nor (_27921_, _27920_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_27922_, _27921_, _27919_);
  or (_27923_, _27922_, _27918_);
  or (_27924_, _27923_, _27587_);
  and (_27925_, _27924_, _27651_);
  and (_27926_, _27925_, _27911_);
  or (_26060_, _27926_, _27910_);
  and (_27927_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_27928_, _27587_, _26489_);
  and (_27929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_27930_, _27914_, _27929_);
  or (_27931_, _27915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_27932_, _27931_, _27583_);
  nor (_27933_, _27932_, _27930_);
  and (_27934_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not (_27935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_27936_, _27894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_27937_, _27936_, _27935_);
  or (_27938_, _27936_, _27935_);
  and (_27939_, _27938_, _27937_);
  and (_27940_, _27939_, _27641_);
  or (_27941_, _27940_, _27934_);
  or (_27942_, _27941_, _27933_);
  or (_27943_, _27942_, _27587_);
  and (_27944_, _27943_, _27651_);
  and (_27945_, _27944_, _27928_);
  or (_26062_, _27945_, _27927_);
  and (_27946_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand (_27947_, _27587_, _26482_);
  not (_27948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_27949_, _27630_, _27641_);
  and (_27950_, _27930_, _27583_);
  nor (_27951_, _27950_, _27949_);
  and (_27952_, _27951_, _27948_);
  nor (_27953_, _27951_, _27948_);
  nor (_27954_, _27953_, _27952_);
  or (_27955_, _27954_, _27587_);
  and (_27956_, _27955_, _27651_);
  and (_27957_, _27956_, _27947_);
  or (_26064_, _27957_, _27946_);
  and (_27958_, _27624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_27959_, _27587_, _26475_);
  not (_27960_, _27953_);
  nor (_27961_, _27960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_27962_, _27960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_27963_, _27962_, _27961_);
  or (_27964_, _27963_, _27587_);
  and (_27965_, _27964_, _27651_);
  and (_27966_, _27965_, _27959_);
  or (_26066_, _27966_, _27958_);
  nor (_27967_, _27681_, _27670_);
  or (_27968_, _27967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_27969_, _27680_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_27970_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_27971_, _27970_, _27734_);
  nand (_27972_, _27971_, _27969_);
  or (_27973_, _27972_, _27670_);
  and (_27974_, _27973_, _27968_);
  or (_27975_, _27974_, _27667_);
  nand (_27976_, _27667_, _26521_);
  and (_27977_, _27976_, _27355_);
  and (_26068_, _27977_, _27975_);
  nor (_27978_, _27969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_27979_, _27969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_27980_, _27979_, _27978_);
  and (_27981_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_27982_, _27981_, _27700_);
  nor (_27983_, _27982_, _27980_);
  nor (_27984_, _27983_, _27670_);
  and (_27985_, _27670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_27986_, _27985_, _27984_);
  and (_27987_, _27986_, _27668_);
  nor (_27988_, _27668_, _26512_);
  or (_27989_, _27988_, _27987_);
  and (_26070_, _27989_, _27355_);
  nand (_27990_, _27667_, _26505_);
  nor (_27991_, _27979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_27992_, _27969_, _27684_);
  nor (_27993_, _27992_, _27991_);
  and (_27994_, _27721_, _27700_);
  and (_27995_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_27996_, _27995_, _27993_);
  nor (_27997_, _27996_, _27670_);
  and (_27998_, _27670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_27999_, _27998_, _27997_);
  or (_28000_, _27999_, _27667_);
  and (_28001_, _28000_, _27355_);
  and (_26072_, _28001_, _27990_);
  nand (_28002_, _27667_, _26497_);
  and (_28003_, _27686_, _27680_);
  nor (_28004_, _27992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_28005_, _28004_, _28003_);
  and (_28006_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_28007_, _28006_, _28005_);
  nor (_28008_, _28007_, _27670_);
  and (_28009_, _27670_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_28010_, _28009_, _28008_);
  or (_28011_, _28010_, _27667_);
  and (_28012_, _28011_, _27355_);
  and (_26074_, _28012_, _28002_);
  nor (_28013_, _28003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_28014_, _28013_, _27688_);
  and (_28015_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_28016_, _28015_, _28014_);
  or (_28017_, _28016_, _27670_);
  or (_28018_, _27714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_28019_, _28018_, _27668_);
  and (_28020_, _28019_, _28017_);
  nor (_28021_, _27668_, _26489_);
  or (_28022_, _28021_, _28020_);
  and (_26076_, _28022_, _27355_);
  nand (_28023_, _27667_, _26482_);
  or (_28024_, _27714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_28025_, _27994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_28026_, _27688_, _27707_);
  or (_28027_, _28026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_28028_, _28026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_28029_, _28028_);
  or (_28030_, _28029_, _27670_);
  and (_28031_, _28030_, _28027_);
  or (_28032_, _28031_, _28025_);
  and (_28033_, _28032_, _28024_);
  or (_28034_, _28033_, _27667_);
  and (_28035_, _28034_, _27355_);
  and (_26078_, _28035_, _28023_);
  and (_28036_, _27721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_28037_, _28036_, _27680_);
  and (_28038_, _28037_, _27734_);
  nor (_28039_, _28029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_28040_, _28039_, _28038_);
  nor (_28041_, _28040_, _27670_);
  and (_28042_, _28030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_28043_, _28042_, _28041_);
  and (_28044_, _28043_, _27668_);
  nor (_28045_, _27668_, _26475_);
  or (_28046_, _28045_, _28044_);
  and (_26080_, _28046_, _27355_);
  nor (_28047_, _27736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_28048_, _27736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_28049_, _28048_, _28047_);
  and (_28050_, _28049_, _27732_);
  and (_28051_, _27744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_28052_, _27744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_28053_, _28052_, _27743_);
  nor (_28054_, _28053_, _28051_);
  and (_28055_, _27688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_28056_, _27688_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_28057_, _28056_, _27671_);
  nor (_28058_, _28057_, _28055_);
  or (_28059_, _28058_, _28054_);
  nor (_28060_, _28059_, _28050_);
  nand (_28061_, _28060_, _27714_);
  nand (_28062_, _27670_, _26521_);
  and (_28063_, _28062_, _27668_);
  and (_28064_, _28063_, _28061_);
  and (_28065_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_28066_, _28065_, _28064_);
  and (_26082_, _28066_, _27355_);
  nand (_28067_, _27670_, _26512_);
  or (_28068_, _28048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_28069_, _27734_, _27680_);
  and (_28070_, _28069_, _27690_);
  not (_28071_, _28070_);
  or (_28072_, _28071_, _27721_);
  and (_28073_, _28072_, _27732_);
  and (_28074_, _28073_, _28068_);
  and (_28075_, _27744_, _27690_);
  or (_28076_, _28051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_28077_, _28076_, _27743_);
  nor (_28078_, _28077_, _28075_);
  and (_28079_, _28055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_28080_, _28055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_28081_, _28080_, _27671_);
  nor (_28082_, _28081_, _28079_);
  or (_28083_, _28082_, _28078_);
  or (_28084_, _28083_, _28074_);
  or (_28085_, _28084_, _27670_);
  and (_28086_, _28085_, _27668_);
  and (_28087_, _28086_, _28067_);
  and (_28088_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_28089_, _28088_, _28087_);
  and (_26084_, _28089_, _27355_);
  nand (_28090_, _27670_, _26505_);
  or (_28091_, _28070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_28092_, _28069_, _27691_);
  not (_28093_, _28092_);
  and (_28094_, _28093_, _27702_);
  and (_28095_, _28094_, _28091_);
  or (_28096_, _28079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_28097_, _27691_, _27688_);
  nor (_28098_, _28097_, _27707_);
  and (_28099_, _28098_, _28096_);
  and (_28100_, _28075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_28101_, _28100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_28102_, _27744_, _27691_);
  nand (_28103_, _28102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_28104_, _28103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_28105_, _28104_, _28101_);
  or (_28106_, _28105_, _28099_);
  or (_28107_, _28106_, _28095_);
  or (_28108_, _28107_, _27670_);
  and (_28109_, _28108_, _27668_);
  and (_28110_, _28109_, _28090_);
  and (_28111_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_28112_, _28111_, _28110_);
  and (_26086_, _28112_, _27355_);
  nand (_28113_, _27670_, _26497_);
  not (_28114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_28115_, _28092_, _27701_);
  nor (_28116_, _28115_, _28114_);
  and (_28117_, _28115_, _28114_);
  or (_28118_, _28117_, _28116_);
  and (_28119_, _28118_, _27732_);
  or (_28120_, _28102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_28121_, _27745_);
  and (_28122_, _28121_, _27743_);
  and (_28123_, _28122_, _28120_);
  or (_28124_, _28097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_28125_, _27692_, _27688_);
  nor (_28126_, _28125_, _27707_);
  and (_28127_, _28126_, _28124_);
  or (_28128_, _28127_, _28123_);
  or (_28129_, _28128_, _28119_);
  or (_28130_, _28129_, _27670_);
  and (_28131_, _28130_, _27668_);
  and (_28132_, _28131_, _28113_);
  and (_28133_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_28134_, _28133_, _28132_);
  and (_26088_, _28134_, _27355_);
  nand (_28135_, _27670_, _26489_);
  or (_28136_, _28125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_28137_, _28079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_28138_, _28137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_28139_, _28138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_28140_, _28139_, _27707_);
  and (_28141_, _28140_, _28136_);
  and (_28142_, _28069_, _27692_);
  nand (_28143_, _28142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_28144_, _28142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_28145_, _28144_, _27702_);
  and (_28146_, _28145_, _28143_);
  and (_28147_, _27745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_28148_, _28147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_28149_, _28148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_28150_, _27745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_28151_, _28150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_28152_, _28151_, _28149_);
  or (_28153_, _28152_, _28146_);
  or (_28154_, _28153_, _28141_);
  or (_28155_, _28154_, _27670_);
  and (_28156_, _28155_, _27668_);
  and (_28157_, _28156_, _28135_);
  and (_28158_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_28159_, _28158_, _28157_);
  and (_26090_, _28159_, _27355_);
  nand (_28160_, _27670_, _26482_);
  nor (_28161_, _28143_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_28162_, _28161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_28163_, _28161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_28164_, _28163_, _27732_);
  and (_28165_, _28164_, _28162_);
  not (_28166_, _27746_);
  and (_28167_, _28166_, _27743_);
  or (_28168_, _28150_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_28169_, _28168_, _28167_);
  not (_28170_, _28139_);
  nor (_28171_, _28170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_28172_, _28170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_28173_, _28172_, _28171_);
  and (_28174_, _28173_, _27671_);
  or (_28175_, _28174_, _28169_);
  or (_28176_, _28175_, _28165_);
  or (_28177_, _28176_, _27670_);
  and (_28178_, _28177_, _27668_);
  and (_28179_, _28178_, _28160_);
  and (_28180_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_28181_, _28180_, _28179_);
  and (_26092_, _28181_, _27355_);
  nand (_28182_, _27670_, _26475_);
  or (_28183_, _27737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_28184_, _28183_, _27732_);
  nor (_28185_, _28184_, _27738_);
  or (_28186_, _27746_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_28187_, _27747_);
  and (_28188_, _28187_, _27743_);
  and (_28189_, _28188_, _28186_);
  or (_28190_, _27694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_28191_, _27752_, _27707_);
  and (_28192_, _28191_, _28190_);
  or (_28193_, _28192_, _28189_);
  or (_28194_, _28193_, _28185_);
  or (_28195_, _28194_, _27670_);
  and (_28196_, _28195_, _27668_);
  and (_28197_, _28196_, _28182_);
  and (_28198_, _27667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_28199_, _28198_, _28197_);
  and (_26094_, _28199_, _27355_);
  nor (_28200_, _27770_, _27720_);
  and (_00002_, _27770_, _26522_);
  or (_00003_, _00002_, _28200_);
  and (_26096_, _00003_, _27355_);
  or (_00004_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00005_, _00004_, _27355_);
  nand (_00006_, _27770_, _26512_);
  and (_26098_, _00006_, _00005_);
  or (_00007_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00008_, _00007_, _27355_);
  nand (_00009_, _27770_, _26505_);
  and (_26100_, _00009_, _00008_);
  or (_00010_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_00011_, _00010_, _27355_);
  nand (_00012_, _27770_, _26497_);
  and (_26102_, _00012_, _00011_);
  or (_00013_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00014_, _00013_, _27355_);
  nand (_00015_, _27770_, _26489_);
  and (_26104_, _00015_, _00014_);
  or (_00016_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00017_, _00016_, _27355_);
  nand (_00018_, _27770_, _26482_);
  and (_26106_, _00018_, _00017_);
  or (_00019_, _27770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00020_, _00019_, _27355_);
  nand (_00021_, _27770_, _26475_);
  and (_26108_, _00021_, _00020_);
  nor (_00022_, _25128_, _25115_);
  and (_00023_, _00022_, _27048_);
  and (_00024_, _00023_, _27179_);
  and (_00025_, _00024_, _25517_);
  nand (_00026_, _00025_, _25514_);
  and (_00027_, _26456_, _25517_);
  and (_00028_, _00027_, _27203_);
  not (_00029_, _00028_);
  or (_00030_, _00025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_00031_, _00030_, _00029_);
  and (_00032_, _00031_, _00026_);
  nor (_00033_, _00029_, _26543_);
  or (_00034_, _00033_, _00032_);
  and (_27294_, _00034_, _27355_);
  and (_00035_, _27576_, _25055_);
  and (_00036_, _00035_, _27186_);
  and (_00037_, _25128_, _25116_);
  and (_00038_, _00037_, _27048_);
  and (_00039_, _00038_, _27179_);
  and (_00040_, _00039_, _25517_);
  nand (_00041_, _00040_, _25514_);
  or (_00042_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_00043_, _00042_, _00041_);
  or (_00044_, _00043_, _00036_);
  nand (_00045_, _00036_, _26543_);
  and (_00046_, _00045_, _27355_);
  and (_27296_, _00046_, _00044_);
  and (_00047_, _00035_, _26460_);
  and (_00048_, _00038_, _27147_);
  nand (_00049_, _00048_, _25053_);
  and (_00050_, _00049_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_00051_, _00050_, _00047_);
  nor (_00052_, _27047_, _25115_);
  and (_00053_, _00052_, _25128_);
  and (_00054_, _00053_, _25102_);
  and (_00055_, _00054_, _27147_);
  or (_00056_, _25054_, _25715_);
  and (_00057_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_00058_, _00057_, _27025_);
  and (_00059_, _00058_, _00055_);
  or (_00060_, _00059_, _00051_);
  nand (_00061_, _00047_, _26475_);
  and (_00062_, _00061_, _27355_);
  and (_27298_, _00062_, _00060_);
  not (_00063_, _00047_);
  nor (_00064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_00065_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_00066_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_00067_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_00069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00068_);
  and (_00070_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00071_, _00070_, _00069_);
  nor (_00072_, _00071_, _00067_);
  or (_00073_, _00072_, _00066_);
  and (_00074_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_00075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_00076_, _00075_, _00074_);
  nor (_00077_, _00076_, _00067_);
  and (_00078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00068_);
  and (_00079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00080_, _00079_, _00078_);
  nand (_00081_, _00080_, _00077_);
  or (_00082_, _00081_, _00073_);
  and (_00083_, _00082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_00084_, _00083_, _00065_);
  and (_00085_, _26460_, _25517_);
  and (_00086_, _00085_, _00052_);
  or (_00087_, _00086_, _00084_);
  and (_00088_, _00087_, _00063_);
  nand (_00089_, _00086_, _25514_);
  and (_00090_, _00089_, _00088_);
  nor (_00091_, _00063_, _26543_);
  or (_00092_, _00091_, _00090_);
  and (_27301_, _00092_, _27355_);
  and (_00093_, _27586_, _25521_);
  nand (_00094_, _00093_, _25514_);
  not (_00095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_00096_, _00095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_00097_, _00080_, _00067_);
  not (_00098_, _00097_);
  or (_00099_, _00098_, _00077_);
  or (_00100_, _00099_, _00073_);
  and (_00101_, _00100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_00102_, _00101_, _00096_);
  or (_00103_, _00102_, _00093_);
  and (_00104_, _00103_, _00063_);
  and (_00105_, _00104_, _00094_);
  nor (_00106_, _00063_, _26482_);
  or (_00107_, _00106_, _00105_);
  and (_27303_, _00107_, _27355_);
  not (_00108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_00109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _00108_);
  nand (_00110_, _00072_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_00111_, _00097_, _00077_);
  or (_00112_, _00111_, _00110_);
  and (_00113_, _00112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_00114_, _00113_, _00109_);
  and (_00115_, _00052_, _26462_);
  or (_00116_, _00115_, _00114_);
  and (_00117_, _00116_, _00063_);
  nand (_00118_, _00115_, _25514_);
  and (_00119_, _00118_, _00117_);
  nor (_00120_, _00063_, _26512_);
  or (_00121_, _00120_, _00119_);
  and (_27305_, _00121_, _27355_);
  and (_00122_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_00123_, _00110_, _00099_);
  and (_00124_, _00123_, _00122_);
  and (_00125_, _00052_, _26592_);
  or (_00126_, _00125_, _00124_);
  and (_00127_, _00126_, _00063_);
  nand (_00128_, _00125_, _25514_);
  and (_00129_, _00128_, _00127_);
  nor (_00130_, _00063_, _26497_);
  or (_00131_, _00130_, _00129_);
  and (_27307_, _00131_, _27355_);
  nand (_00132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_00133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00068_);
  and (_00134_, _00133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_00135_, _00134_, _00132_);
  or (_00136_, _00135_, _00067_);
  and (_00137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_00138_, _00137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_00139_, _00138_);
  and (_00140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_00141_, _00140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_00143_, _00141_);
  and (_00145_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_00147_, _00145_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_00151_, _00149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_00153_, _00151_, _00147_);
  and (_00155_, _00153_, _00143_);
  and (_00157_, _00155_, _00139_);
  not (_00159_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_00161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_00163_, _00161_, _00159_);
  nand (_00165_, _00163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_00167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_00171_, _00169_, _00167_);
  and (_00173_, _00171_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_00175_, _00173_);
  and (_00177_, _00175_, _00165_);
  nand (_00179_, _00177_, _00157_);
  and (_00181_, _00179_, _00136_);
  and (_00183_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_00185_, _00183_, _00068_);
  and (_00187_, _00185_, _00181_);
  not (_00189_, _00187_);
  not (_00191_, _00185_);
  and (_00193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _00067_);
  not (_00195_, _00193_);
  not (_00197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_00199_, _00140_, _00197_);
  not (_00201_, _00199_);
  not (_00203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00204_, _00145_, _00203_);
  not (_00205_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_00206_, _00149_, _00205_);
  nor (_00207_, _00206_, _00204_);
  and (_00208_, _00207_, _00201_);
  nor (_00209_, _00208_, _00195_);
  not (_00210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_00211_, _00163_, _00210_);
  not (_00212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_00213_, _00171_, _00212_);
  nor (_00214_, _00213_, _00211_);
  not (_00215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_00216_, _00137_, _00215_);
  not (_00217_, _00216_);
  and (_00218_, _00217_, _00214_);
  nor (_00219_, _00218_, _00195_);
  nor (_00220_, _00219_, _00209_);
  or (_00221_, _00220_, _00191_);
  and (_00222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _27355_);
  and (_00223_, _00222_, _00221_);
  and (_27341_, _00223_, _00189_);
  nor (_00224_, _00183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_00225_, _00224_);
  not (_00226_, _00181_);
  and (_00227_, _00220_, _00226_);
  nor (_00228_, _00227_, _00225_);
  nand (_00229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _27355_);
  nor (_27343_, _00229_, _00228_);
  and (_00230_, _00177_, _00139_);
  nand (_00231_, _00230_, _00181_);
  or (_00232_, _00219_, _00181_);
  and (_00233_, _00232_, _00185_);
  and (_00234_, _00233_, _00231_);
  or (_00235_, _00234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_00236_, _00189_, _00155_);
  nor (_00237_, _00191_, _00181_);
  nand (_00238_, _00237_, _00209_);
  and (_00239_, _00238_, _27355_);
  and (_00240_, _00239_, _00236_);
  and (_27345_, _00240_, _00235_);
  and (_00241_, _00231_, _00224_);
  or (_00242_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_00243_, _00224_, _00181_);
  not (_00244_, _00243_);
  or (_00245_, _00244_, _00155_);
  or (_00246_, _00219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_00247_, _00224_, _00209_);
  and (_00248_, _00247_, _00246_);
  or (_00249_, _00248_, _00181_);
  and (_00250_, _00249_, _27355_);
  and (_00251_, _00250_, _00245_);
  and (_27347_, _00251_, _00242_);
  nand (_00252_, _00227_, _00067_);
  nor (_00253_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_00254_, _00253_, _00183_);
  and (_00255_, _00254_, _27355_);
  and (_27349_, _00255_, _00252_);
  and (_00256_, _00227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_00257_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_00258_, _00257_, _00253_);
  nor (_00259_, _00258_, _00226_);
  or (_00260_, _00259_, _00183_);
  or (_00261_, _00260_, _00256_);
  not (_00262_, _00183_);
  or (_00263_, _00258_, _00262_);
  and (_00264_, _00263_, _27355_);
  and (_27351_, _00264_, _00261_);
  and (_00265_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _27355_);
  and (_27353_, _00265_, _00183_);
  nor (_27357_, _00064_, rst);
  and (_27359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _27355_);
  nor (_00266_, _00227_, _00183_);
  and (_00267_, _00183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_00268_, _00267_, _00266_);
  and (_00142_, _00268_, _27355_);
  and (_00269_, _00183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_00270_, _00269_, _00266_);
  and (_00144_, _00270_, _27355_);
  and (_00271_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _27355_);
  and (_00146_, _00271_, _00183_);
  nor (_00272_, _00220_, _00181_);
  not (_00273_, _00206_);
  nor (_00274_, _00213_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_00275_, _00274_, _00211_);
  or (_00276_, _00275_, _00216_);
  and (_00277_, _00276_, _00273_);
  or (_00278_, _00277_, _00204_);
  and (_00279_, _00278_, _00201_);
  and (_00280_, _00279_, _00272_);
  not (_00281_, _00151_);
  or (_00282_, _00173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_00283_, _00282_, _00165_);
  or (_00284_, _00283_, _00138_);
  and (_00285_, _00284_, _00281_);
  or (_00286_, _00285_, _00147_);
  and (_00287_, _00181_, _00143_);
  and (_00288_, _00287_, _00286_);
  or (_00289_, _00288_, _00183_);
  or (_00290_, _00289_, _00280_);
  or (_00291_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_00292_, _00291_, _27355_);
  and (_00148_, _00292_, _00290_);
  nor (_00293_, _00204_, _00199_);
  or (_00294_, _00216_, _00206_);
  and (_00295_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_00296_, _00295_, _00294_);
  and (_00297_, _00296_, _00293_);
  and (_00298_, _00297_, _00272_);
  not (_00299_, _00147_);
  or (_00300_, _00151_, _00138_);
  and (_00301_, _00177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_00302_, _00301_, _00300_);
  and (_00303_, _00302_, _00299_);
  and (_00304_, _00303_, _00287_);
  or (_00305_, _00304_, _00183_);
  or (_00306_, _00305_, _00298_);
  or (_00307_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_00308_, _00307_, _27355_);
  and (_00150_, _00308_, _00306_);
  and (_00309_, _00217_, _00193_);
  nand (_00310_, _00309_, _00208_);
  or (_00311_, _00310_, _00214_);
  nor (_00312_, _00311_, _00181_);
  nand (_00313_, _00157_, _00136_);
  nor (_00314_, _00313_, _00177_);
  or (_00315_, _00314_, _00183_);
  or (_00316_, _00315_, _00312_);
  or (_00317_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_00318_, _00317_, _27355_);
  and (_00152_, _00318_, _00316_);
  and (_00319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _27355_);
  and (_00154_, _00319_, _00183_);
  and (_00320_, _00183_, _00068_);
  or (_00321_, _00320_, _00228_);
  or (_00322_, _00321_, _00237_);
  and (_00156_, _00322_, _27355_);
  not (_00323_, _00266_);
  and (_00324_, _00323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_00325_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00068_);
  or (_00326_, _00325_, _00143_);
  and (_00327_, _00326_, _00181_);
  not (_00328_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_00329_, _00173_, _00068_);
  or (_00330_, _00329_, _00328_);
  nor (_00331_, _00165_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00332_, _00331_, _00138_);
  nand (_00333_, _00332_, _00330_);
  or (_00334_, _00139_, _00070_);
  and (_00335_, _00334_, _00333_);
  or (_00336_, _00335_, _00151_);
  or (_00337_, _00325_, _00281_);
  and (_00338_, _00337_, _00299_);
  and (_00339_, _00338_, _00336_);
  and (_00340_, _00147_, _00070_);
  or (_00341_, _00340_, _00141_);
  or (_00342_, _00341_, _00339_);
  and (_00343_, _00342_, _00327_);
  or (_00344_, _00325_, _00201_);
  and (_00345_, _00213_, _00068_);
  or (_00346_, _00345_, _00328_);
  and (_00347_, _00211_, _00068_);
  nor (_00348_, _00347_, _00216_);
  nand (_00349_, _00348_, _00346_);
  or (_00350_, _00217_, _00070_);
  and (_00351_, _00350_, _00349_);
  or (_00352_, _00351_, _00206_);
  not (_00353_, _00204_);
  or (_00354_, _00325_, _00273_);
  and (_00355_, _00354_, _00353_);
  and (_00356_, _00355_, _00352_);
  and (_00357_, _00204_, _00070_);
  or (_00358_, _00357_, _00199_);
  or (_00359_, _00358_, _00356_);
  and (_00360_, _00359_, _00272_);
  and (_00361_, _00360_, _00344_);
  or (_00362_, _00361_, _00343_);
  and (_00363_, _00362_, _00262_);
  or (_00364_, _00363_, _00324_);
  and (_00158_, _00364_, _27355_);
  or (_00365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00068_);
  and (_00366_, _00365_, _00143_);
  or (_00367_, _00366_, _00155_);
  or (_00368_, _00329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_00369_, _00368_, _00332_);
  nand (_00370_, _00138_, _00079_);
  nand (_00371_, _00370_, _00153_);
  or (_00372_, _00371_, _00369_);
  and (_00373_, _00372_, _00367_);
  nand (_00374_, _00141_, _00079_);
  nand (_00375_, _00374_, _00181_);
  or (_00376_, _00375_, _00373_);
  or (_00377_, _00345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_00378_, _00377_, _00348_);
  and (_00379_, _00216_, _00079_);
  or (_00380_, _00379_, _00378_);
  and (_00381_, _00380_, _00207_);
  not (_00382_, _00207_);
  and (_00383_, _00365_, _00382_);
  or (_00384_, _00383_, _00199_);
  or (_00385_, _00384_, _00381_);
  or (_00386_, _00201_, _00079_);
  nand (_00387_, _00386_, _00385_);
  nand (_00388_, _00387_, _00272_);
  and (_00389_, _00388_, _00376_);
  or (_00390_, _00389_, _00183_);
  or (_00391_, _00266_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_00392_, _00391_, _27355_);
  and (_00160_, _00392_, _00390_);
  and (_00393_, _00323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_00394_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00395_, _00394_, _00143_);
  and (_00396_, _00395_, _00181_);
  not (_00397_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_00398_, _00173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00399_, _00398_, _00397_);
  nor (_00400_, _00165_, _00068_);
  nor (_00401_, _00400_, _00138_);
  nand (_00402_, _00401_, _00399_);
  or (_00403_, _00139_, _00069_);
  and (_00404_, _00403_, _00402_);
  or (_00405_, _00404_, _00151_);
  or (_00406_, _00394_, _00281_);
  and (_00407_, _00406_, _00299_);
  and (_00408_, _00407_, _00405_);
  and (_00409_, _00147_, _00069_);
  or (_00410_, _00409_, _00141_);
  or (_00411_, _00410_, _00408_);
  and (_00412_, _00411_, _00396_);
  or (_00413_, _00394_, _00201_);
  and (_00414_, _00213_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00415_, _00414_, _00397_);
  and (_00416_, _00211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00417_, _00416_, _00216_);
  nand (_00418_, _00417_, _00415_);
  or (_00419_, _00217_, _00069_);
  and (_00420_, _00419_, _00418_);
  or (_00421_, _00420_, _00206_);
  or (_00422_, _00394_, _00273_);
  and (_00423_, _00422_, _00353_);
  and (_00424_, _00423_, _00421_);
  and (_00425_, _00204_, _00069_);
  or (_00426_, _00425_, _00199_);
  or (_00427_, _00426_, _00424_);
  and (_00428_, _00427_, _00272_);
  and (_00429_, _00428_, _00413_);
  or (_00430_, _00429_, _00412_);
  and (_00431_, _00430_, _00262_);
  or (_00432_, _00431_, _00393_);
  and (_00162_, _00432_, _27355_);
  and (_00433_, _00199_, _00078_);
  or (_00434_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_00435_, _00434_, _00201_);
  or (_00436_, _00435_, _00208_);
  and (_00437_, _00216_, _00078_);
  or (_00438_, _00414_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00439_, _00438_, _00417_);
  or (_00440_, _00439_, _00382_);
  or (_00441_, _00440_, _00437_);
  and (_00442_, _00441_, _00436_);
  or (_00443_, _00442_, _00433_);
  and (_00444_, _00443_, _00272_);
  or (_00445_, _00398_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00446_, _00445_, _00401_);
  and (_00447_, _00138_, _00078_);
  or (_00448_, _00447_, _00446_);
  and (_00449_, _00448_, _00153_);
  not (_00450_, _00153_);
  and (_00451_, _00434_, _00450_);
  or (_00452_, _00451_, _00141_);
  or (_00453_, _00452_, _00449_);
  or (_00454_, _00143_, _00078_);
  and (_00455_, _00454_, _00181_);
  and (_00456_, _00455_, _00453_);
  and (_00457_, _00227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_00458_, _00457_, _00183_);
  or (_00459_, _00458_, _00456_);
  or (_00460_, _00459_, _00444_);
  or (_00461_, _00262_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00462_, _00461_, _27355_);
  and (_00164_, _00462_, _00460_);
  or (_00463_, _00225_, _00220_);
  and (_00464_, _00463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_00465_, _00464_, _00243_);
  and (_00166_, _00465_, _27355_);
  and (_00466_, _00221_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_00467_, _00466_, _00187_);
  and (_00168_, _00467_, _27355_);
  or (_00468_, _00049_, _25719_);
  or (_00469_, _00468_, _25574_);
  nand (_00470_, _00468_, _00108_);
  and (_00471_, _00470_, _00063_);
  and (_00472_, _00471_, _00469_);
  nor (_00473_, _00063_, _26521_);
  or (_00474_, _00473_, _00472_);
  and (_00170_, _00474_, _27355_);
  nand (_00475_, _00055_, _25716_);
  nor (_00476_, _00475_, _25514_);
  and (_00477_, _00475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_00478_, _00477_, _00047_);
  or (_00479_, _00478_, _00476_);
  nand (_00480_, _00047_, _26505_);
  and (_00481_, _00480_, _27355_);
  and (_00172_, _00481_, _00479_);
  and (_00482_, _00055_, _25838_);
  or (_00483_, _00482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_00484_, _00483_, _00063_);
  nand (_00485_, _00482_, _25514_);
  and (_00486_, _00485_, _00484_);
  nor (_00487_, _00063_, _26489_);
  or (_00488_, _00487_, _00486_);
  and (_00174_, _00488_, _27355_);
  and (_00489_, _00039_, _25055_);
  nand (_00490_, _00489_, _25514_);
  not (_00491_, _00036_);
  or (_00492_, _00489_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_00493_, _00492_, _00491_);
  and (_00494_, _00493_, _00490_);
  nor (_00495_, _00491_, _26521_);
  or (_00496_, _00495_, _00494_);
  and (_00176_, _00496_, _27355_);
  and (_00497_, _00039_, _26947_);
  or (_00498_, _00497_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_00499_, _00498_, _00491_);
  nand (_00500_, _00497_, _25514_);
  and (_00501_, _00500_, _00499_);
  nor (_00502_, _00491_, _26512_);
  or (_00503_, _00502_, _00501_);
  and (_00178_, _00503_, _27355_);
  nand (_00504_, _00039_, _27237_);
  and (_00505_, _00504_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00506_, _00505_, _00036_);
  and (_00507_, _27240_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00508_, _00507_, _25718_);
  and (_00509_, _00508_, _00039_);
  or (_00510_, _00509_, _00506_);
  nand (_00511_, _00036_, _26505_);
  and (_00512_, _00511_, _27355_);
  and (_00180_, _00512_, _00510_);
  and (_00513_, _00039_, _25778_);
  or (_00514_, _00513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_00515_, _00514_, _00491_);
  nand (_00516_, _00513_, _25514_);
  and (_00517_, _00516_, _00515_);
  nor (_00518_, _00491_, _26497_);
  or (_00519_, _00518_, _00517_);
  and (_00182_, _00519_, _27355_);
  and (_00520_, _00039_, _25838_);
  nand (_00521_, _00520_, _25514_);
  or (_00522_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_00523_, _00522_, _00521_);
  or (_00524_, _00523_, _00036_);
  nand (_00525_, _00036_, _26489_);
  and (_00526_, _00525_, _27355_);
  and (_00184_, _00526_, _00524_);
  and (_00527_, _00039_, _25905_);
  or (_00528_, _00527_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_00529_, _00528_, _00491_);
  nand (_00530_, _00527_, _25514_);
  and (_00531_, _00530_, _00529_);
  nor (_00532_, _00491_, _26482_);
  or (_00533_, _00532_, _00531_);
  and (_00186_, _00533_, _27355_);
  and (_00534_, _00039_, _25972_);
  or (_00535_, _00534_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_00536_, _00535_, _00491_);
  nand (_00537_, _00534_, _25514_);
  and (_00538_, _00537_, _00536_);
  nor (_00539_, _00491_, _26475_);
  or (_00540_, _00539_, _00538_);
  and (_00188_, _00540_, _27355_);
  and (_00541_, _00024_, _25055_);
  nand (_00542_, _00541_, _25514_);
  or (_00543_, _00541_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_00544_, _00028_, rst);
  and (_00545_, _00544_, _00543_);
  and (_00546_, _00545_, _00542_);
  and (_00547_, _00028_, _27774_);
  or (_00190_, _00547_, _00546_);
  and (_00548_, _00024_, _26947_);
  nand (_00549_, _00548_, _25514_);
  or (_00550_, _00548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00551_, _00550_, _00029_);
  and (_00552_, _00551_, _00549_);
  nor (_00553_, _00029_, _26512_);
  or (_00554_, _00553_, _00552_);
  and (_00192_, _00554_, _27355_);
  nor (_00555_, _25719_, _00205_);
  or (_00556_, _00555_, _25718_);
  and (_00557_, _00556_, _00024_);
  nand (_00558_, _00024_, _27237_);
  and (_00559_, _00558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_00560_, _00559_, _00028_);
  or (_00561_, _00560_, _00557_);
  nand (_00562_, _00028_, _26505_);
  and (_00563_, _00562_, _27355_);
  and (_00194_, _00563_, _00561_);
  and (_00564_, _00024_, _25778_);
  nand (_00565_, _00564_, _25514_);
  or (_00566_, _00564_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_00567_, _00566_, _00565_);
  or (_00568_, _00567_, _00028_);
  nand (_00569_, _00028_, _26497_);
  and (_00570_, _00569_, _27355_);
  and (_00196_, _00570_, _00568_);
  and (_00571_, _00024_, _25838_);
  nand (_00572_, _00571_, _25514_);
  or (_00573_, _00571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_00574_, _00573_, _00572_);
  or (_00575_, _00574_, _00028_);
  nand (_00576_, _00028_, _26489_);
  and (_00577_, _00576_, _27355_);
  and (_00198_, _00577_, _00575_);
  and (_00578_, _00024_, _25905_);
  nand (_00579_, _00578_, _25514_);
  or (_00580_, _00578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_00581_, _00580_, _00579_);
  or (_00582_, _00581_, _00028_);
  nand (_00583_, _00028_, _26482_);
  and (_00584_, _00583_, _27355_);
  and (_00200_, _00584_, _00582_);
  and (_00585_, _00024_, _25972_);
  nand (_00586_, _00585_, _25514_);
  or (_00588_, _00585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_00589_, _00588_, _00029_);
  and (_00591_, _00589_, _00586_);
  nor (_00592_, _00029_, _26475_);
  or (_00594_, _00592_, _00591_);
  and (_00202_, _00594_, _27355_);
  and (_00596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_00597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_00599_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_00600_, _00599_, _00597_);
  not (_00602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_00603_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_00605_, _00603_, _00600_);
  nor (_00606_, _00605_, _00596_);
  or (_00608_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_00609_, _00608_, _27355_);
  nor (_00590_, _00609_, _00606_);
  nor (_00611_, _00606_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_00613_, _00611_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_00614_, _00611_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_00616_, _00614_, _27355_);
  and (_00593_, _00616_, _00613_);
  not (_00618_, rxd_i);
  and (_00619_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00618_);
  nor (_00621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_00622_, _00621_);
  and (_00624_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_00625_, _00624_, _00622_);
  and (_00627_, _00625_, _00619_);
  not (_00628_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_00630_, _00628_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_00631_, _00630_, _00621_);
  or (_00633_, _00631_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_00634_, _00633_, _00627_);
  and (_00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _27355_);
  and (_00595_, _00636_, _00634_);
  and (_00638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_00639_, _00638_, _00622_);
  nor (_00640_, _00621_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_00641_, _00640_, _00628_);
  nor (_00642_, _00641_, _00639_);
  not (_00643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_00644_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _00643_);
  not (_00645_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_00646_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _00645_);
  and (_00647_, _00646_, _00644_);
  not (_00648_, _00647_);
  or (_00649_, _00648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_00650_, _00647_, _00639_);
  and (_00651_, _00639_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00652_, _00651_, _00650_);
  and (_00653_, _00652_, _00649_);
  or (_00654_, _00653_, _00642_);
  and (_00655_, _00621_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_00656_, _00655_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not (_00657_, _00656_);
  or (_00658_, _00657_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_00659_, _00658_, _00654_);
  nand (_00598_, _00659_, _00636_);
  not (_00660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_00661_, _00639_);
  nor (_00662_, _00628_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_00663_, _00662_);
  not (_00664_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_00665_, _00621_, _00664_);
  and (_00666_, _00665_, _00663_);
  and (_00667_, _00666_, _00661_);
  nor (_00668_, _00667_, _00660_);
  and (_00669_, _00667_, rxd_i);
  or (_00670_, _00669_, rst);
  or (_00601_, _00670_, _00668_);
  nor (_00671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_00672_, _00671_, _00644_);
  and (_00673_, _00672_, _00651_);
  nand (_00674_, _00673_, _00618_);
  or (_00675_, _00673_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_00676_, _00675_, _27355_);
  and (_00604_, _00676_, _00674_);
  and (_00677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_00678_, _00677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_00679_, _00678_, _00643_);
  and (_00680_, _00679_, _00651_);
  and (_00681_, _00625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_00682_, _00681_, _00651_);
  nor (_00683_, _00678_, _00661_);
  or (_00684_, _00683_, _00682_);
  and (_00685_, _00684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_00686_, _00685_, _00680_);
  and (_00607_, _00686_, _27355_);
  and (_00687_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _27355_);
  nand (_00688_, _00687_, _00664_);
  nand (_00689_, _00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_00610_, _00689_, _00688_);
  and (_00690_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00664_);
  not (_00691_, _00625_);
  not (_00692_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_00693_, _00631_, _00692_);
  and (_00694_, _00693_, _00691_);
  and (_00695_, _00694_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_00696_, _00695_, _00639_);
  or (_00697_, _00647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_00698_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_00699_, _00698_, _00650_);
  and (_00700_, _00699_, _00697_);
  and (_00701_, _00700_, _00696_);
  or (_00702_, _00701_, _00656_);
  nand (_00703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_00704_, _00703_, _00639_);
  or (_00705_, _00704_, _00648_);
  and (_00706_, _00705_, _00657_);
  or (_00707_, _00706_, rxd_i);
  and (_00708_, _00707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_00709_, _00708_, _00702_);
  or (_00710_, _00709_, _00690_);
  and (_00612_, _00710_, _27355_);
  and (_00711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_00712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_00713_, _00599_, _00712_);
  or (_00714_, _00713_, _00603_);
  nor (_00715_, _00714_, _00711_);
  or (_00716_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_00717_, _00716_, _27355_);
  nor (_00615_, _00717_, _00715_);
  nor (_00718_, _00715_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_00719_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_00720_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_00721_, _00720_, _27355_);
  and (_00617_, _00721_, _00719_);
  and (_00722_, _00655_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_00723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_00724_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_00725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_00726_, _00725_, _00724_);
  and (_00727_, _00726_, _00723_);
  not (_00728_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_00729_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_00730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_00731_, _00730_, _00729_);
  and (_00732_, _00731_, _00728_);
  and (_00733_, _00732_, _00727_);
  or (_00734_, _00733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_00735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_00736_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_00737_, _00736_, _00735_);
  and (_00738_, _00622_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_00739_, _00738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_00740_, _00739_, _00737_);
  not (_00741_, _00740_);
  or (_00742_, _00741_, _00734_);
  and (_00743_, _00737_, _00738_);
  not (_00744_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or (_00745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00744_);
  or (_00746_, _00745_, _00743_);
  and (_00747_, _00746_, _00742_);
  or (_00748_, _00747_, _00722_);
  not (_00749_, _00722_);
  not (_00750_, _00733_);
  or (_00751_, _00750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_00752_, _00751_, _00734_);
  or (_00753_, _00752_, _00749_);
  nand (_00754_, _00753_, _00748_);
  nand (_00755_, _26947_, _25116_);
  nor (_00756_, _00755_, _27575_);
  and (_00757_, _00756_, _27170_);
  nor (_00758_, _00757_, rst);
  nand (_00759_, _00758_, _00754_);
  not (_00760_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_00761_, _00757_, _27355_);
  nand (_00762_, _00761_, _00760_);
  and (_00620_, _00762_, _00759_);
  nor (_00763_, _00750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_00764_, _00743_, _00763_);
  and (_00765_, _00733_, _00722_);
  or (_00766_, _00744_, rst);
  nor (_00767_, _00766_, _00765_);
  and (_00768_, _00767_, _00764_);
  or (_00623_, _00768_, _00761_);
  or (_00769_, _00741_, _00763_);
  or (_00770_, _00743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_00771_, _00655_, _00744_);
  and (_00772_, _00771_, _00770_);
  and (_00773_, _00772_, _00769_);
  or (_00774_, _00773_, _00765_);
  and (_00626_, _00774_, _00758_);
  and (_00775_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_00776_, _00775_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_00777_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_00779_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_00780_, _00779_, _00778_);
  and (_00629_, _00780_, _00758_);
  nor (_00781_, _00740_, _00722_);
  and (_00782_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_00783_, _00782_, _00758_);
  and (_00784_, _00761_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_00632_, _00784_, _00783_);
  and (_00785_, _00027_, _26460_);
  or (_00786_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_00787_, _00786_, _27355_);
  nand (_00788_, _00785_, _26543_);
  and (_00635_, _00788_, _00787_);
  and (_00789_, _00023_, _27147_);
  and (_00790_, _00789_, _25517_);
  nand (_00791_, _00790_, _25514_);
  and (_00792_, _00035_, _27170_);
  not (_00793_, _00792_);
  or (_00794_, _00790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_00795_, _00794_, _00793_);
  and (_00796_, _00795_, _00791_);
  nor (_00797_, _00793_, _26543_);
  or (_00798_, _00797_, _00796_);
  and (_00637_, _00798_, _27355_);
  nor (_00799_, _00656_, _00650_);
  not (_00800_, _00799_);
  nor (_00801_, _00694_, _00639_);
  nor (_00802_, _00801_, _00800_);
  nor (_00803_, _00802_, _00664_);
  or (_00804_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_00805_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _00664_);
  or (_00806_, _00805_, _00799_);
  and (_00807_, _00806_, _27355_);
  and (_01239_, _00807_, _00804_);
  or (_00808_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_00809_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _00664_);
  or (_00810_, _00809_, _00799_);
  and (_00811_, _00810_, _27355_);
  and (_01241_, _00811_, _00808_);
  or (_00812_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_00813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _00664_);
  or (_00814_, _00813_, _00799_);
  and (_00815_, _00814_, _27355_);
  and (_01243_, _00815_, _00812_);
  or (_00816_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_00817_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _00664_);
  or (_00818_, _00817_, _00799_);
  and (_00819_, _00818_, _27355_);
  and (_01245_, _00819_, _00816_);
  or (_00820_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_00821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _00664_);
  or (_00822_, _00821_, _00799_);
  and (_00823_, _00822_, _27355_);
  and (_01247_, _00823_, _00820_);
  or (_00824_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_00825_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _00664_);
  or (_00826_, _00825_, _00799_);
  and (_00827_, _00826_, _27355_);
  and (_01248_, _00827_, _00824_);
  or (_00828_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_00829_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _00664_);
  or (_00830_, _00829_, _00799_);
  and (_00831_, _00830_, _27355_);
  and (_01250_, _00831_, _00828_);
  or (_00832_, _00803_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_00833_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _00664_);
  or (_00834_, _00833_, _00799_);
  and (_00835_, _00834_, _27355_);
  and (_01252_, _00835_, _00832_);
  nor (_00836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_00837_, _00836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_00838_, _00648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_00839_, _00647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_00840_, _00839_, _00639_);
  and (_00841_, _00840_, _00838_);
  or (_00842_, _00625_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_00843_, _00842_, _00693_);
  and (_00844_, _00843_, _00661_);
  or (_00845_, _00844_, _00841_);
  or (_00846_, _00845_, _00656_);
  or (_00847_, _00657_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_00848_, _00847_, _00636_);
  and (_00849_, _00848_, _00846_);
  or (_01254_, _00849_, _00837_);
  and (_00850_, _00647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_00851_, _00850_, _00694_);
  or (_00852_, _00851_, _00802_);
  and (_00853_, _00852_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_00854_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _00664_);
  nand (_00855_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_00856_, _00855_, _00799_);
  or (_00857_, _00856_, _00854_);
  or (_00858_, _00857_, _00853_);
  and (_01256_, _00858_, _27355_);
  not (_00859_, _00803_);
  and (_00860_, _00859_, _00687_);
  or (_00861_, _00851_, _00800_);
  and (_00862_, _00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_00863_, _00862_, _00861_);
  or (_01258_, _00863_, _00860_);
  or (_00864_, _00680_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_00865_, _00680_, _00618_);
  and (_00866_, _00865_, _27355_);
  and (_01260_, _00866_, _00864_);
  or (_00867_, _00682_, _00645_);
  or (_00868_, _00651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_00869_, _00868_, _27355_);
  and (_01262_, _00869_, _00867_);
  and (_00870_, _00682_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_00871_, _00671_, _00677_);
  and (_00872_, _00871_, _00651_);
  or (_00873_, _00872_, _00870_);
  and (_01264_, _00873_, _27355_);
  and (_00874_, _00684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_00875_, _00677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_00876_, _00875_, _00683_);
  or (_00877_, _00876_, _00874_);
  and (_01266_, _00877_, _27355_);
  and (_00878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _00664_);
  and (_00879_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00880_, _00879_, _00878_);
  and (_01267_, _00880_, _27355_);
  and (_00881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _00664_);
  and (_00882_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00883_, _00882_, _00881_);
  and (_01269_, _00883_, _27355_);
  and (_00884_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _00664_);
  and (_00885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00886_, _00885_, _00884_);
  and (_01271_, _00886_, _27355_);
  and (_00887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _00664_);
  and (_00888_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00889_, _00888_, _00887_);
  and (_01273_, _00889_, _27355_);
  and (_00890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _00664_);
  and (_00891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00892_, _00891_, _00890_);
  and (_01275_, _00892_, _27355_);
  and (_00893_, _00636_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01277_, _00893_, _00837_);
  and (_00894_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00895_, _00894_, _00854_);
  and (_01279_, _00895_, _27355_);
  nor (_00896_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_00897_, _00896_, _00775_);
  and (_01281_, _00897_, _00758_);
  nor (_00898_, _00775_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_00899_, _00898_, _00776_);
  and (_01282_, _00899_, _00758_);
  nor (_00900_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_00901_, _00900_, _00777_);
  and (_01284_, _00901_, _00758_);
  or (_00902_, _00740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_00903_, _00741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_00904_, _00903_, _00902_);
  and (_00905_, _00904_, _00749_);
  and (_00906_, _00733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_00907_, _00906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_00908_, _00907_, _00722_);
  or (_00909_, _00908_, _00905_);
  and (_00910_, _00909_, _00758_);
  nor (_00911_, _00622_, _26521_);
  and (_00912_, _00911_, _00761_);
  or (_01286_, _00912_, _00910_);
  not (_00913_, _00781_);
  and (_00914_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_00915_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_00916_, _00915_, _00914_);
  and (_00917_, _00916_, _00758_);
  nand (_00918_, _00621_, _26512_);
  nand (_00919_, _00622_, _26521_);
  and (_00920_, _00919_, _00761_);
  and (_00921_, _00920_, _00918_);
  or (_01288_, _00921_, _00917_);
  nor (_00922_, _00781_, _00728_);
  and (_00923_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_00924_, _00923_, _00922_);
  and (_00925_, _00924_, _00758_);
  nand (_00926_, _00621_, _26505_);
  nand (_00927_, _00622_, _26512_);
  and (_00928_, _00927_, _00761_);
  and (_00929_, _00928_, _00926_);
  or (_01290_, _00929_, _00925_);
  nor (_00930_, _00781_, _00724_);
  and (_00931_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_00932_, _00931_, _00930_);
  and (_00933_, _00932_, _00758_);
  nand (_00934_, _00622_, _26505_);
  nand (_00935_, _00621_, _26497_);
  and (_00936_, _00935_, _00761_);
  and (_00937_, _00936_, _00934_);
  or (_01292_, _00937_, _00933_);
  and (_00938_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_00939_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or (_00940_, _00939_, _00938_);
  and (_00941_, _00940_, _00758_);
  nand (_00942_, _00621_, _26489_);
  nand (_00943_, _00622_, _26497_);
  and (_00944_, _00943_, _00761_);
  and (_00945_, _00944_, _00942_);
  or (_01294_, _00945_, _00941_);
  and (_00946_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_00947_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_00948_, _00947_, _00946_);
  and (_00949_, _00948_, _00758_);
  nand (_00950_, _00622_, _26489_);
  nand (_00951_, _00621_, _26482_);
  and (_00952_, _00951_, _00761_);
  and (_00953_, _00952_, _00950_);
  or (_01296_, _00953_, _00949_);
  and (_00954_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_00955_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_00956_, _00955_, _00954_);
  and (_00957_, _00956_, _00758_);
  nand (_00959_, _00621_, _26475_);
  nand (_00960_, _00622_, _26482_);
  and (_00961_, _00960_, _00761_);
  and (_00962_, _00961_, _00959_);
  or (_01297_, _00962_, _00957_);
  and (_00963_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_00964_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_00965_, _00964_, _00963_);
  and (_00966_, _00965_, _00758_);
  nand (_00967_, _00621_, _26543_);
  nand (_00968_, _00622_, _26475_);
  and (_00969_, _00968_, _00761_);
  and (_00970_, _00969_, _00967_);
  or (_01299_, _00970_, _00966_);
  and (_00971_, _00757_, _00622_);
  nand (_00972_, _00971_, _26543_);
  and (_00973_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_00974_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_00975_, _00974_, _00973_);
  or (_00976_, _00975_, _00757_);
  and (_00977_, _00976_, _27355_);
  and (_01301_, _00977_, _00972_);
  and (_00978_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_00979_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_00980_, _00979_, _00978_);
  and (_00981_, _00980_, _00758_);
  or (_00982_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_00983_, _00982_, _00622_);
  and (_00984_, _00983_, _00761_);
  or (_01303_, _00984_, _00981_);
  nand (_00986_, _00785_, _26521_);
  or (_00987_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_00988_, _00987_, _27355_);
  and (_01305_, _00988_, _00986_);
  or (_00989_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_00990_, _00989_, _27355_);
  nand (_00991_, _00785_, _26512_);
  and (_01307_, _00991_, _00990_);
  or (_00992_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_00993_, _00992_, _27355_);
  nand (_00994_, _00785_, _26505_);
  and (_01309_, _00994_, _00993_);
  or (_00995_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_00996_, _00995_, _27355_);
  nand (_00997_, _00785_, _26497_);
  and (_01310_, _00997_, _00996_);
  or (_00998_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_00999_, _00998_, _27355_);
  nand (_01000_, _00785_, _26489_);
  and (_01312_, _01000_, _00999_);
  or (_01002_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_01003_, _01002_, _27355_);
  nand (_01004_, _00785_, _26482_);
  and (_01314_, _01004_, _01003_);
  or (_01005_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_01006_, _01005_, _27355_);
  nand (_01007_, _00785_, _26475_);
  and (_01316_, _01007_, _01006_);
  nand (_01008_, _25514_, _25055_);
  or (_01009_, _25055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_01010_, _01009_, _00789_);
  and (_01011_, _01010_, _01008_);
  not (_01012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_01013_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01012_);
  or (_01014_, _01013_, _00621_);
  nor (_01015_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_01016_, _01015_, _01014_);
  nor (_01017_, _01016_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_01018_, _01017_, _00789_);
  or (_01019_, _01018_, _00792_);
  or (_01020_, _01019_, _01011_);
  nand (_01021_, _00792_, _26521_);
  and (_01022_, _01021_, _27355_);
  and (_01318_, _01022_, _01020_);
  or (_01023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_01024_, _01023_, _00789_);
  nand (_01025_, _27079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_01026_, _01025_, _00789_);
  or (_01027_, _01026_, _27080_);
  and (_01028_, _01027_, _01024_);
  or (_01029_, _01028_, _00792_);
  nand (_01030_, _00792_, _26512_);
  and (_01031_, _01030_, _27355_);
  and (_01320_, _01031_, _01029_);
  not (_01032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not (_01033_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_01034_, _00640_, _01033_);
  nor (_01035_, _01034_, _01032_);
  and (_01036_, _01034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_01037_, _01036_, _01035_);
  or (_01038_, _01037_, _00789_);
  or (_01039_, _25716_, _01032_);
  nand (_01040_, _01039_, _00789_);
  or (_01041_, _01040_, _25718_);
  and (_01042_, _01041_, _01038_);
  or (_01043_, _01042_, _00792_);
  nand (_01044_, _00792_, _26505_);
  and (_01045_, _01044_, _27355_);
  and (_01322_, _01045_, _01043_);
  and (_01046_, _00789_, _25778_);
  nand (_01047_, _01046_, _25514_);
  or (_01048_, _01046_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_01049_, _01048_, _00793_);
  and (_01050_, _01049_, _01047_);
  nor (_01051_, _00793_, _26497_);
  or (_01052_, _01051_, _01050_);
  and (_01323_, _01052_, _27355_);
  and (_01053_, _00789_, _25838_);
  nand (_01054_, _01053_, _25514_);
  or (_01055_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_01056_, _01055_, _00793_);
  and (_01057_, _01056_, _01054_);
  nor (_01058_, _00793_, _26489_);
  or (_01059_, _01058_, _01057_);
  and (_01325_, _01059_, _27355_);
  and (_01060_, _00789_, _25905_);
  nand (_01061_, _01060_, _25514_);
  or (_01062_, _01060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_01063_, _01062_, _01061_);
  or (_01064_, _01063_, _00792_);
  nand (_01065_, _00792_, _26482_);
  and (_01066_, _01065_, _27355_);
  and (_01327_, _01066_, _01064_);
  and (_01067_, _00789_, _25972_);
  nand (_01068_, _01067_, _25514_);
  or (_01069_, _01067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_01070_, _01069_, _00793_);
  and (_01071_, _01070_, _01068_);
  nor (_01072_, _00793_, _26475_);
  or (_01073_, _01072_, _01071_);
  and (_01329_, _01073_, _27355_);
  and (_01640_, t2_i, _27355_);
  nor (_01074_, t2_i, rst);
  and (_01643_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_01075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _27355_);
  nor (_01646_, _01075_, t2ex_i);
  and (_01649_, t2ex_i, _27355_);
  and (_01076_, _26457_, _26939_);
  and (_01077_, _01076_, _27666_);
  nand (_01078_, _01077_, _26543_);
  and (_01079_, _01076_, _27577_);
  not (_01080_, _01079_);
  and (_01081_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_01083_, _01082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_01084_, _01083_, _01081_);
  not (_01085_, _01084_);
  and (_01086_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01087_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_01088_, _01087_, _01086_);
  or (_01089_, _01077_, _01088_);
  and (_01090_, _01089_, _01080_);
  and (_01091_, _01090_, _01078_);
  and (_01092_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_01093_, _01092_, _01091_);
  and (_01652_, _01093_, _27355_);
  nand (_01094_, _01079_, _26543_);
  nor (_01095_, _01077_, _01085_);
  or (_01096_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_01097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_01098_, _01095_, _01097_);
  and (_01099_, _01098_, _01096_);
  or (_01100_, _01099_, _01079_);
  and (_01101_, _01100_, _27355_);
  and (_01655_, _01101_, _01094_);
  not (_01102_, _01082_);
  or (_01103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_01104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_01105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01104_);
  and (_01106_, _01105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_01107_, _01106_, _01103_);
  and (_01108_, _01076_, _25905_);
  and (_01109_, _01108_, _27576_);
  and (_01110_, _01076_, _27669_);
  nor (_01111_, _01110_, _01109_);
  and (_01112_, _01111_, _01107_);
  and (_01113_, _01112_, _01102_);
  and (_01114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_01115_, _01114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_01116_, _01115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_01117_, _01116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_01118_, _01117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_01119_, _01118_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_01120_, _01119_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01121_, _01120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_01122_, _01121_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_01123_, _01122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_01124_, _01123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_01125_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_01126_, _01125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_01127_, _01126_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_01128_, _01127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_01129_, _01128_);
  nand (_01130_, _01129_, _01113_);
  or (_01131_, _01113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_01132_, _01131_, _27355_);
  and (_01658_, _01132_, _01130_);
  nand (_01133_, _01110_, _26543_);
  not (_01134_, _01109_);
  not (_01135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_01136_, _01081_, _01135_);
  and (_01137_, _01136_, _01082_);
  and (_01138_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not (_01139_, _01137_);
  not (_01140_, _01083_);
  and (_01141_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01142_, _01128_, _01107_);
  and (_01143_, _01142_, _01141_);
  and (_01144_, _01119_, _01107_);
  or (_01145_, _01144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_01146_, _01144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01147_, _01146_, _01145_);
  or (_01148_, _01147_, _01143_);
  and (_01149_, _01148_, _01139_);
  or (_01150_, _01149_, _01138_);
  or (_01151_, _01150_, _01110_);
  and (_01152_, _01151_, _01134_);
  and (_01153_, _01152_, _01133_);
  and (_01154_, _01109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_01155_, _01154_, _01153_);
  and (_01661_, _01155_, _27355_);
  nand (_01156_, _01109_, _26543_);
  nor (_01157_, _01137_, _01097_);
  and (_01158_, _01139_, _01107_);
  and (_01159_, _01158_, _01127_);
  or (_01160_, _01159_, _01157_);
  nand (_01161_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_01162_, _01161_, _01142_);
  and (_01163_, _01162_, _01160_);
  nand (_01164_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_01165_, _01164_, _01111_);
  or (_01166_, _01165_, _01163_);
  nand (_01167_, _01110_, _01097_);
  and (_01168_, _01167_, _27355_);
  and (_01169_, _01168_, _01166_);
  and (_01664_, _01169_, _01156_);
  not (_01170_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor (_01171_, _01111_, _01170_);
  and (_01172_, _01158_, _01082_);
  and (_01173_, _01172_, _01111_);
  and (_01174_, _01173_, _01128_);
  or (_01175_, _01174_, _01171_);
  and (_01667_, _01175_, _27355_);
  or (_01176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_01177_, _00038_, _26923_);
  or (_01178_, _01177_, _01176_);
  nand (_01179_, _26926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_01180_, _01179_, _01177_);
  or (_01181_, _01180_, _26927_);
  and (_01182_, _01181_, _01178_);
  and (_01183_, _01076_, _00035_);
  or (_01184_, _01183_, _01182_);
  nand (_01185_, _01183_, _26543_);
  and (_01186_, _01185_, _27355_);
  and (_01670_, _01186_, _01184_);
  or (_01187_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not (_01188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_01189_, _01084_, _01188_);
  and (_01190_, _01189_, _01187_);
  or (_01191_, _01190_, _01077_);
  nand (_01192_, _01077_, _26521_);
  and (_01193_, _01192_, _01191_);
  or (_01194_, _01193_, _01079_);
  not (_01195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_01196_, _01079_, _01195_);
  and (_01197_, _01196_, _27355_);
  and (_02203_, _01197_, _01194_);
  nand (_01198_, _01077_, _26512_);
  and (_01199_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_01200_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_01201_, _01200_, _01199_);
  or (_01202_, _01201_, _01077_);
  and (_01203_, _01202_, _01080_);
  and (_01204_, _01203_, _01198_);
  and (_01205_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_01206_, _01205_, _01204_);
  and (_02205_, _01206_, _27355_);
  nand (_01207_, _01077_, _26505_);
  and (_01208_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_01209_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_01210_, _01209_, _01208_);
  or (_01211_, _01210_, _01077_);
  and (_01212_, _01211_, _01080_);
  and (_01213_, _01212_, _01207_);
  and (_01214_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_01215_, _01214_, _01213_);
  and (_02207_, _01215_, _27355_);
  nand (_01216_, _01077_, _26497_);
  and (_01217_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_01218_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_01219_, _01218_, _01217_);
  or (_01220_, _01219_, _01077_);
  and (_01221_, _01220_, _01080_);
  and (_01222_, _01221_, _01216_);
  and (_01223_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_01224_, _01223_, _01222_);
  and (_02209_, _01224_, _27355_);
  nand (_01225_, _01077_, _26489_);
  and (_01226_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_01227_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_01228_, _01227_, _01226_);
  or (_01229_, _01228_, _01077_);
  and (_01230_, _01229_, _01080_);
  and (_01231_, _01230_, _01225_);
  and (_01232_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_01233_, _01232_, _01231_);
  and (_02211_, _01233_, _27355_);
  nand (_01234_, _01077_, _26482_);
  and (_01235_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_01236_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_01237_, _01236_, _01235_);
  or (_01238_, _01237_, _01077_);
  and (_01240_, _01238_, _01080_);
  and (_01242_, _01240_, _01234_);
  and (_01244_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_01246_, _01244_, _01242_);
  and (_02213_, _01246_, _27355_);
  nand (_01249_, _01077_, _26475_);
  and (_01251_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_01253_, _01084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_01255_, _01253_, _01251_);
  or (_01257_, _01255_, _01077_);
  and (_01259_, _01257_, _01080_);
  and (_01261_, _01259_, _01249_);
  and (_01263_, _01079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_01265_, _01263_, _01261_);
  and (_02215_, _01265_, _27355_);
  and (_01268_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  not (_01270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_01272_, _01095_, _01270_);
  or (_01274_, _01272_, _01268_);
  or (_01276_, _01274_, _01079_);
  nand (_01278_, _01079_, _26521_);
  and (_01280_, _01278_, _27355_);
  and (_02217_, _01280_, _01276_);
  nand (_01283_, _01079_, _26512_);
  and (_01285_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  not (_01287_, _01095_);
  and (_01289_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_01291_, _01289_, _01285_);
  or (_01293_, _01291_, _01079_);
  and (_01295_, _01293_, _27355_);
  and (_02219_, _01295_, _01283_);
  nand (_01298_, _01079_, _26505_);
  and (_01300_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_01302_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_01304_, _01302_, _01300_);
  or (_01306_, _01304_, _01079_);
  and (_01308_, _01306_, _27355_);
  and (_02221_, _01308_, _01298_);
  nand (_01311_, _01079_, _26497_);
  and (_01313_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_01315_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_01317_, _01315_, _01313_);
  or (_01319_, _01317_, _01079_);
  and (_01321_, _01319_, _27355_);
  and (_02223_, _01321_, _01311_);
  nand (_01324_, _01079_, _26489_);
  and (_01326_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_01328_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_01330_, _01328_, _01326_);
  or (_01331_, _01330_, _01079_);
  and (_01332_, _01331_, _27355_);
  and (_02225_, _01332_, _01324_);
  nand (_01333_, _01079_, _26482_);
  and (_01334_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_01335_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_01336_, _01335_, _01334_);
  or (_01337_, _01336_, _01079_);
  and (_01338_, _01337_, _27355_);
  and (_02227_, _01338_, _01333_);
  nand (_01339_, _01079_, _26475_);
  and (_01340_, _01287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_01341_, _01095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_01342_, _01341_, _01340_);
  or (_01343_, _01342_, _01079_);
  and (_01344_, _01343_, _27355_);
  and (_02229_, _01344_, _01339_);
  and (_01345_, _01107_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_01346_, _01083_, _01195_);
  nand (_01347_, _01346_, _01128_);
  nand (_01348_, _01347_, _01345_);
  or (_01349_, _01107_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_01350_, _01349_, _01139_);
  and (_01351_, _01350_, _01348_);
  nand (_01352_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_01353_, _01352_, _01111_);
  or (_01354_, _01353_, _01351_);
  nand (_01355_, _01109_, _01188_);
  nand (_01356_, _01110_, _26521_);
  and (_01357_, _01356_, _27355_);
  and (_01358_, _01357_, _01355_);
  and (_02231_, _01358_, _01354_);
  and (_01359_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_01360_, _01359_, _01158_);
  and (_01361_, _01360_, _01128_);
  and (_01362_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_01363_, _01345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_01364_, _01114_, _01107_);
  nor (_01365_, _01364_, _01137_);
  and (_01366_, _01365_, _01363_);
  nor (_01367_, _01366_, _01362_);
  nand (_01368_, _01367_, _01111_);
  or (_01369_, _01368_, _01361_);
  nand (_01370_, _01110_, _26512_);
  or (_01371_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_01372_, _01371_, _27355_);
  and (_01373_, _01372_, _01370_);
  and (_02233_, _01373_, _01369_);
  and (_01374_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_01375_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_01376_, _01375_, _01142_);
  not (_01377_, _01364_);
  nor (_01378_, _01377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_01379_, _01377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_01380_, _01379_, _01378_);
  or (_01381_, _01380_, _01376_);
  and (_01382_, _01381_, _01139_);
  or (_01383_, _01382_, _01374_);
  or (_01384_, _01383_, _01110_);
  nand (_01385_, _01110_, _26505_);
  and (_01386_, _01385_, _01134_);
  and (_01387_, _01386_, _01384_);
  and (_01388_, _01109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_01389_, _01388_, _01387_);
  and (_02235_, _01389_, _27355_);
  not (_01390_, _01110_);
  nor (_01391_, _01390_, _26497_);
  and (_01392_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_01393_, _01392_, _01142_);
  nand (_01394_, _01115_, _01107_);
  and (_01395_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_01396_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_01397_, _01396_, _01137_);
  or (_01398_, _01397_, _01395_);
  or (_01399_, _01398_, _01393_);
  or (_01400_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_01401_, _01400_, _01111_);
  and (_01402_, _01401_, _01399_);
  and (_01403_, _01109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_01404_, _01403_, _01402_);
  or (_01405_, _01404_, _01391_);
  and (_02237_, _01405_, _27355_);
  and (_01406_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_01407_, _01406_, _01142_);
  nand (_01408_, _01116_, _01107_);
  and (_01409_, _01408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_01410_, _01408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_01411_, _01410_, _01137_);
  or (_01412_, _01411_, _01409_);
  or (_01413_, _01412_, _01407_);
  nor (_01414_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_01415_, _01414_, _01110_);
  and (_01416_, _01415_, _01413_);
  nor (_01417_, _01390_, _26489_);
  or (_01418_, _01417_, _01416_);
  or (_01419_, _01418_, _01109_);
  or (_01420_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_01421_, _01420_, _27355_);
  and (_02239_, _01421_, _01419_);
  and (_01422_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_01423_, _01422_, _01142_);
  nand (_01424_, _01117_, _01107_);
  and (_01425_, _01424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_01426_, _01424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_01427_, _01426_, _01137_);
  or (_01428_, _01427_, _01425_);
  or (_01429_, _01428_, _01423_);
  nor (_01430_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_01431_, _01430_, _01110_);
  and (_01432_, _01431_, _01429_);
  nor (_01433_, _01390_, _26482_);
  or (_01434_, _01433_, _01432_);
  or (_01435_, _01434_, _01109_);
  or (_01436_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_01437_, _01436_, _27355_);
  and (_02241_, _01437_, _01435_);
  nor (_01438_, _01390_, _26475_);
  and (_01439_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_01440_, _01439_, _01142_);
  and (_01441_, _01118_, _01107_);
  nor (_01442_, _01441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_01443_, _01442_, _01144_);
  or (_01444_, _01443_, _01137_);
  or (_01445_, _01444_, _01440_);
  nor (_01446_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_01447_, _01446_, _01110_);
  and (_01448_, _01447_, _01445_);
  or (_01449_, _01448_, _01109_);
  or (_01450_, _01449_, _01438_);
  or (_01451_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_01452_, _01451_, _27355_);
  and (_02243_, _01452_, _01450_);
  nor (_01453_, _01083_, _01270_);
  and (_01454_, _01453_, _01142_);
  and (_01455_, _01120_, _01107_);
  or (_01456_, _01455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_01457_, _01455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_01458_, _01457_, _01456_);
  or (_01459_, _01458_, _01137_);
  or (_01460_, _01459_, _01454_);
  and (_01461_, _01137_, _01270_);
  nor (_01462_, _01461_, _01110_);
  and (_01463_, _01462_, _01460_);
  and (_01464_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_01465_, _01464_, _01109_);
  or (_01466_, _01465_, _01463_);
  nand (_01467_, _01109_, _26521_);
  and (_01468_, _01467_, _27355_);
  and (_02245_, _01468_, _01466_);
  and (_01469_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_01470_, _01469_, _01142_);
  and (_01471_, _01121_, _01107_);
  or (_01472_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_01473_, _01471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_01474_, _01473_, _01472_);
  or (_01475_, _01474_, _01137_);
  or (_01476_, _01475_, _01470_);
  nor (_01477_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_01478_, _01477_, _01110_);
  and (_01479_, _01478_, _01476_);
  and (_01480_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_01481_, _01480_, _01109_);
  or (_01482_, _01481_, _01479_);
  nand (_01483_, _01109_, _26512_);
  and (_01484_, _01483_, _27355_);
  and (_02247_, _01484_, _01482_);
  and (_01485_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_01486_, _01485_, _01142_);
  nand (_01487_, _01122_, _01107_);
  and (_01488_, _01487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_01489_, _01487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_01490_, _01489_, _01137_);
  or (_01491_, _01490_, _01488_);
  or (_01492_, _01491_, _01486_);
  nor (_01493_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_01494_, _01493_, _01110_);
  and (_01495_, _01494_, _01492_);
  and (_01496_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_01497_, _01496_, _01109_);
  or (_01498_, _01497_, _01495_);
  nand (_01499_, _01109_, _26505_);
  and (_01500_, _01499_, _27355_);
  and (_02249_, _01500_, _01498_);
  and (_01501_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_01502_, _01501_, _01142_);
  nand (_01503_, _01123_, _01107_);
  and (_01504_, _01503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_01505_, _01503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_01506_, _01505_, _01137_);
  or (_01507_, _01506_, _01504_);
  or (_01508_, _01507_, _01502_);
  nor (_01509_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_01510_, _01509_, _01110_);
  and (_01511_, _01510_, _01508_);
  and (_01512_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_01513_, _01512_, _01109_);
  or (_01514_, _01513_, _01511_);
  nand (_01515_, _01109_, _26497_);
  and (_01516_, _01515_, _27355_);
  and (_02251_, _01516_, _01514_);
  nand (_01517_, _01109_, _26489_);
  and (_01518_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_01519_, _01518_, _01142_);
  nand (_01520_, _01124_, _01107_);
  and (_01521_, _01520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_01522_, _01520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_01523_, _01522_, _01137_);
  or (_01524_, _01523_, _01521_);
  or (_01525_, _01524_, _01519_);
  nor (_01526_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_01527_, _01526_, _01110_);
  and (_01528_, _01527_, _01525_);
  and (_01529_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_01530_, _01529_, _01109_);
  or (_01531_, _01530_, _01528_);
  and (_01532_, _01531_, _27355_);
  and (_02253_, _01532_, _01517_);
  and (_01533_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_01534_, _01533_, _01142_);
  nand (_01535_, _01125_, _01107_);
  and (_01536_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_01537_, _01535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_01538_, _01537_, _01137_);
  or (_01539_, _01538_, _01536_);
  or (_01540_, _01539_, _01534_);
  nor (_01541_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_01542_, _01541_, _01110_);
  and (_01543_, _01542_, _01540_);
  and (_01544_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_01545_, _01544_, _01109_);
  or (_01546_, _01545_, _01543_);
  nand (_01547_, _01109_, _26482_);
  and (_01548_, _01547_, _27355_);
  and (_02255_, _01548_, _01546_);
  and (_01549_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_01550_, _01549_, _01142_);
  nand (_01551_, _01126_, _01107_);
  and (_01552_, _01551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_01553_, _01551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_01554_, _01553_, _01137_);
  or (_01555_, _01554_, _01552_);
  or (_01556_, _01555_, _01550_);
  nor (_01557_, _01139_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_01558_, _01557_, _01110_);
  and (_01559_, _01558_, _01556_);
  and (_01560_, _01110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_01561_, _01560_, _01109_);
  or (_01562_, _01561_, _01559_);
  nand (_01563_, _01109_, _26475_);
  and (_01564_, _01563_, _27355_);
  and (_02257_, _01564_, _01562_);
  and (_01565_, _01177_, _25055_);
  nand (_01566_, _01565_, _25514_);
  not (_01567_, _01183_);
  or (_01568_, _01565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_01569_, _01568_, _01567_);
  and (_01570_, _01569_, _01566_);
  nor (_01571_, _01567_, _26521_);
  or (_01572_, _01571_, _01570_);
  and (_02259_, _01572_, _27355_);
  and (_01573_, _01177_, _26947_);
  nand (_01574_, _01573_, _25514_);
  or (_01575_, _01573_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_01576_, _01575_, _01574_);
  or (_01577_, _01576_, _01183_);
  nand (_01578_, _01183_, _26512_);
  and (_01579_, _01578_, _27355_);
  and (_02261_, _01579_, _01577_);
  nand (_01580_, _01177_, _27237_);
  and (_01581_, _01580_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_01582_, _01581_, _01183_);
  and (_01583_, _27240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_01584_, _01583_, _25718_);
  and (_01585_, _01584_, _01177_);
  or (_01586_, _01585_, _01582_);
  nand (_01587_, _01183_, _26505_);
  and (_01588_, _01587_, _27355_);
  and (_02263_, _01588_, _01586_);
  and (_01589_, _01177_, _25778_);
  or (_01590_, _01589_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_01591_, _01590_, _01567_);
  nand (_01592_, _01589_, _25514_);
  and (_01593_, _01592_, _01591_);
  nor (_01594_, _01567_, _26497_);
  or (_01595_, _01594_, _01593_);
  and (_02265_, _01595_, _27355_);
  and (_01596_, _01177_, _25838_);
  or (_01597_, _01596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_01598_, _01597_, _01567_);
  nand (_01599_, _01596_, _25514_);
  and (_01600_, _01599_, _01598_);
  nor (_01601_, _01567_, _26489_);
  or (_01602_, _01601_, _01600_);
  and (_02267_, _01602_, _27355_);
  and (_01603_, _01177_, _25905_);
  or (_01604_, _01603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_01605_, _01604_, _01567_);
  nand (_01606_, _01603_, _25514_);
  and (_01607_, _01606_, _01605_);
  nor (_01608_, _01567_, _26482_);
  or (_01609_, _01608_, _01607_);
  and (_02269_, _01609_, _27355_);
  and (_01610_, _01081_, _01170_);
  or (_01611_, _01610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_01612_, _01611_, _01177_);
  nand (_01613_, _27024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_01614_, _01613_, _01177_);
  or (_01615_, _01614_, _27025_);
  and (_01616_, _01615_, _01612_);
  or (_01617_, _01616_, _01183_);
  nand (_01618_, _01183_, _26475_);
  and (_01619_, _01618_, _27355_);
  and (_02271_, _01619_, _01617_);
  and (_01620_, _25101_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_01621_, _01620_, _25116_);
  nor (_01622_, _25053_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_01623_, _01622_, _01621_);
  nor (_01624_, _26436_, _26389_);
  and (_01625_, _01624_, _26454_);
  nand (_01626_, _26545_, _01625_);
  nor (_01627_, _26436_, _26390_);
  and (_01628_, _26938_, _26939_);
  and (_01629_, _01628_, _26940_);
  not (_01630_, _01629_);
  and (_01631_, _01630_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_01632_, _01631_, _26996_);
  and (_01633_, _01632_, _25116_);
  nor (_01634_, _01632_, _25116_);
  or (_01635_, _01634_, _01633_);
  not (_01636_, _01635_);
  not (_01637_, _25128_);
  and (_01638_, _01630_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_01639_, _01638_, _27006_);
  nor (_01641_, _01639_, _01637_);
  and (_01642_, _01639_, _01637_);
  nor (_01644_, _01642_, _01641_);
  and (_01645_, _26033_, _25053_);
  not (_01647_, _01645_);
  nor (_01648_, _26033_, _25053_);
  and (_01650_, _25073_, _25101_);
  and (_01651_, _01650_, _26938_);
  not (_01653_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_01654_, _25446_, _01653_);
  not (_01656_, _01654_);
  nor (_01657_, _01656_, _00755_);
  and (_01659_, _01657_, _01651_);
  not (_01660_, _01659_);
  and (_01662_, _25055_, _25116_);
  and (_01663_, _01651_, _01662_);
  not (_01665_, _01663_);
  and (_01666_, _01650_, _26457_);
  and (_01668_, _01666_, _01662_);
  not (_01669_, _01668_);
  and (_01671_, _01666_, _27035_);
  and (_01672_, _01666_, _27224_);
  nor (_01673_, _01672_, _01671_);
  and (_01674_, _01673_, _01669_);
  not (_01675_, _01666_);
  nor (_01676_, _01675_, _00755_);
  not (_01677_, _01676_);
  and (_01678_, _01651_, _27035_);
  and (_01679_, _01651_, _27224_);
  nor (_01680_, _01679_, _01678_);
  and (_01681_, _01680_, _01677_);
  and (_01682_, _01681_, _01674_);
  and (_01683_, _01682_, _01665_);
  or (_01684_, _01683_, _01656_);
  and (_01685_, _01684_, _01660_);
  nor (_01686_, _01685_, _01648_);
  and (_01687_, _01686_, _01647_);
  and (_01688_, _01687_, _01644_);
  and (_01689_, _01688_, _01636_);
  and (_01690_, _01689_, _26543_);
  not (_01691_, _01639_);
  and (_01692_, _01632_, _26034_);
  and (_01693_, _01692_, _01691_);
  and (_01694_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_01695_, _01632_, _26033_);
  and (_01696_, _01695_, _01639_);
  and (_01697_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_01698_, _01697_, _01694_);
  nor (_01699_, _01632_, _26034_);
  and (_01700_, _01699_, _01691_);
  and (_01701_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_01702_, _01632_, _26033_);
  and (_01703_, _01702_, _01639_);
  and (_01704_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_01705_, _01704_, _01701_);
  and (_01706_, _01705_, _01698_);
  not (_01707_, _01689_);
  and (_01708_, _01702_, _01691_);
  nand (_01709_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_01710_, _01692_, _01639_);
  nand (_01711_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_01712_, _01711_, _01709_);
  and (_01713_, _01695_, _01691_);
  nand (_01714_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_01715_, _01699_, _01639_);
  nand (_01716_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_01717_, _01716_, _01714_);
  and (_01718_, _01717_, _01712_);
  and (_01719_, _01718_, _01707_);
  and (_01720_, _01719_, _01706_);
  nor (_01721_, _01720_, _01690_);
  nand (_01722_, _01721_, _01627_);
  and (_01723_, _26454_, _26436_);
  not (_01724_, _01723_);
  nor (_01725_, _01724_, _26389_);
  not (_01726_, _25987_);
  and (_01727_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  nor (_01728_, _25996_, _26190_);
  nor (_01729_, _26018_, _26193_);
  nor (_01730_, _01729_, _01728_);
  and (_01731_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_01732_, _26002_, _26186_);
  nor (_01733_, _01732_, _01731_);
  and (_01734_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not (_01735_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_01736_, _26009_, _01735_);
  nor (_01737_, _01736_, _01734_);
  and (_01738_, _01737_, _01733_);
  and (_01739_, _01738_, _01730_);
  and (_01740_, _25993_, _25987_);
  not (_01741_, _01740_);
  nor (_01742_, _01741_, _01739_);
  nor (_01743_, _01742_, _01727_);
  not (_01744_, _01743_);
  nand (_01745_, _01744_, _01725_);
  and (_01746_, _01745_, _26454_);
  and (_01747_, _01746_, _01722_);
  and (_01748_, _01747_, _01626_);
  and (_01749_, _26286_, _26266_);
  or (_01750_, _01749_, _26337_);
  and (_01751_, _26359_, _26273_);
  and (_01752_, _26287_, _26269_);
  or (_01753_, _01752_, _26300_);
  or (_01754_, _01753_, _01751_);
  nor (_01755_, _01754_, _01750_);
  nor (_01756_, _26318_, _26275_);
  and (_01757_, _01756_, _26310_);
  and (_01758_, _01757_, _01755_);
  nor (_01759_, _01758_, _26393_);
  or (_01760_, _26316_, _26313_);
  and (_01761_, _26372_, _01760_);
  nor (_01762_, _01761_, _01759_);
  not (_01763_, _01762_);
  and (_01764_, _01763_, _01748_);
  not (_01765_, _01764_);
  and (_01766_, _01627_, _26454_);
  and (_01767_, _01689_, _26497_);
  and (_01768_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_01769_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_01770_, _01769_, _01768_);
  and (_01771_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_01772_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_01773_, _01772_, _01771_);
  and (_01774_, _01773_, _01770_);
  and (_01775_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_01776_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_01777_, _01776_, _01775_);
  and (_01778_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_01779_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_01780_, _01779_, _01778_);
  and (_01781_, _01780_, _01777_);
  and (_01782_, _01781_, _01707_);
  and (_01783_, _01782_, _01774_);
  nor (_01784_, _01783_, _01767_);
  and (_01785_, _01784_, _01766_);
  not (_01786_, _01785_);
  not (_01787_, _01625_);
  or (_01788_, _26571_, _01787_);
  not (_01789_, _01632_);
  and (_01790_, _01723_, _26389_);
  nand (_01791_, _01790_, _01789_);
  and (_01792_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_01793_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not (_01794_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_01795_, _26009_, _01794_);
  nor (_01796_, _01795_, _01793_);
  and (_01797_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_01798_, _26018_, _26057_);
  nor (_01799_, _01798_, _01797_);
  nor (_01800_, _25996_, _26051_);
  nor (_01801_, _26002_, _26043_);
  nor (_01802_, _01801_, _01800_);
  and (_01803_, _01802_, _01799_);
  and (_01804_, _01803_, _01796_);
  nor (_01805_, _01804_, _01741_);
  nor (_01806_, _01805_, _01792_);
  not (_01807_, _01806_);
  nand (_01808_, _01807_, _01725_);
  and (_01809_, _01808_, _01791_);
  and (_01810_, _01809_, _01788_);
  and (_01811_, _01810_, _01786_);
  or (_01812_, _01811_, _01765_);
  and (_01813_, _01689_, _26521_);
  and (_01814_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_01815_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_01816_, _01815_, _01814_);
  and (_01817_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_01818_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_01819_, _01818_, _01817_);
  and (_01820_, _01819_, _01816_);
  and (_01821_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_01822_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_01823_, _01822_, _01821_);
  and (_01824_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_01825_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_01826_, _01825_, _01824_);
  and (_01827_, _01826_, _01823_);
  and (_01828_, _01827_, _01707_);
  and (_01829_, _01828_, _01820_);
  nor (_01830_, _01829_, _01813_);
  and (_01831_, _01830_, _01766_);
  not (_01832_, _01831_);
  and (_01833_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  nor (_01834_, _25996_, _26008_);
  nor (_01835_, _26018_, _25994_);
  nor (_01836_, _01835_, _01834_);
  and (_01837_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_01838_, _26002_, _26015_);
  nor (_01839_, _01838_, _01837_);
  and (_01840_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not (_01841_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_01842_, _26009_, _01841_);
  nor (_01843_, _01842_, _01840_);
  and (_01844_, _01843_, _01839_);
  and (_01845_, _01844_, _01836_);
  nor (_01846_, _01845_, _01741_);
  nor (_01847_, _01846_, _01833_);
  not (_01848_, _01847_);
  and (_01849_, _01848_, _01725_);
  or (_01850_, _26553_, _01787_);
  nand (_01851_, _01790_, _26033_);
  nand (_01852_, _01851_, _01850_);
  nor (_01853_, _01852_, _01849_);
  and (_01854_, _01853_, _01832_);
  or (_01855_, _01854_, _01763_);
  nand (_01856_, _01855_, _01812_);
  and (_01857_, _01856_, _01623_);
  nor (_01858_, _01856_, _01623_);
  nor (_01859_, _01858_, _01857_);
  and (_01860_, _01620_, _01637_);
  nor (_01861_, _25042_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_01862_, _01861_, _01860_);
  and (_01863_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_01864_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_01865_, _01864_, _01863_);
  and (_01866_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_01867_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_01868_, _01867_, _01866_);
  and (_01869_, _01868_, _01865_);
  and (_01870_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_01871_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_01872_, _01871_, _01870_);
  and (_01873_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_01874_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_01875_, _01874_, _01873_);
  and (_01876_, _01875_, _01872_);
  and (_01877_, _01876_, _01707_);
  and (_01878_, _01877_, _01869_);
  and (_01879_, _01689_, _26489_);
  nor (_01880_, _01879_, _01878_);
  and (_01881_, _01880_, _01766_);
  not (_01882_, _01881_);
  not (_01883_, _26454_);
  and (_01884_, _01883_, _26436_);
  nor (_01885_, _26577_, _01787_);
  nor (_01886_, _01885_, _01884_);
  and (_01887_, _01790_, _01691_);
  and (_01888_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  nor (_01889_, _25996_, _26157_);
  nor (_01890_, _26018_, _26159_);
  nor (_01891_, _01890_, _01889_);
  not (_01892_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_01893_, _26009_, _01892_);
  nor (_01894_, _26002_, _26167_);
  nor (_01895_, _01894_, _01893_);
  and (_01896_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_01897_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_01898_, _01897_, _01896_);
  and (_01899_, _01898_, _01895_);
  and (_01900_, _01899_, _01891_);
  nor (_01901_, _01900_, _01741_);
  nor (_01902_, _01901_, _01888_);
  not (_01903_, _01902_);
  and (_01904_, _01903_, _01725_);
  nor (_01905_, _01904_, _01887_);
  and (_01906_, _01905_, _01886_);
  and (_01907_, _01906_, _01882_);
  or (_01908_, _01907_, _01765_);
  and (_01909_, _01689_, _26512_);
  and (_01910_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_01911_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_01912_, _01911_, _01910_);
  and (_01913_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_01914_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_01915_, _01914_, _01913_);
  and (_01916_, _01915_, _01912_);
  and (_01917_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_01918_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_01919_, _01918_, _01917_);
  and (_01920_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_01921_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_01922_, _01921_, _01920_);
  and (_01923_, _01922_, _01919_);
  and (_01924_, _01923_, _01707_);
  and (_01925_, _01924_, _01916_);
  nor (_01926_, _01925_, _01909_);
  and (_01927_, _01926_, _01766_);
  not (_01928_, _01927_);
  and (_01929_, _01627_, _01883_);
  nor (_01930_, _26559_, _01787_);
  nor (_01931_, _01930_, _01929_);
  and (_01932_, _01790_, _26153_);
  and (_01933_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_01934_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  not (_01935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_01936_, _26009_, _01935_);
  nor (_01937_, _01936_, _01934_);
  nor (_01938_, _25996_, _26127_);
  nor (_01939_, _26002_, _26132_);
  nor (_01940_, _01939_, _01938_);
  and (_01941_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_01942_, _26018_, _26129_);
  nor (_01943_, _01942_, _01941_);
  and (_01944_, _01943_, _01940_);
  and (_01945_, _01944_, _01937_);
  nor (_01946_, _01945_, _01741_);
  nor (_01947_, _01946_, _01933_);
  not (_01948_, _01947_);
  and (_01949_, _01948_, _01725_);
  nor (_01950_, _01949_, _01932_);
  and (_01951_, _01950_, _01931_);
  and (_01952_, _01951_, _01928_);
  or (_01953_, _01952_, _01763_);
  and (_01954_, _01953_, _01908_);
  and (_01955_, _01954_, _01862_);
  nor (_01956_, _01954_, _01862_);
  or (_01957_, _01956_, _01955_);
  and (_01958_, _01957_, _01859_);
  nor (_01959_, _01620_, _26922_);
  not (_01960_, _01959_);
  and (_01961_, _01884_, _26389_);
  nor (_01962_, _26583_, _01787_);
  nor (_01963_, _01962_, _01961_);
  and (_01964_, _01624_, _01883_);
  not (_01965_, _01964_);
  and (_01966_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  nor (_01967_, _25996_, _26218_);
  nor (_01968_, _26018_, _26212_);
  nor (_01969_, _01968_, _01967_);
  and (_01970_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  not (_01971_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_01972_, _26009_, _01971_);
  nor (_01973_, _01972_, _01970_);
  and (_01974_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_01975_, _26002_, _26222_);
  nor (_01976_, _01975_, _01974_);
  and (_01977_, _01976_, _01973_);
  and (_01978_, _01977_, _01969_);
  nor (_01979_, _01978_, _01741_);
  nor (_01980_, _01979_, _01966_);
  not (_01981_, _01980_);
  and (_01982_, _01981_, _01725_);
  and (_01983_, _01689_, _26482_);
  and (_01984_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_01985_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_01986_, _01985_, _01984_);
  and (_01987_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_01988_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_01989_, _01988_, _01987_);
  and (_01990_, _01989_, _01986_);
  and (_01991_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_01992_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_01993_, _01992_, _01991_);
  and (_01994_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_01995_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_01996_, _01995_, _01994_);
  and (_01997_, _01996_, _01993_);
  and (_01998_, _01997_, _01707_);
  and (_01999_, _01998_, _01990_);
  nor (_02000_, _01999_, _01983_);
  and (_02001_, _02000_, _01766_);
  nor (_02002_, _02001_, _01982_);
  and (_02003_, _02002_, _01965_);
  and (_02004_, _02003_, _01963_);
  and (_02005_, _02004_, _01765_);
  nor (_02006_, _02005_, _01960_);
  not (_02007_, _02006_);
  nor (_02008_, _01620_, _25073_);
  not (_02009_, _02008_);
  nor (_02010_, _26589_, _01787_);
  not (_02011_, _02010_);
  and (_02012_, _01689_, _26475_);
  and (_02013_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02014_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_02015_, _02014_, _02013_);
  and (_02016_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_02017_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_02018_, _02017_, _02016_);
  and (_02019_, _02018_, _02015_);
  and (_02020_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_02021_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_02022_, _02021_, _02020_);
  and (_02023_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_02024_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor (_02025_, _02024_, _02023_);
  and (_02026_, _02025_, _02022_);
  and (_02027_, _02026_, _01707_);
  and (_02028_, _02027_, _02019_);
  nor (_02029_, _02028_, _02012_);
  and (_02030_, _02029_, _01766_);
  not (_02031_, _02030_);
  and (_02032_, _26436_, _26390_);
  and (_02033_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_02034_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  not (_02035_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_02036_, _26009_, _02035_);
  nor (_02037_, _02036_, _02034_);
  nor (_02038_, _25996_, _26251_);
  nor (_02039_, _26002_, _26247_);
  nor (_02040_, _02039_, _02038_);
  and (_02041_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_02042_, _26018_, _26245_);
  nor (_02043_, _02042_, _02041_);
  and (_02044_, _02043_, _02040_);
  and (_02045_, _02044_, _02037_);
  nor (_02046_, _02045_, _01741_);
  nor (_02047_, _02046_, _02033_);
  not (_02048_, _02047_);
  and (_02049_, _02048_, _02032_);
  nor (_02050_, _01627_, _26454_);
  nor (_02051_, _02050_, _02049_);
  and (_02052_, _02051_, _02031_);
  and (_02053_, _02052_, _02011_);
  nor (_02054_, _02053_, _01764_);
  nor (_02055_, _02054_, _02009_);
  and (_02056_, _02054_, _02009_);
  nor (_02057_, _02056_, _02055_);
  and (_02058_, _02057_, _02007_);
  nor (_02059_, _01748_, _25101_);
  and (_02060_, _01748_, _25101_);
  nor (_02061_, _02060_, _02059_);
  not (_02062_, _02061_);
  nor (_02063_, _01620_, _25128_);
  not (_02064_, _02063_);
  nor (_02065_, _01907_, _01764_);
  and (_02066_, _02065_, _02064_);
  and (_02067_, _02005_, _01960_);
  nor (_02068_, _02067_, _02066_);
  and (_02069_, _02068_, _02062_);
  and (_02070_, _02069_, _02058_);
  and (_02071_, _02070_, _01958_);
  and (_02072_, _01620_, _26458_);
  nor (_02073_, _01620_, _25115_);
  nor (_02074_, _02073_, _02072_);
  and (_02075_, _02053_, _01764_);
  and (_02076_, _01811_, _01765_);
  nor (_02077_, _02076_, _02075_);
  and (_02078_, _02077_, _02074_);
  nor (_02079_, _02077_, _02074_);
  or (_02080_, _02079_, _02078_);
  not (_02081_, _02080_);
  and (_02082_, _01620_, _26922_);
  nor (_02083_, _25020_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_02084_, _02083_, _02082_);
  not (_02085_, _02084_);
  nor (_02086_, _02004_, _01765_);
  and (_02087_, _01715_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_02088_, _01710_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_02089_, _02088_, _02087_);
  and (_02090_, _01700_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_02091_, _01708_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_02092_, _02091_, _02090_);
  and (_02093_, _02092_, _02089_);
  and (_02094_, _01693_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_02095_, _01703_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_02096_, _02095_, _02094_);
  and (_02097_, _01713_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_02098_, _01696_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_02099_, _02098_, _02097_);
  and (_02100_, _02099_, _02096_);
  and (_02101_, _02100_, _01707_);
  and (_02102_, _02101_, _02093_);
  and (_02103_, _01689_, _26505_);
  nor (_02104_, _02103_, _02102_);
  and (_02105_, _02104_, _01766_);
  not (_02106_, _02105_);
  and (_02107_, _01790_, _26125_);
  not (_02108_, _26565_);
  and (_02109_, _02108_, _01625_);
  and (_02110_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_02111_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not (_02112_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_02113_, _26009_, _02112_);
  nor (_02114_, _02113_, _02111_);
  nor (_02115_, _26018_, _26111_);
  nor (_02116_, _26002_, _26097_);
  nor (_02117_, _02116_, _02115_);
  and (_02118_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_02119_, _25996_, _26105_);
  nor (_02120_, _02119_, _02118_);
  and (_02121_, _02120_, _02117_);
  and (_02122_, _02121_, _02114_);
  nor (_02123_, _02122_, _01741_);
  nor (_02124_, _02123_, _02110_);
  not (_02125_, _02124_);
  and (_02126_, _02125_, _01725_);
  or (_02127_, _02126_, _02109_);
  nor (_02128_, _02127_, _02107_);
  and (_02129_, _02128_, _02106_);
  nor (_02130_, _02129_, _01763_);
  nor (_02131_, _02130_, _02086_);
  nor (_02132_, _02131_, _02085_);
  and (_02133_, _02131_, _02085_);
  nor (_02134_, _02133_, _02132_);
  and (_02135_, _02134_, _02081_);
  nor (_02136_, _02065_, _02064_);
  and (_02137_, _25446_, _25099_);
  not (_02138_, _02137_);
  nor (_02139_, _02138_, _02136_);
  and (_02140_, _02139_, _02135_);
  and (_02141_, _02140_, _02071_);
  not (_02142_, _01748_);
  not (_02143_, _02005_);
  not (_02144_, _02131_);
  and (_02145_, _01855_, _01812_);
  and (_02146_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_02147_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_02148_, _02147_, _02146_);
  and (_02149_, _02148_, _01954_);
  not (_02150_, _01954_);
  and (_02151_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_02152_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_02153_, _02152_, _02151_);
  and (_02154_, _02153_, _02150_);
  or (_02155_, _02154_, _02149_);
  or (_02156_, _02155_, _02144_);
  not (_02157_, _02077_);
  and (_02158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and (_02159_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_02160_, _02159_, _02158_);
  and (_02161_, _02160_, _01954_);
  and (_02162_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_02163_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_02164_, _02163_, _02162_);
  and (_02165_, _02164_, _02150_);
  or (_02166_, _02165_, _02161_);
  or (_02167_, _02166_, _02131_);
  and (_02168_, _02167_, _02157_);
  and (_02169_, _02168_, _02156_);
  or (_02170_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_02171_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_02172_, _02171_, _02170_);
  and (_02173_, _02172_, _01954_);
  or (_02174_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_02175_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_02176_, _02175_, _02174_);
  and (_02177_, _02176_, _02150_);
  or (_02178_, _02177_, _02173_);
  or (_02179_, _02178_, _02144_);
  or (_02180_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_02181_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_02182_, _02181_, _02180_);
  and (_02183_, _02182_, _01954_);
  or (_02184_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_02185_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and (_02186_, _02185_, _02184_);
  and (_02187_, _02186_, _02150_);
  or (_02188_, _02187_, _02183_);
  or (_02189_, _02188_, _02131_);
  and (_02190_, _02189_, _02077_);
  and (_02191_, _02190_, _02179_);
  or (_02192_, _02191_, _02169_);
  and (_02193_, _02192_, _02065_);
  not (_02194_, _02065_);
  and (_02195_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_02196_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_02197_, _02196_, _02195_);
  and (_02198_, _02197_, _01954_);
  and (_02199_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_02200_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_02201_, _02200_, _02199_);
  and (_02202_, _02201_, _02150_);
  or (_02204_, _02202_, _02198_);
  or (_02206_, _02204_, _02144_);
  and (_02208_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_02210_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_02212_, _02210_, _02208_);
  and (_02214_, _02212_, _01954_);
  and (_02216_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_02218_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_02220_, _02218_, _02216_);
  and (_02222_, _02220_, _02150_);
  or (_02224_, _02222_, _02214_);
  or (_02226_, _02224_, _02131_);
  and (_02228_, _02226_, _02157_);
  and (_02230_, _02228_, _02206_);
  or (_02232_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_02234_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_02236_, _02234_, _02150_);
  and (_02238_, _02236_, _02232_);
  or (_02240_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_02242_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_02244_, _02242_, _01954_);
  and (_02246_, _02244_, _02240_);
  or (_02248_, _02246_, _02238_);
  or (_02250_, _02248_, _02144_);
  or (_02252_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_02254_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and (_02256_, _02254_, _02150_);
  and (_02258_, _02256_, _02252_);
  or (_02260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_02262_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and (_02264_, _02262_, _01954_);
  and (_02266_, _02264_, _02260_);
  or (_02268_, _02266_, _02258_);
  or (_02270_, _02268_, _02131_);
  and (_02272_, _02270_, _02077_);
  and (_02273_, _02272_, _02250_);
  or (_02274_, _02273_, _02230_);
  and (_02275_, _02274_, _02194_);
  or (_02276_, _02275_, _02193_);
  and (_02277_, _02276_, _02143_);
  and (_02278_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_02279_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_02280_, _02279_, _02278_);
  and (_02281_, _02280_, _01954_);
  and (_02282_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_02283_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_02284_, _02283_, _02282_);
  and (_02285_, _02284_, _02150_);
  or (_02286_, _02285_, _02281_);
  and (_02287_, _02286_, _02131_);
  and (_02288_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_02289_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_02290_, _02289_, _02288_);
  and (_02291_, _02290_, _01954_);
  and (_02292_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_02293_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_02294_, _02293_, _02292_);
  and (_02295_, _02294_, _02150_);
  or (_02296_, _02295_, _02291_);
  and (_02297_, _02296_, _02144_);
  or (_02298_, _02297_, _02287_);
  and (_02299_, _02298_, _02157_);
  or (_02300_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_02301_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_02302_, _02301_, _02150_);
  and (_02303_, _02302_, _02300_);
  or (_02304_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_02305_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_02306_, _02305_, _01954_);
  and (_02307_, _02306_, _02304_);
  or (_02308_, _02307_, _02303_);
  and (_02309_, _02308_, _02131_);
  or (_02310_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_02311_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_02312_, _02311_, _02150_);
  and (_02313_, _02312_, _02310_);
  or (_02314_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_02315_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_02316_, _02315_, _01954_);
  and (_02317_, _02316_, _02314_);
  or (_02318_, _02317_, _02313_);
  and (_02319_, _02318_, _02144_);
  or (_02320_, _02319_, _02309_);
  and (_02321_, _02320_, _02077_);
  or (_02322_, _02321_, _02299_);
  and (_02323_, _02322_, _02194_);
  and (_02324_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_02325_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_02326_, _02325_, _02324_);
  and (_02327_, _02326_, _01954_);
  and (_02328_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_02329_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_02330_, _02329_, _02328_);
  and (_02331_, _02330_, _02150_);
  or (_02332_, _02331_, _02327_);
  and (_02333_, _02332_, _02131_);
  and (_02334_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and (_02335_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_02336_, _02335_, _02334_);
  and (_02337_, _02336_, _01954_);
  and (_02338_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_02339_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_02340_, _02339_, _02338_);
  and (_02341_, _02340_, _02150_);
  or (_02342_, _02341_, _02337_);
  and (_02343_, _02342_, _02144_);
  or (_02344_, _02343_, _02333_);
  and (_02345_, _02344_, _02157_);
  or (_02346_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_02347_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_02348_, _02347_, _02346_);
  and (_02349_, _02348_, _01954_);
  or (_02350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_02351_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_02352_, _02351_, _02350_);
  and (_02353_, _02352_, _02150_);
  or (_02354_, _02353_, _02349_);
  and (_02355_, _02354_, _02131_);
  or (_02356_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_02357_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_02358_, _02357_, _02356_);
  and (_02359_, _02358_, _01954_);
  or (_02360_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_02361_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_02362_, _02361_, _02360_);
  and (_02363_, _02362_, _02150_);
  or (_02364_, _02363_, _02359_);
  and (_02365_, _02364_, _02144_);
  or (_02366_, _02365_, _02355_);
  and (_02367_, _02366_, _02077_);
  or (_02368_, _02367_, _02345_);
  and (_02369_, _02368_, _02065_);
  or (_02370_, _02369_, _02323_);
  and (_02371_, _02370_, _02005_);
  or (_02372_, _02371_, _02277_);
  or (_02373_, _02372_, _02054_);
  not (_02374_, _02054_);
  and (_02375_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and (_02376_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_02377_, _02376_, _02375_);
  and (_02378_, _02377_, _01954_);
  and (_02379_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_02380_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_02381_, _02380_, _02379_);
  and (_02382_, _02381_, _02150_);
  or (_02383_, _02382_, _02378_);
  or (_02384_, _02383_, _02144_);
  and (_02385_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and (_02386_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_02387_, _02386_, _02385_);
  and (_02388_, _02387_, _01954_);
  and (_02389_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_02390_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_02391_, _02390_, _02389_);
  and (_02392_, _02391_, _02150_);
  or (_02393_, _02392_, _02388_);
  or (_02394_, _02393_, _02131_);
  and (_02395_, _02394_, _02157_);
  and (_02396_, _02395_, _02384_);
  or (_02397_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_02398_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_02399_, _02398_, _02150_);
  and (_02400_, _02399_, _02397_);
  or (_02401_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_02402_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and (_02403_, _02402_, _01954_);
  and (_02404_, _02403_, _02401_);
  or (_02405_, _02404_, _02400_);
  or (_02406_, _02405_, _02144_);
  or (_02407_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_02408_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_02409_, _02408_, _02150_);
  and (_02410_, _02409_, _02407_);
  or (_02411_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_02412_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and (_02413_, _02412_, _01954_);
  and (_02414_, _02413_, _02411_);
  or (_02415_, _02414_, _02410_);
  or (_02416_, _02415_, _02131_);
  and (_02417_, _02416_, _02077_);
  and (_02418_, _02417_, _02406_);
  or (_02419_, _02418_, _02396_);
  and (_02420_, _02419_, _02194_);
  and (_02421_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_02422_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_02423_, _02422_, _02421_);
  and (_02424_, _02423_, _01954_);
  and (_02425_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_02426_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_02427_, _02426_, _02425_);
  and (_02428_, _02427_, _02150_);
  or (_02429_, _02428_, _02424_);
  or (_02430_, _02429_, _02144_);
  and (_02431_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_02432_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_02433_, _02432_, _02431_);
  and (_02434_, _02433_, _01954_);
  and (_02435_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_02436_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_02437_, _02436_, _02435_);
  and (_02438_, _02437_, _02150_);
  or (_02439_, _02438_, _02434_);
  or (_02440_, _02439_, _02131_);
  and (_02441_, _02440_, _02157_);
  and (_02442_, _02441_, _02430_);
  or (_02443_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_02444_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_02445_, _02444_, _02443_);
  and (_02446_, _02445_, _01954_);
  or (_02447_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_02448_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_02449_, _02448_, _02447_);
  and (_02450_, _02449_, _02150_);
  or (_02451_, _02450_, _02446_);
  or (_02452_, _02451_, _02144_);
  or (_02453_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_02454_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_02455_, _02454_, _02453_);
  and (_02456_, _02455_, _01954_);
  or (_02457_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_02458_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_02459_, _02458_, _02457_);
  and (_02460_, _02459_, _02150_);
  or (_02461_, _02460_, _02456_);
  or (_02462_, _02461_, _02131_);
  and (_02463_, _02462_, _02077_);
  and (_02464_, _02463_, _02452_);
  or (_02465_, _02464_, _02442_);
  and (_02466_, _02465_, _02065_);
  or (_02467_, _02466_, _02420_);
  and (_02468_, _02467_, _02143_);
  or (_02469_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_02470_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_02471_, _02470_, _02469_);
  and (_02472_, _02471_, _01954_);
  or (_02473_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_02474_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and (_02475_, _02474_, _02473_);
  and (_02476_, _02475_, _02150_);
  or (_02477_, _02476_, _02472_);
  and (_02478_, _02477_, _02144_);
  or (_02479_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_02480_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_02481_, _02480_, _02479_);
  and (_02482_, _02481_, _01954_);
  or (_02483_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_02484_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_02485_, _02484_, _02483_);
  and (_02486_, _02485_, _02150_);
  or (_02487_, _02486_, _02482_);
  and (_02488_, _02487_, _02131_);
  or (_02489_, _02488_, _02478_);
  and (_02490_, _02489_, _02077_);
  and (_02491_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_02492_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_02493_, _02492_, _02491_);
  and (_02494_, _02493_, _01954_);
  and (_02495_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_02496_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_02497_, _02496_, _02495_);
  and (_02498_, _02497_, _02150_);
  or (_02499_, _02498_, _02494_);
  and (_02500_, _02499_, _02144_);
  and (_02501_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and (_02502_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_02503_, _02502_, _02501_);
  and (_02504_, _02503_, _01954_);
  and (_02505_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and (_02506_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_02507_, _02506_, _02505_);
  and (_02508_, _02507_, _02150_);
  or (_02509_, _02508_, _02504_);
  and (_02510_, _02509_, _02131_);
  or (_02511_, _02510_, _02500_);
  and (_02512_, _02511_, _02157_);
  or (_02513_, _02512_, _02490_);
  and (_02514_, _02513_, _02065_);
  or (_02515_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_02516_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_02517_, _02516_, _02150_);
  and (_02518_, _02517_, _02515_);
  or (_02519_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_02520_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_02521_, _02520_, _01954_);
  and (_02522_, _02521_, _02519_);
  or (_02523_, _02522_, _02518_);
  and (_02524_, _02523_, _02144_);
  or (_02525_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_02526_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and (_02527_, _02526_, _02150_);
  and (_02528_, _02527_, _02525_);
  or (_02529_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_02530_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_02531_, _02530_, _01954_);
  and (_02532_, _02531_, _02529_);
  or (_02533_, _02532_, _02528_);
  and (_02534_, _02533_, _02131_);
  or (_02535_, _02534_, _02524_);
  and (_02536_, _02535_, _02077_);
  and (_02537_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and (_02538_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_02539_, _02538_, _02537_);
  and (_02540_, _02539_, _01954_);
  and (_02541_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_02542_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_02543_, _02542_, _02541_);
  and (_02544_, _02543_, _02150_);
  or (_02545_, _02544_, _02540_);
  and (_02546_, _02545_, _02144_);
  and (_02547_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_02548_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_02549_, _02548_, _02547_);
  and (_02550_, _02549_, _01954_);
  and (_02551_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_02552_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_02553_, _02552_, _02551_);
  and (_02554_, _02553_, _02150_);
  or (_02555_, _02554_, _02550_);
  and (_02556_, _02555_, _02131_);
  or (_02557_, _02556_, _02546_);
  and (_02558_, _02557_, _02157_);
  or (_02559_, _02558_, _02536_);
  and (_02560_, _02559_, _02194_);
  or (_02561_, _02560_, _02514_);
  and (_02562_, _02561_, _02005_);
  or (_02563_, _02562_, _02468_);
  or (_02564_, _02563_, _02374_);
  and (_02565_, _02564_, _02373_);
  or (_02566_, _02565_, _02142_);
  and (_02567_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and (_02568_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_02569_, _02568_, _02567_);
  and (_02570_, _02569_, _01954_);
  and (_02571_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and (_02572_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_02573_, _02572_, _02571_);
  and (_02574_, _02573_, _02150_);
  or (_02575_, _02574_, _02570_);
  and (_02576_, _02575_, _02131_);
  and (_02577_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and (_02578_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_02579_, _02578_, _02577_);
  and (_02580_, _02579_, _01954_);
  and (_02581_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and (_02582_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_02583_, _02582_, _02581_);
  and (_02584_, _02583_, _02150_);
  or (_02585_, _02584_, _02580_);
  and (_02586_, _02585_, _02144_);
  or (_02587_, _02586_, _02576_);
  and (_02588_, _02587_, _02157_);
  or (_02589_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_02590_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_02591_, _02590_, _02150_);
  and (_02592_, _02591_, _02589_);
  or (_02593_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_02594_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and (_02595_, _02594_, _01954_);
  and (_02596_, _02595_, _02593_);
  or (_02597_, _02596_, _02592_);
  and (_02598_, _02597_, _02131_);
  or (_02599_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_02600_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and (_02601_, _02600_, _02150_);
  and (_02602_, _02601_, _02599_);
  or (_02603_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_02604_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and (_02605_, _02604_, _01954_);
  and (_02606_, _02605_, _02603_);
  or (_02607_, _02606_, _02602_);
  and (_02608_, _02607_, _02144_);
  or (_02609_, _02608_, _02598_);
  and (_02610_, _02609_, _02077_);
  or (_02611_, _02610_, _02588_);
  and (_02612_, _02611_, _02194_);
  and (_02613_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_02614_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_02615_, _02614_, _02613_);
  and (_02616_, _02615_, _01954_);
  and (_02617_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_02618_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_02619_, _02618_, _02617_);
  and (_02620_, _02619_, _02150_);
  or (_02621_, _02620_, _02616_);
  and (_02622_, _02621_, _02131_);
  and (_02623_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_02624_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_02625_, _02624_, _02623_);
  and (_02626_, _02625_, _01954_);
  and (_02627_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_02628_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_02629_, _02628_, _02627_);
  and (_02630_, _02629_, _02150_);
  or (_02631_, _02630_, _02626_);
  and (_02632_, _02631_, _02144_);
  or (_02633_, _02632_, _02622_);
  and (_02634_, _02633_, _02157_);
  or (_02635_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_02636_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_02637_, _02636_, _02635_);
  and (_02638_, _02637_, _01954_);
  or (_02639_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_02640_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_02641_, _02640_, _02639_);
  and (_02642_, _02641_, _02150_);
  or (_02643_, _02642_, _02638_);
  and (_02644_, _02643_, _02131_);
  or (_02645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_02646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_02647_, _02646_, _02645_);
  and (_02648_, _02647_, _01954_);
  or (_02649_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_02650_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_02651_, _02650_, _02649_);
  and (_02652_, _02651_, _02150_);
  or (_02653_, _02652_, _02648_);
  and (_02654_, _02653_, _02144_);
  or (_02655_, _02654_, _02644_);
  and (_02656_, _02655_, _02077_);
  or (_02657_, _02656_, _02634_);
  and (_02658_, _02657_, _02065_);
  or (_02659_, _02658_, _02612_);
  and (_02660_, _02659_, _02005_);
  and (_02661_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_02662_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_02663_, _02662_, _02661_);
  and (_02664_, _02663_, _01954_);
  and (_02665_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_02666_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_02667_, _02666_, _02665_);
  and (_02668_, _02667_, _02150_);
  or (_02669_, _02668_, _02664_);
  or (_02670_, _02669_, _02144_);
  and (_02671_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_02672_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_02673_, _02672_, _02671_);
  and (_02674_, _02673_, _01954_);
  and (_02675_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_02676_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_02677_, _02676_, _02675_);
  and (_02678_, _02677_, _02150_);
  or (_02679_, _02678_, _02674_);
  or (_02680_, _02679_, _02131_);
  and (_02681_, _02680_, _02157_);
  and (_02682_, _02681_, _02670_);
  or (_02683_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_02684_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_02685_, _02684_, _02683_);
  and (_02686_, _02685_, _01954_);
  or (_02687_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_02688_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_02689_, _02688_, _02687_);
  and (_02690_, _02689_, _02150_);
  or (_02691_, _02690_, _02686_);
  or (_02692_, _02691_, _02144_);
  or (_02693_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_02694_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_02695_, _02694_, _02693_);
  and (_02696_, _02695_, _01954_);
  or (_02697_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_02698_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_02699_, _02698_, _02697_);
  and (_02700_, _02699_, _02150_);
  or (_02701_, _02700_, _02696_);
  or (_02702_, _02701_, _02131_);
  and (_02703_, _02702_, _02077_);
  and (_02704_, _02703_, _02692_);
  or (_02705_, _02704_, _02682_);
  and (_02707_, _02705_, _02065_);
  and (_02708_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_02709_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_02710_, _02709_, _02708_);
  and (_02711_, _02710_, _01954_);
  and (_02712_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_02713_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_02714_, _02713_, _02712_);
  and (_02716_, _02714_, _02150_);
  or (_02717_, _02716_, _02711_);
  or (_02718_, _02717_, _02144_);
  and (_02719_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_02720_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_02721_, _02720_, _02719_);
  and (_02722_, _02721_, _01954_);
  and (_02723_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_02724_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_02725_, _02724_, _02723_);
  and (_02726_, _02725_, _02150_);
  or (_02727_, _02726_, _02722_);
  or (_02728_, _02727_, _02131_);
  and (_02729_, _02728_, _02157_);
  and (_02730_, _02729_, _02718_);
  or (_02731_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_02732_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_02733_, _02732_, _02150_);
  and (_02734_, _02733_, _02731_);
  or (_02735_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_02736_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_02737_, _02736_, _01954_);
  and (_02738_, _02737_, _02735_);
  or (_02739_, _02738_, _02734_);
  or (_02740_, _02739_, _02144_);
  or (_02741_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_02742_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_02743_, _02742_, _02150_);
  and (_02744_, _02743_, _02741_);
  or (_02745_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_02746_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_02747_, _02746_, _01954_);
  and (_02748_, _02747_, _02745_);
  or (_02749_, _02748_, _02744_);
  or (_02750_, _02749_, _02131_);
  and (_02751_, _02750_, _02077_);
  and (_02752_, _02751_, _02740_);
  or (_02753_, _02752_, _02730_);
  and (_02754_, _02753_, _02194_);
  or (_02755_, _02754_, _02707_);
  and (_02756_, _02755_, _02143_);
  or (_02757_, _02756_, _02660_);
  or (_02758_, _02757_, _02054_);
  and (_02759_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_02760_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_02761_, _02760_, _02759_);
  and (_02762_, _02761_, _02150_);
  and (_02763_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_02764_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_02765_, _02764_, _02763_);
  and (_02766_, _02765_, _01954_);
  or (_02767_, _02766_, _02762_);
  or (_02768_, _02767_, _02144_);
  and (_02769_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_02770_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_02771_, _02770_, _02769_);
  and (_02772_, _02771_, _02150_);
  and (_02773_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_02774_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_02775_, _02774_, _02773_);
  and (_02776_, _02775_, _01954_);
  or (_02777_, _02776_, _02772_);
  or (_02778_, _02777_, _02131_);
  and (_02779_, _02778_, _02157_);
  and (_02780_, _02779_, _02768_);
  or (_02781_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_02782_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_02783_, _02782_, _01954_);
  and (_02785_, _02783_, _02781_);
  or (_02786_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_02787_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_02788_, _02787_, _02150_);
  and (_02789_, _02788_, _02786_);
  or (_02790_, _02789_, _02785_);
  or (_02791_, _02790_, _02144_);
  or (_02792_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_02793_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_02794_, _02793_, _01954_);
  and (_02795_, _02794_, _02792_);
  or (_02796_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_02797_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_02798_, _02797_, _02150_);
  and (_02799_, _02798_, _02796_);
  or (_02800_, _02799_, _02795_);
  or (_02801_, _02800_, _02131_);
  and (_02802_, _02801_, _02077_);
  and (_02803_, _02802_, _02791_);
  or (_02804_, _02803_, _02780_);
  and (_02805_, _02804_, _02194_);
  and (_02806_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_02807_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_02808_, _02807_, _01954_);
  or (_02809_, _02808_, _02806_);
  and (_02810_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_02811_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_02812_, _02811_, _02150_);
  or (_02813_, _02812_, _02810_);
  and (_02814_, _02813_, _02809_);
  or (_02815_, _02814_, _02144_);
  and (_02816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_02817_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_02818_, _02817_, _01954_);
  or (_02819_, _02818_, _02816_);
  and (_02820_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_02821_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_02822_, _02821_, _02150_);
  or (_02823_, _02822_, _02820_);
  and (_02824_, _02823_, _02819_);
  or (_02825_, _02824_, _02131_);
  and (_02826_, _02825_, _02157_);
  and (_02827_, _02826_, _02815_);
  or (_02828_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_02829_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_02830_, _02829_, _02828_);
  or (_02831_, _02830_, _02150_);
  or (_02832_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_02833_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_02834_, _02833_, _02832_);
  or (_02835_, _02834_, _01954_);
  and (_02836_, _02835_, _02831_);
  or (_02837_, _02836_, _02144_);
  or (_02838_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_02839_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_02840_, _02839_, _02838_);
  or (_02841_, _02840_, _02150_);
  or (_02842_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_02843_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_02844_, _02843_, _02842_);
  or (_02845_, _02844_, _01954_);
  and (_02846_, _02845_, _02841_);
  or (_02847_, _02846_, _02131_);
  and (_02848_, _02847_, _02077_);
  and (_02849_, _02848_, _02837_);
  or (_02850_, _02849_, _02827_);
  and (_02851_, _02850_, _02065_);
  or (_02852_, _02851_, _02805_);
  and (_02853_, _02852_, _02143_);
  and (_02854_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_02855_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_02856_, _02855_, _02854_);
  and (_02857_, _02856_, _01954_);
  and (_02858_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_02859_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_02860_, _02859_, _02858_);
  and (_02861_, _02860_, _02150_);
  or (_02862_, _02861_, _02857_);
  and (_02863_, _02862_, _02131_);
  and (_02864_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_02865_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_02866_, _02865_, _02864_);
  and (_02867_, _02866_, _01954_);
  and (_02868_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_02869_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_02870_, _02869_, _02868_);
  and (_02871_, _02870_, _02150_);
  or (_02872_, _02871_, _02867_);
  and (_02873_, _02872_, _02144_);
  or (_02874_, _02873_, _02863_);
  and (_02875_, _02874_, _02157_);
  or (_02876_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_02877_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_02878_, _02877_, _02876_);
  and (_02879_, _02878_, _01954_);
  or (_02880_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_02881_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_02882_, _02881_, _02880_);
  and (_02883_, _02882_, _02150_);
  or (_02884_, _02883_, _02879_);
  and (_02885_, _02884_, _02131_);
  or (_02886_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_02887_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_02888_, _02887_, _02886_);
  and (_02889_, _02888_, _01954_);
  or (_02890_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_02891_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_02892_, _02891_, _02890_);
  and (_02893_, _02892_, _02150_);
  or (_02894_, _02893_, _02889_);
  and (_02895_, _02894_, _02144_);
  or (_02896_, _02895_, _02885_);
  and (_02897_, _02896_, _02077_);
  or (_02898_, _02897_, _02875_);
  and (_02899_, _02898_, _02065_);
  and (_02900_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and (_02901_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or (_02902_, _02901_, _02900_);
  and (_02903_, _02902_, _01954_);
  and (_02904_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  and (_02905_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or (_02906_, _02905_, _02904_);
  and (_02907_, _02906_, _02150_);
  or (_02908_, _02907_, _02903_);
  and (_02909_, _02908_, _02131_);
  and (_02910_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  and (_02911_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or (_02912_, _02911_, _02910_);
  and (_02913_, _02912_, _01954_);
  and (_02914_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and (_02915_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or (_02916_, _02915_, _02914_);
  and (_02917_, _02916_, _02150_);
  or (_02918_, _02917_, _02913_);
  and (_02919_, _02918_, _02144_);
  or (_02920_, _02919_, _02909_);
  and (_02921_, _02920_, _02157_);
  or (_02922_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_02923_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  and (_02924_, _02923_, _02922_);
  and (_02925_, _02924_, _01954_);
  or (_02926_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or (_02927_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and (_02928_, _02927_, _02926_);
  and (_02929_, _02928_, _02150_);
  or (_02930_, _02929_, _02925_);
  and (_02931_, _02930_, _02131_);
  or (_02932_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or (_02933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  and (_02934_, _02933_, _02932_);
  and (_02935_, _02934_, _01954_);
  or (_02936_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or (_02937_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and (_02938_, _02937_, _02936_);
  and (_02939_, _02938_, _02150_);
  or (_02940_, _02939_, _02935_);
  and (_02941_, _02940_, _02144_);
  or (_02942_, _02941_, _02931_);
  and (_02943_, _02942_, _02077_);
  or (_02944_, _02943_, _02921_);
  and (_02945_, _02944_, _02194_);
  or (_02946_, _02945_, _02899_);
  and (_02947_, _02946_, _02005_);
  or (_02948_, _02947_, _02853_);
  or (_02949_, _02948_, _02374_);
  and (_02950_, _02949_, _02758_);
  or (_02951_, _02950_, _01748_);
  and (_02952_, _02951_, _02566_);
  or (_02953_, _02952_, _02141_);
  not (_02954_, _02141_);
  or (_02955_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_02956_, _02955_, _27355_);
  and (_02715_, _02956_, _02953_);
  nor (_02957_, _02138_, _01623_);
  nor (_02958_, _02138_, _01862_);
  nor (_02959_, _02958_, _02957_);
  nor (_02960_, _02138_, _02084_);
  nor (_02961_, _02138_, _02074_);
  nor (_02962_, _02961_, _02960_);
  and (_02963_, _02962_, _02959_);
  and (_02964_, _02137_, _02063_);
  nor (_02965_, _02138_, _01959_);
  nor (_02966_, _02965_, _02964_);
  nor (_02967_, _01650_, _01620_);
  and (_02968_, _02967_, _02137_);
  not (_02969_, _02968_);
  and (_02970_, _02969_, _02966_);
  and (_02971_, _02970_, _02137_);
  and (_02972_, _02971_, _02963_);
  not (_02973_, _02972_);
  and (_02974_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_02975_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25182_);
  and (_02976_, _02975_, _25168_);
  and (_02977_, _02976_, _25574_);
  nor (_02978_, _26521_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not (_02979_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_02980_, _02976_, _02979_);
  and (_02981_, _02980_, _24073_);
  or (_02982_, _02981_, _02978_);
  or (_02983_, _02982_, _02977_);
  and (_02985_, _02983_, _02972_);
  or (_03577_, _02985_, _02974_);
  and (_02986_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nand (_02987_, _02975_, _25172_);
  nor (_02988_, _02987_, _25514_);
  nor (_02989_, _26512_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_02990_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_02991_, _02975_, _25177_);
  or (_02992_, _02991_, _02990_);
  and (_02993_, _02975_, _25174_);
  or (_02994_, _02993_, _02992_);
  and (_02995_, _02994_, _24023_);
  or (_02996_, _02995_, _02989_);
  or (_02997_, _02996_, _02988_);
  and (_02998_, _02997_, _02972_);
  or (_03581_, _02998_, _02986_);
  and (_02999_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_03000_, _02975_, _25175_);
  nor (_03001_, _03000_, _25514_);
  nor (_03002_, _26505_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_03003_, _25175_, _25182_);
  and (_03004_, _24059_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_03005_, _03004_, _03003_);
  or (_03006_, _03005_, _03002_);
  or (_03007_, _03006_, _03001_);
  and (_03008_, _03007_, _02972_);
  or (_03587_, _03008_, _02999_);
  and (_03009_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_03010_, _02991_, _25574_);
  nor (_03011_, _26497_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_03012_, _25177_, _25182_);
  and (_03013_, _24009_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_03014_, _03013_, _03012_);
  or (_03015_, _03014_, _03011_);
  or (_03016_, _03015_, _03010_);
  and (_03017_, _03016_, _02972_);
  or (_03591_, _03017_, _03009_);
  and (_03018_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_03019_, _02990_, _25168_);
  nor (_03020_, _03019_, _25514_);
  nor (_03021_, _26489_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_03022_, _25168_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_03023_, _23958_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_03024_, _03023_, _03022_);
  or (_03025_, _03024_, _03021_);
  or (_03026_, _03025_, _03020_);
  and (_03027_, _03026_, _02972_);
  or (_03595_, _03027_, _03018_);
  and (_03028_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_03029_, _02990_, _25172_);
  nor (_03030_, _03029_, _25514_);
  nor (_03031_, _26482_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_03032_, _25172_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_03033_, _23995_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_03034_, _03033_, _03032_);
  or (_03035_, _03034_, _03031_);
  or (_03036_, _03035_, _03030_);
  and (_03037_, _03036_, _02972_);
  or (_03600_, _03037_, _03028_);
  and (_03038_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand (_03040_, _02990_, _25175_);
  nor (_03041_, _03040_, _25514_);
  nor (_03042_, _26475_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_03043_, _25175_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_03044_, _24040_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_03045_, _03044_, _03043_);
  or (_03046_, _03045_, _03042_);
  or (_03047_, _03046_, _03041_);
  and (_03048_, _03047_, _02972_);
  or (_03605_, _03048_, _03038_);
  and (_03050_, _02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_03051_, _02990_, _25177_);
  not (_03052_, _03051_);
  nor (_03053_, _03052_, _25514_);
  nand (_03054_, _26543_, _02979_);
  or (_03055_, _23978_, _02979_);
  and (_03056_, _03055_, _03052_);
  and (_03057_, _03056_, _03054_);
  or (_03058_, _03057_, _03053_);
  and (_03059_, _03058_, _02972_);
  or (_03607_, _03059_, _03050_);
  and (_03060_, _02983_, _02137_);
  and (_03061_, _02957_, _01862_);
  and (_03062_, _03061_, _02962_);
  and (_03063_, _03062_, _02970_);
  and (_03064_, _03063_, _03060_);
  not (_03065_, _03063_);
  and (_03066_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_03613_, _03066_, _03064_);
  and (_03067_, _02997_, _02137_);
  and (_03069_, _03063_, _03067_);
  and (_03070_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_03616_, _03070_, _03069_);
  and (_03071_, _03007_, _02137_);
  and (_03072_, _03063_, _03071_);
  and (_03073_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_03619_, _03073_, _03072_);
  and (_03074_, _03016_, _02137_);
  and (_03075_, _03063_, _03074_);
  and (_03076_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_03622_, _03076_, _03075_);
  and (_03077_, _03026_, _02137_);
  and (_03078_, _03063_, _03077_);
  and (_03079_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_03626_, _03079_, _03078_);
  and (_03080_, _03036_, _02137_);
  and (_03081_, _03063_, _03080_);
  and (_03082_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_03629_, _03082_, _03081_);
  and (_03083_, _03047_, _02137_);
  and (_03085_, _03063_, _03083_);
  and (_03086_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_03632_, _03086_, _03085_);
  and (_03087_, _03058_, _02137_);
  and (_03088_, _03063_, _03087_);
  and (_03089_, _03065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_03634_, _03089_, _03088_);
  and (_03090_, _02958_, _01623_);
  and (_03091_, _03090_, _02962_);
  and (_03092_, _03091_, _02970_);
  and (_03093_, _03092_, _03060_);
  not (_03094_, _03092_);
  and (_03095_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_03641_, _03095_, _03093_);
  and (_03096_, _03092_, _03067_);
  and (_03097_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_03644_, _03097_, _03096_);
  and (_03098_, _03092_, _03071_);
  and (_03099_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_03647_, _03099_, _03098_);
  and (_03101_, _03092_, _03074_);
  and (_03102_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_03650_, _03102_, _03101_);
  and (_03103_, _03092_, _03077_);
  and (_03104_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_03653_, _03104_, _03103_);
  and (_03105_, _03092_, _03080_);
  and (_03106_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_03656_, _03106_, _03105_);
  and (_03107_, _03092_, _03083_);
  and (_03109_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_03659_, _03109_, _03107_);
  and (_03110_, _03092_, _03087_);
  and (_03111_, _03094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_03662_, _03111_, _03110_);
  and (_03112_, _02958_, _02957_);
  and (_03113_, _03112_, _02962_);
  and (_03114_, _03113_, _02970_);
  and (_03115_, _03114_, _03060_);
  not (_03116_, _03114_);
  and (_03118_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_03667_, _03118_, _03115_);
  and (_03119_, _03114_, _03067_);
  and (_03120_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_03670_, _03120_, _03119_);
  and (_03121_, _03114_, _03071_);
  and (_03122_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_03673_, _03122_, _03121_);
  and (_03123_, _03114_, _03074_);
  and (_03124_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_03676_, _03124_, _03123_);
  and (_03126_, _03114_, _03077_);
  and (_03127_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_03679_, _03127_, _03126_);
  and (_03128_, _03114_, _03080_);
  and (_03129_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_03682_, _03129_, _03128_);
  and (_03130_, _03114_, _03083_);
  and (_03131_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_03685_, _03131_, _03130_);
  and (_03133_, _03114_, _03087_);
  and (_03134_, _03116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_03688_, _03134_, _03133_);
  and (_03135_, _02960_, _02074_);
  and (_03136_, _03135_, _02959_);
  and (_03137_, _03136_, _02970_);
  and (_03138_, _03137_, _03060_);
  not (_03139_, _03137_);
  and (_03140_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_03694_, _03140_, _03138_);
  and (_03142_, _03137_, _03067_);
  and (_03143_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_03697_, _03143_, _03142_);
  and (_03144_, _03137_, _03071_);
  and (_03145_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_03700_, _03145_, _03144_);
  and (_03146_, _03137_, _03074_);
  and (_03147_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_03704_, _03147_, _03146_);
  and (_03148_, _03137_, _03077_);
  and (_03150_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_03707_, _03150_, _03148_);
  and (_03151_, _03137_, _03080_);
  and (_03152_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_03710_, _03152_, _03151_);
  and (_03153_, _03137_, _03083_);
  and (_03154_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_03713_, _03154_, _03153_);
  and (_03155_, _03137_, _03087_);
  and (_03156_, _03139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_03716_, _03156_, _03155_);
  and (_03159_, _03135_, _03061_);
  and (_03160_, _03159_, _02970_);
  and (_03161_, _03160_, _03060_);
  not (_03162_, _03160_);
  and (_03163_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_03720_, _03163_, _03161_);
  and (_03164_, _03160_, _03067_);
  and (_03165_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_03723_, _03165_, _03164_);
  and (_03167_, _03160_, _03071_);
  and (_03168_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_03726_, _03168_, _03167_);
  and (_03169_, _03160_, _03074_);
  and (_03170_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_03729_, _03170_, _03169_);
  and (_03171_, _03160_, _03077_);
  and (_03172_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_03733_, _03172_, _03171_);
  and (_03173_, _03160_, _03080_);
  and (_03174_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_03736_, _03174_, _03173_);
  and (_03175_, _03160_, _03083_);
  and (_03176_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_03739_, _03176_, _03175_);
  and (_03177_, _03160_, _03087_);
  and (_03178_, _03162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_03741_, _03178_, _03177_);
  and (_03179_, _03135_, _03090_);
  and (_03180_, _03179_, _02970_);
  and (_03181_, _03180_, _03060_);
  not (_03182_, _03180_);
  and (_03183_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_03745_, _03183_, _03181_);
  and (_03184_, _03180_, _03067_);
  and (_03185_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_03748_, _03185_, _03184_);
  and (_03186_, _03180_, _03071_);
  and (_03187_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_03751_, _03187_, _03186_);
  and (_03188_, _03180_, _03074_);
  and (_03189_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_03754_, _03189_, _03188_);
  and (_03190_, _03180_, _03077_);
  and (_03191_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_03758_, _03191_, _03190_);
  and (_03192_, _03180_, _03080_);
  and (_03193_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_03761_, _03193_, _03192_);
  and (_03194_, _03180_, _03083_);
  and (_03195_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_03764_, _03195_, _03194_);
  and (_03196_, _03180_, _03087_);
  and (_03197_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_03766_, _03197_, _03196_);
  and (_03198_, _03135_, _03112_);
  and (_03199_, _03198_, _02970_);
  and (_03200_, _03199_, _03060_);
  not (_03201_, _03199_);
  and (_03202_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_03771_, _03202_, _03200_);
  and (_03203_, _03199_, _03067_);
  and (_03204_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_03774_, _03204_, _03203_);
  and (_03205_, _03199_, _03071_);
  and (_03206_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_03777_, _03206_, _03205_);
  and (_03207_, _03199_, _03074_);
  and (_03208_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_03780_, _03208_, _03207_);
  and (_03209_, _03199_, _03077_);
  and (_03210_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_03784_, _03210_, _03209_);
  and (_03211_, _03199_, _03080_);
  and (_03212_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_03787_, _03212_, _03211_);
  and (_03213_, _03199_, _03083_);
  and (_03214_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_03790_, _03214_, _03213_);
  and (_03215_, _03199_, _03087_);
  and (_03216_, _03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_03793_, _03216_, _03215_);
  and (_03217_, _02961_, _02084_);
  and (_03218_, _03217_, _02959_);
  and (_03219_, _03218_, _02970_);
  and (_03220_, _03219_, _03060_);
  not (_03221_, _03219_);
  and (_03222_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_03799_, _03222_, _03220_);
  and (_03223_, _03219_, _03067_);
  and (_03224_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_03802_, _03224_, _03223_);
  and (_03225_, _03219_, _03071_);
  and (_03226_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_03805_, _03226_, _03225_);
  and (_03227_, _03219_, _03074_);
  and (_03228_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_03808_, _03228_, _03227_);
  and (_03229_, _03219_, _03077_);
  and (_03230_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_03812_, _03230_, _03229_);
  and (_03231_, _03219_, _03080_);
  and (_03232_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_03815_, _03232_, _03231_);
  and (_03233_, _03219_, _03083_);
  and (_03234_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_03818_, _03234_, _03233_);
  and (_03235_, _03219_, _03087_);
  and (_03236_, _03221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_03820_, _03236_, _03235_);
  and (_03237_, _03217_, _03061_);
  and (_03238_, _03237_, _02970_);
  and (_03239_, _03238_, _03060_);
  not (_03240_, _03238_);
  and (_03241_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_03824_, _03241_, _03239_);
  and (_03242_, _03238_, _03067_);
  and (_03243_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_03827_, _03243_, _03242_);
  and (_03244_, _03238_, _03071_);
  and (_03245_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_03830_, _03245_, _03244_);
  and (_03246_, _03238_, _03074_);
  and (_03247_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_03833_, _03247_, _03246_);
  and (_03248_, _03238_, _03077_);
  and (_03249_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_03837_, _03249_, _03248_);
  and (_03250_, _03238_, _03080_);
  and (_03251_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_03840_, _03251_, _03250_);
  and (_03252_, _03238_, _03083_);
  and (_03253_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_03843_, _03253_, _03252_);
  and (_03254_, _03238_, _03087_);
  and (_03255_, _03240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_03845_, _03255_, _03254_);
  and (_03256_, _03217_, _03090_);
  and (_03257_, _03256_, _02970_);
  and (_03258_, _03257_, _03060_);
  not (_03259_, _03257_);
  and (_03260_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_03850_, _03260_, _03258_);
  and (_03261_, _03257_, _03067_);
  and (_03262_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_03853_, _03262_, _03261_);
  and (_03263_, _03257_, _03071_);
  and (_03264_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_03856_, _03264_, _03263_);
  and (_03265_, _03257_, _03074_);
  and (_03266_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_03859_, _03266_, _03265_);
  and (_03267_, _03257_, _03077_);
  and (_03268_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_03862_, _03268_, _03267_);
  and (_03269_, _03257_, _03080_);
  and (_03270_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_03865_, _03270_, _03269_);
  and (_03271_, _03257_, _03083_);
  and (_03272_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_03868_, _03272_, _03271_);
  and (_03273_, _03257_, _03087_);
  and (_03274_, _03259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_03871_, _03274_, _03273_);
  and (_03275_, _03217_, _03112_);
  and (_03276_, _03275_, _02970_);
  and (_03277_, _03276_, _03060_);
  not (_03278_, _03276_);
  and (_03279_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_03875_, _03279_, _03277_);
  and (_03280_, _03276_, _03067_);
  and (_03281_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_03878_, _03281_, _03280_);
  and (_03282_, _03276_, _03071_);
  and (_03283_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_03881_, _03283_, _03282_);
  and (_03284_, _03276_, _03074_);
  and (_03285_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_03884_, _03285_, _03284_);
  and (_03286_, _03276_, _03077_);
  and (_03287_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_03887_, _03287_, _03286_);
  and (_03288_, _03276_, _03080_);
  and (_03289_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_03891_, _03289_, _03288_);
  and (_03290_, _03276_, _03083_);
  and (_03291_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_03894_, _03291_, _03290_);
  and (_03292_, _03276_, _03087_);
  and (_03293_, _03278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_03896_, _03293_, _03292_);
  and (_03294_, _02961_, _02960_);
  and (_03295_, _03294_, _02959_);
  and (_03296_, _03295_, _02970_);
  and (_03297_, _03296_, _03060_);
  not (_03298_, _03296_);
  and (_03299_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_03901_, _03299_, _03297_);
  and (_03300_, _03296_, _03067_);
  and (_03301_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_03904_, _03301_, _03300_);
  and (_03303_, _03296_, _03071_);
  and (_03304_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_03907_, _03304_, _03303_);
  and (_03305_, _03296_, _03074_);
  and (_03306_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_03910_, _03306_, _03305_);
  and (_03307_, _03296_, _03077_);
  and (_03308_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_03913_, _03308_, _03307_);
  and (_03309_, _03296_, _03080_);
  and (_03310_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_03917_, _03310_, _03309_);
  and (_03311_, _03296_, _03083_);
  and (_03312_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_03920_, _03312_, _03311_);
  and (_03313_, _03296_, _03087_);
  and (_03314_, _03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_03922_, _03314_, _03313_);
  and (_03315_, _03294_, _03061_);
  and (_03316_, _03315_, _02970_);
  and (_03317_, _03316_, _03060_);
  not (_03318_, _03316_);
  and (_03319_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_03926_, _03319_, _03317_);
  and (_03320_, _03316_, _03067_);
  and (_03321_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_03929_, _03321_, _03320_);
  and (_03322_, _03316_, _03071_);
  and (_03323_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_03932_, _03323_, _03322_);
  and (_03324_, _03316_, _03074_);
  and (_03325_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_03935_, _03325_, _03324_);
  and (_03326_, _03316_, _03077_);
  and (_03327_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_03938_, _03327_, _03326_);
  and (_03328_, _03316_, _03080_);
  and (_03329_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_03942_, _03329_, _03328_);
  and (_03330_, _03316_, _03083_);
  and (_03331_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_03945_, _03331_, _03330_);
  and (_03332_, _03316_, _03087_);
  and (_03333_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_03947_, _03333_, _03332_);
  and (_03334_, _03294_, _03090_);
  and (_03335_, _03334_, _02970_);
  and (_03336_, _03335_, _03060_);
  not (_03337_, _03335_);
  and (_03338_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_03952_, _03338_, _03336_);
  and (_03339_, _03335_, _03067_);
  and (_03340_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_03955_, _03340_, _03339_);
  and (_03341_, _03335_, _03071_);
  and (_03342_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_03958_, _03342_, _03341_);
  and (_03343_, _03335_, _03074_);
  and (_03344_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_03961_, _03344_, _03343_);
  and (_03345_, _03335_, _03077_);
  and (_03346_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_03964_, _03346_, _03345_);
  and (_03347_, _03335_, _03080_);
  and (_03348_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_03967_, _03348_, _03347_);
  and (_03349_, _03335_, _03083_);
  and (_03350_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_03970_, _03350_, _03349_);
  and (_03351_, _03335_, _03087_);
  and (_03352_, _03337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_03973_, _03352_, _03351_);
  and (_03353_, _03294_, _03112_);
  and (_03354_, _03353_, _02970_);
  and (_03355_, _03354_, _03060_);
  not (_03356_, _03354_);
  and (_03357_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_03977_, _03357_, _03355_);
  and (_03358_, _03354_, _03067_);
  and (_03359_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_03980_, _03359_, _03358_);
  and (_03360_, _03354_, _03071_);
  and (_03361_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_03983_, _03361_, _03360_);
  and (_03362_, _03354_, _03074_);
  and (_03363_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_03987_, _03363_, _03362_);
  and (_03364_, _03354_, _03077_);
  and (_03365_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_03990_, _03365_, _03364_);
  and (_03366_, _03354_, _03080_);
  and (_03367_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_03993_, _03367_, _03366_);
  and (_03368_, _03354_, _03083_);
  and (_03369_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_03997_, _03369_, _03368_);
  and (_03370_, _03354_, _03087_);
  and (_03371_, _03356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_03999_, _03371_, _03370_);
  not (_03372_, _02967_);
  and (_03373_, _02964_, _25085_);
  and (_03374_, _03373_, _03372_);
  and (_03375_, _03374_, _02963_);
  and (_03376_, _03375_, _03060_);
  not (_03377_, _03375_);
  and (_03378_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or (_04005_, _03378_, _03376_);
  and (_03379_, _03375_, _03067_);
  and (_03380_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or (_04008_, _03380_, _03379_);
  and (_03381_, _03375_, _03071_);
  and (_03382_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or (_04011_, _03382_, _03381_);
  and (_03383_, _03375_, _03074_);
  and (_03384_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or (_04014_, _03384_, _03383_);
  and (_03385_, _03375_, _03077_);
  and (_03386_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or (_04017_, _03386_, _03385_);
  and (_03387_, _03375_, _03080_);
  and (_03388_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or (_04021_, _03388_, _03387_);
  and (_03389_, _03375_, _03083_);
  and (_03390_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or (_04024_, _03390_, _03389_);
  and (_03391_, _03375_, _03087_);
  and (_03392_, _03377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or (_04026_, _03392_, _03391_);
  and (_03393_, _03374_, _03062_);
  and (_03394_, _03393_, _03060_);
  not (_03395_, _03393_);
  and (_03396_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_04030_, _03396_, _03394_);
  and (_03397_, _03393_, _03067_);
  and (_03398_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_04033_, _03398_, _03397_);
  and (_03399_, _03393_, _03071_);
  and (_03400_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_04036_, _03400_, _03399_);
  and (_03401_, _03393_, _03074_);
  and (_03402_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_04039_, _03402_, _03401_);
  and (_03403_, _03393_, _03077_);
  and (_03404_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_04042_, _03404_, _03403_);
  and (_03405_, _03393_, _03080_);
  and (_03406_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_04045_, _03406_, _03405_);
  and (_03407_, _03393_, _03083_);
  and (_03408_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_04049_, _03408_, _03407_);
  and (_03409_, _03393_, _03087_);
  and (_03410_, _03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_04051_, _03410_, _03409_);
  and (_03411_, _03374_, _03091_);
  and (_03412_, _03411_, _03060_);
  not (_03413_, _03411_);
  and (_03414_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_04055_, _03414_, _03412_);
  and (_03415_, _03411_, _03067_);
  and (_03416_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_04058_, _03416_, _03415_);
  and (_03417_, _03411_, _03071_);
  and (_03418_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_04061_, _03418_, _03417_);
  and (_03419_, _03411_, _03074_);
  and (_03420_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_04064_, _03420_, _03419_);
  and (_03421_, _03411_, _03077_);
  and (_03422_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_04067_, _03422_, _03421_);
  and (_03423_, _03411_, _03080_);
  and (_03424_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_04070_, _03424_, _03423_);
  and (_03425_, _03411_, _03083_);
  and (_03426_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_04073_, _03426_, _03425_);
  and (_03427_, _03411_, _03087_);
  and (_03428_, _03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_04076_, _03428_, _03427_);
  and (_03429_, _03374_, _03113_);
  and (_03430_, _03429_, _03060_);
  not (_03431_, _03429_);
  and (_03432_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or (_04079_, _03432_, _03430_);
  and (_03433_, _03429_, _03067_);
  and (_03434_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or (_04082_, _03434_, _03433_);
  and (_03435_, _03429_, _03071_);
  and (_03436_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or (_04085_, _03436_, _03435_);
  and (_03437_, _03429_, _03074_);
  and (_03438_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or (_04088_, _03438_, _03437_);
  and (_03439_, _03429_, _03077_);
  and (_03440_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or (_04091_, _03440_, _03439_);
  and (_03441_, _03429_, _03080_);
  and (_03442_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or (_04094_, _03442_, _03441_);
  and (_03444_, _03429_, _03083_);
  and (_03445_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or (_04097_, _03445_, _03444_);
  and (_03446_, _03429_, _03087_);
  and (_03447_, _03431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or (_04100_, _03447_, _03446_);
  and (_03448_, _03374_, _03136_);
  and (_03449_, _03448_, _03060_);
  not (_03450_, _03448_);
  and (_03451_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or (_04104_, _03451_, _03449_);
  and (_03452_, _03448_, _03067_);
  and (_03453_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or (_04107_, _03453_, _03452_);
  and (_03454_, _03448_, _03071_);
  and (_03455_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or (_04110_, _03455_, _03454_);
  and (_03456_, _03448_, _03074_);
  and (_03457_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or (_04113_, _03457_, _03456_);
  and (_03458_, _03448_, _03077_);
  and (_03459_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or (_04116_, _03459_, _03458_);
  and (_03460_, _03448_, _03080_);
  and (_03461_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or (_04119_, _03461_, _03460_);
  and (_03462_, _03448_, _03083_);
  and (_03463_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or (_04122_, _03463_, _03462_);
  and (_03464_, _03448_, _03087_);
  and (_03465_, _03450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_04124_, _03465_, _03464_);
  and (_03466_, _03374_, _03159_);
  and (_03467_, _03466_, _03060_);
  not (_03468_, _03466_);
  and (_03469_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_04129_, _03469_, _03467_);
  and (_03470_, _03466_, _03067_);
  and (_03471_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_04132_, _03471_, _03470_);
  and (_03472_, _03466_, _03071_);
  and (_03473_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_04135_, _03473_, _03472_);
  and (_03474_, _03466_, _03074_);
  and (_03475_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_04138_, _03475_, _03474_);
  and (_03476_, _03466_, _03077_);
  and (_03477_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_04141_, _03477_, _03476_);
  and (_03478_, _03466_, _03080_);
  and (_03479_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_04144_, _03479_, _03478_);
  and (_03480_, _03466_, _03083_);
  and (_03481_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_04147_, _03481_, _03480_);
  and (_03482_, _03466_, _03087_);
  and (_03483_, _03468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_04150_, _03483_, _03482_);
  and (_03484_, _03374_, _03179_);
  and (_03485_, _03484_, _03060_);
  not (_03486_, _03484_);
  and (_03487_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_04153_, _03487_, _03485_);
  and (_03488_, _03484_, _03067_);
  and (_03489_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_04157_, _03489_, _03488_);
  and (_03490_, _03484_, _03071_);
  and (_03491_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_04160_, _03491_, _03490_);
  and (_03492_, _03484_, _03074_);
  and (_03493_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_04163_, _03493_, _03492_);
  and (_03494_, _03484_, _03077_);
  and (_03495_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_04166_, _03495_, _03494_);
  and (_03496_, _03484_, _03080_);
  and (_03497_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_04169_, _03497_, _03496_);
  and (_03498_, _03484_, _03083_);
  and (_03499_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_04172_, _03499_, _03498_);
  and (_03500_, _03484_, _03087_);
  and (_03501_, _03486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_04174_, _03501_, _03500_);
  and (_03502_, _03374_, _03198_);
  and (_03503_, _03502_, _03060_);
  not (_03504_, _03502_);
  and (_03505_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or (_04178_, _03505_, _03503_);
  and (_03506_, _03502_, _03067_);
  and (_03507_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or (_04181_, _03507_, _03506_);
  and (_03508_, _03502_, _03071_);
  and (_03509_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or (_04185_, _03509_, _03508_);
  and (_03510_, _03502_, _03074_);
  and (_03511_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or (_04188_, _03511_, _03510_);
  and (_03512_, _03502_, _03077_);
  and (_03513_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or (_04192_, _03513_, _03512_);
  and (_03514_, _03502_, _03080_);
  and (_03515_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or (_04195_, _03515_, _03514_);
  and (_03516_, _03502_, _03083_);
  and (_03517_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or (_04198_, _03517_, _03516_);
  and (_03518_, _03502_, _03087_);
  and (_03519_, _03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or (_04200_, _03519_, _03518_);
  and (_03520_, _03374_, _03218_);
  and (_03521_, _03520_, _03060_);
  not (_03522_, _03520_);
  and (_03523_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_04204_, _03523_, _03521_);
  and (_03524_, _03520_, _03067_);
  and (_03525_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_04207_, _03525_, _03524_);
  and (_03526_, _03520_, _03071_);
  and (_03527_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_04210_, _03527_, _03526_);
  and (_03528_, _03520_, _03074_);
  and (_03529_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_04213_, _03529_, _03528_);
  and (_03530_, _03520_, _03077_);
  and (_03531_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_04216_, _03531_, _03530_);
  and (_03532_, _03520_, _03080_);
  and (_03533_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_04219_, _03533_, _03532_);
  and (_03534_, _03520_, _03083_);
  and (_03535_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_04222_, _03535_, _03534_);
  and (_03536_, _03520_, _03087_);
  and (_03537_, _03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_04225_, _03537_, _03536_);
  and (_03538_, _03374_, _03237_);
  and (_03539_, _03538_, _03060_);
  not (_03540_, _03538_);
  and (_03541_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or (_04228_, _03541_, _03539_);
  and (_03542_, _03538_, _03067_);
  and (_03543_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or (_04231_, _03543_, _03542_);
  and (_03544_, _03538_, _03071_);
  and (_03545_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or (_04234_, _03545_, _03544_);
  and (_03546_, _03538_, _03074_);
  and (_03547_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or (_04238_, _03547_, _03546_);
  and (_03548_, _03538_, _03077_);
  and (_03549_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or (_04241_, _03549_, _03548_);
  and (_03550_, _03538_, _03080_);
  and (_03551_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or (_04244_, _03551_, _03550_);
  and (_03552_, _03538_, _03083_);
  and (_03553_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or (_04247_, _03553_, _03552_);
  and (_03554_, _03538_, _03087_);
  and (_03555_, _03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or (_04249_, _03555_, _03554_);
  and (_03556_, _03374_, _03256_);
  and (_03557_, _03556_, _03060_);
  not (_03558_, _03556_);
  and (_03559_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or (_04253_, _03559_, _03557_);
  and (_03560_, _03556_, _03067_);
  and (_03561_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or (_04256_, _03561_, _03560_);
  and (_03562_, _03556_, _03071_);
  and (_03563_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or (_04259_, _03563_, _03562_);
  and (_03564_, _03556_, _03074_);
  and (_03565_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or (_04262_, _03565_, _03564_);
  and (_03566_, _03556_, _03077_);
  and (_03567_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or (_04266_, _03567_, _03566_);
  and (_03568_, _03556_, _03080_);
  and (_03569_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or (_04269_, _03569_, _03568_);
  and (_03570_, _03556_, _03083_);
  and (_03571_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or (_04272_, _03571_, _03570_);
  and (_03572_, _03556_, _03087_);
  and (_03573_, _03558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or (_04274_, _03573_, _03572_);
  and (_03574_, _03374_, _03275_);
  and (_03575_, _03574_, _03060_);
  not (_03576_, _03574_);
  and (_03578_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_04278_, _03578_, _03575_);
  and (_03579_, _03574_, _03067_);
  and (_03580_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_04281_, _03580_, _03579_);
  and (_03582_, _03574_, _03071_);
  and (_03583_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_04284_, _03583_, _03582_);
  and (_03585_, _03574_, _03074_);
  and (_03586_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_04287_, _03586_, _03585_);
  and (_03588_, _03574_, _03077_);
  and (_03589_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_04290_, _03589_, _03588_);
  and (_03590_, _03574_, _03080_);
  and (_03592_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_04294_, _03592_, _03590_);
  and (_03593_, _03574_, _03083_);
  and (_03594_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_04297_, _03594_, _03593_);
  and (_03596_, _03574_, _03087_);
  and (_03597_, _03576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_04300_, _03597_, _03596_);
  and (_03598_, _03374_, _03295_);
  and (_03599_, _03598_, _03060_);
  not (_03601_, _03598_);
  and (_03602_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_04303_, _03602_, _03599_);
  and (_03603_, _03598_, _03067_);
  and (_03604_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_04306_, _03604_, _03603_);
  and (_03606_, _03598_, _03071_);
  and (_03608_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_04309_, _03608_, _03606_);
  and (_03609_, _03598_, _03074_);
  and (_03610_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_04312_, _03610_, _03609_);
  and (_03611_, _03598_, _03077_);
  and (_03612_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_04315_, _03612_, _03611_);
  and (_03614_, _03598_, _03080_);
  and (_03615_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_04319_, _03615_, _03614_);
  and (_03617_, _03598_, _03083_);
  and (_03618_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_04322_, _03618_, _03617_);
  and (_03620_, _03598_, _03087_);
  and (_03621_, _03601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_04324_, _03621_, _03620_);
  and (_03623_, _03374_, _03315_);
  and (_03624_, _03623_, _03060_);
  not (_03625_, _03623_);
  and (_03627_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or (_04328_, _03627_, _03624_);
  and (_03628_, _03623_, _03067_);
  and (_03630_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or (_04331_, _03630_, _03628_);
  and (_03631_, _03623_, _03071_);
  and (_03633_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or (_04334_, _03633_, _03631_);
  and (_03635_, _03623_, _03074_);
  and (_03636_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or (_04337_, _03636_, _03635_);
  and (_03637_, _03623_, _03077_);
  and (_03638_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or (_04340_, _03638_, _03637_);
  and (_03639_, _03623_, _03080_);
  and (_03640_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or (_04343_, _03640_, _03639_);
  and (_03642_, _03623_, _03083_);
  and (_03643_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or (_04347_, _03643_, _03642_);
  and (_03645_, _03623_, _03087_);
  and (_03646_, _03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or (_04349_, _03646_, _03645_);
  and (_03648_, _03374_, _03334_);
  and (_03649_, _03648_, _03060_);
  not (_03651_, _03648_);
  and (_03652_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or (_04353_, _03652_, _03649_);
  and (_03654_, _03648_, _03067_);
  and (_03655_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or (_04356_, _03655_, _03654_);
  and (_03657_, _03648_, _03071_);
  and (_03658_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or (_04359_, _03658_, _03657_);
  and (_03660_, _03648_, _03074_);
  and (_03661_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or (_04362_, _03661_, _03660_);
  and (_03663_, _03648_, _03077_);
  and (_03664_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or (_04365_, _03664_, _03663_);
  and (_03665_, _03648_, _03080_);
  and (_03666_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or (_04368_, _03666_, _03665_);
  and (_03668_, _03648_, _03083_);
  and (_03669_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or (_04371_, _03669_, _03668_);
  and (_03671_, _03648_, _03087_);
  and (_03672_, _03651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or (_04374_, _03672_, _03671_);
  and (_03674_, _03374_, _03353_);
  and (_03675_, _03674_, _03060_);
  not (_03677_, _03674_);
  and (_03678_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_04377_, _03678_, _03675_);
  and (_03680_, _03674_, _03067_);
  and (_03681_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_04380_, _03681_, _03680_);
  and (_03683_, _03674_, _03071_);
  and (_03684_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_04383_, _03684_, _03683_);
  and (_03686_, _03674_, _03074_);
  and (_03687_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_04386_, _03687_, _03686_);
  and (_03689_, _03674_, _03077_);
  and (_03690_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_04389_, _03690_, _03689_);
  and (_03691_, _03674_, _03080_);
  and (_03692_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_04392_, _03692_, _03691_);
  and (_03693_, _03674_, _03083_);
  and (_03695_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_04395_, _03695_, _03693_);
  and (_03696_, _03674_, _03087_);
  and (_03698_, _03677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_04399_, _03698_, _03696_);
  and (_03699_, _02965_, _02064_);
  and (_03701_, _03699_, _03372_);
  and (_03702_, _03701_, _02963_);
  and (_03703_, _03702_, _03060_);
  not (_03705_, _03702_);
  and (_03706_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_04406_, _03706_, _03703_);
  and (_03708_, _03702_, _03067_);
  and (_03709_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_04409_, _03709_, _03708_);
  and (_03711_, _03702_, _03071_);
  and (_03712_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_04412_, _03712_, _03711_);
  and (_03714_, _03702_, _03074_);
  and (_03715_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_04415_, _03715_, _03714_);
  and (_03717_, _03702_, _03077_);
  and (_03718_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_04418_, _03718_, _03717_);
  and (_03719_, _03702_, _03080_);
  and (_03721_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_04421_, _03721_, _03719_);
  and (_03722_, _03702_, _03083_);
  and (_03724_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_04424_, _03724_, _03722_);
  and (_03725_, _03702_, _03087_);
  and (_03727_, _03705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_04427_, _03727_, _03725_);
  and (_03728_, _03701_, _03062_);
  and (_03730_, _03728_, _03060_);
  not (_03731_, _03728_);
  and (_03732_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or (_04430_, _03732_, _03730_);
  and (_03734_, _03728_, _03067_);
  and (_03735_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or (_04433_, _03735_, _03734_);
  and (_03737_, _03728_, _03071_);
  and (_03738_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or (_04436_, _03738_, _03737_);
  and (_03740_, _03728_, _03074_);
  and (_03742_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or (_04439_, _03742_, _03740_);
  and (_03743_, _03728_, _03077_);
  and (_03744_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or (_04442_, _03744_, _03743_);
  and (_03746_, _03728_, _03080_);
  and (_03747_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or (_04445_, _03747_, _03746_);
  and (_03749_, _03728_, _03083_);
  and (_03750_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or (_04448_, _03750_, _03749_);
  and (_03752_, _03728_, _03087_);
  and (_03753_, _03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or (_04451_, _03753_, _03752_);
  and (_03755_, _03701_, _03091_);
  and (_03756_, _03755_, _03060_);
  not (_03757_, _03755_);
  and (_03759_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or (_04455_, _03759_, _03756_);
  and (_03760_, _03755_, _03067_);
  and (_03762_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or (_04458_, _03762_, _03760_);
  and (_03763_, _03755_, _03071_);
  and (_03765_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or (_04461_, _03765_, _03763_);
  and (_03767_, _03755_, _03074_);
  and (_03768_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or (_04464_, _03768_, _03767_);
  and (_03769_, _03755_, _03077_);
  and (_03770_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or (_04467_, _03770_, _03769_);
  and (_03772_, _03755_, _03080_);
  and (_03773_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or (_04470_, _03773_, _03772_);
  and (_03775_, _03755_, _03083_);
  and (_03776_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or (_04473_, _03776_, _03775_);
  and (_03778_, _03755_, _03087_);
  and (_03779_, _03757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or (_04475_, _03779_, _03778_);
  and (_03781_, _03701_, _03113_);
  and (_03783_, _03781_, _03060_);
  not (_03785_, _03781_);
  and (_03786_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_04480_, _03786_, _03783_);
  and (_03788_, _03781_, _03067_);
  and (_03789_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_04483_, _03789_, _03788_);
  and (_03791_, _03781_, _03071_);
  and (_03792_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_04486_, _03792_, _03791_);
  and (_03794_, _03781_, _03074_);
  and (_03795_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_04489_, _03795_, _03794_);
  and (_03796_, _03781_, _03077_);
  and (_03797_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_04492_, _03797_, _03796_);
  and (_03798_, _03781_, _03080_);
  and (_03800_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_04495_, _03800_, _03798_);
  and (_03801_, _03781_, _03083_);
  and (_03803_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_04498_, _03803_, _03801_);
  and (_03804_, _03781_, _03087_);
  and (_03806_, _03785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_04501_, _03806_, _03804_);
  and (_03807_, _03701_, _03136_);
  and (_03809_, _03807_, _03060_);
  not (_03810_, _03807_);
  and (_03811_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_04505_, _03811_, _03809_);
  and (_03813_, _03807_, _03067_);
  and (_03814_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_04508_, _03814_, _03813_);
  and (_03816_, _03807_, _03071_);
  and (_03817_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_04511_, _03817_, _03816_);
  and (_03819_, _03807_, _03074_);
  and (_03821_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_04514_, _03821_, _03819_);
  and (_03822_, _03807_, _03077_);
  and (_03823_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_04517_, _03823_, _03822_);
  and (_03825_, _03807_, _03080_);
  and (_03826_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_04520_, _03826_, _03825_);
  and (_03828_, _03807_, _03083_);
  and (_03829_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_04523_, _03829_, _03828_);
  and (_03831_, _03807_, _03087_);
  and (_03832_, _03810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_04526_, _03832_, _03831_);
  and (_03834_, _03701_, _03159_);
  and (_03835_, _03834_, _03060_);
  not (_03836_, _03834_);
  and (_03838_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or (_04529_, _03838_, _03835_);
  and (_03839_, _03834_, _03067_);
  and (_03841_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or (_04533_, _03841_, _03839_);
  and (_03842_, _03834_, _03071_);
  and (_03844_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or (_04536_, _03844_, _03842_);
  and (_03846_, _03834_, _03074_);
  and (_03847_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or (_04539_, _03847_, _03846_);
  and (_03848_, _03834_, _03077_);
  and (_03849_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or (_04542_, _03849_, _03848_);
  and (_03851_, _03834_, _03080_);
  and (_03852_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or (_04545_, _03852_, _03851_);
  and (_03854_, _03834_, _03083_);
  and (_03855_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or (_04548_, _03855_, _03854_);
  and (_03857_, _03834_, _03087_);
  and (_03858_, _03836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or (_04550_, _03858_, _03857_);
  and (_03860_, _03701_, _03179_);
  and (_03861_, _03860_, _03060_);
  not (_03863_, _03860_);
  and (_03864_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or (_04554_, _03864_, _03861_);
  and (_03866_, _03860_, _03067_);
  and (_03867_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or (_04557_, _03867_, _03866_);
  and (_03869_, _03860_, _03071_);
  and (_03870_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or (_04561_, _03870_, _03869_);
  and (_03872_, _03860_, _03074_);
  and (_03873_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or (_04565_, _03873_, _03872_);
  and (_03874_, _03860_, _03077_);
  and (_03876_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or (_04568_, _03876_, _03874_);
  and (_03877_, _03860_, _03080_);
  and (_03879_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or (_04571_, _03879_, _03877_);
  and (_03880_, _03860_, _03083_);
  and (_03882_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or (_04574_, _03882_, _03880_);
  and (_03883_, _03860_, _03087_);
  and (_03885_, _03863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or (_04576_, _03885_, _03883_);
  and (_03886_, _03701_, _03198_);
  and (_03888_, _03886_, _03060_);
  not (_03889_, _03886_);
  and (_03890_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_04580_, _03890_, _03888_);
  and (_03892_, _03886_, _03067_);
  and (_03893_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_04583_, _03893_, _03892_);
  and (_03895_, _03886_, _03071_);
  and (_03897_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_04586_, _03897_, _03895_);
  and (_03898_, _03886_, _03074_);
  and (_03899_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_04589_, _03899_, _03898_);
  and (_03900_, _03886_, _03077_);
  and (_03902_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_04592_, _03902_, _03900_);
  and (_03903_, _03886_, _03080_);
  and (_03905_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_04595_, _03905_, _03903_);
  and (_03906_, _03886_, _03083_);
  and (_03908_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_04598_, _03908_, _03906_);
  and (_03909_, _03886_, _03087_);
  and (_03911_, _03889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_04601_, _03911_, _03909_);
  and (_03912_, _03701_, _03218_);
  and (_03914_, _03912_, _03060_);
  not (_03915_, _03912_);
  and (_03916_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or (_04605_, _03916_, _03914_);
  and (_03918_, _03912_, _03067_);
  and (_03919_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or (_04608_, _03919_, _03918_);
  and (_03921_, _03912_, _03071_);
  and (_03923_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or (_04611_, _03923_, _03921_);
  and (_03924_, _03912_, _03074_);
  and (_03925_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or (_04614_, _03925_, _03924_);
  and (_03927_, _03912_, _03077_);
  and (_03928_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or (_04618_, _03928_, _03927_);
  and (_03930_, _03912_, _03080_);
  and (_03931_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or (_04621_, _03931_, _03930_);
  and (_03933_, _03912_, _03083_);
  and (_03934_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or (_04624_, _03934_, _03933_);
  and (_03936_, _03912_, _03087_);
  and (_03937_, _03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or (_04626_, _03937_, _03936_);
  and (_03939_, _03701_, _03237_);
  and (_03940_, _03939_, _03060_);
  not (_03941_, _03939_);
  and (_03943_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_04630_, _03943_, _03940_);
  and (_03944_, _03939_, _03067_);
  and (_03946_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_04633_, _03946_, _03944_);
  and (_03948_, _03939_, _03071_);
  and (_03949_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_04636_, _03949_, _03948_);
  and (_03950_, _03939_, _03074_);
  and (_03951_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_04639_, _03951_, _03950_);
  and (_03953_, _03939_, _03077_);
  and (_03954_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_04642_, _03954_, _03953_);
  and (_03956_, _03939_, _03080_);
  and (_03957_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_04646_, _03957_, _03956_);
  and (_03959_, _03939_, _03083_);
  and (_03960_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_04649_, _03960_, _03959_);
  and (_03962_, _03939_, _03087_);
  and (_03963_, _03941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_04651_, _03963_, _03962_);
  and (_03965_, _03701_, _03256_);
  and (_03966_, _03965_, _03060_);
  not (_03968_, _03965_);
  and (_03969_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_04655_, _03969_, _03966_);
  and (_03971_, _03965_, _03067_);
  and (_03972_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_04658_, _03972_, _03971_);
  and (_03974_, _03965_, _03071_);
  and (_03975_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_04661_, _03975_, _03974_);
  and (_03976_, _03965_, _03074_);
  and (_03978_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_04664_, _03978_, _03976_);
  and (_03979_, _03965_, _03077_);
  and (_03981_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_04667_, _03981_, _03979_);
  and (_03982_, _03965_, _03080_);
  and (_03984_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_04670_, _03984_, _03982_);
  and (_03986_, _03965_, _03083_);
  and (_03988_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_04673_, _03988_, _03986_);
  and (_03989_, _03965_, _03087_);
  and (_03991_, _03968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_04676_, _03991_, _03989_);
  and (_03992_, _03701_, _03275_);
  and (_03994_, _03992_, _03060_);
  not (_03995_, _03992_);
  and (_03996_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or (_04679_, _03996_, _03994_);
  and (_03998_, _03992_, _03067_);
  and (_04000_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or (_04682_, _04000_, _03998_);
  and (_04001_, _03992_, _03071_);
  and (_04002_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or (_04685_, _04002_, _04001_);
  and (_04003_, _03992_, _03074_);
  and (_04004_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or (_04688_, _04004_, _04003_);
  and (_04006_, _03992_, _03077_);
  and (_04007_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or (_04691_, _04007_, _04006_);
  and (_04009_, _03992_, _03080_);
  and (_04010_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_04694_, _04010_, _04009_);
  and (_04012_, _03992_, _03083_);
  and (_04013_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or (_04698_, _04013_, _04012_);
  and (_04015_, _03992_, _03087_);
  and (_04016_, _03995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or (_04700_, _04016_, _04015_);
  and (_04018_, _03701_, _03295_);
  and (_04019_, _04018_, _03060_);
  not (_04020_, _04018_);
  and (_04022_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or (_04704_, _04022_, _04019_);
  and (_04023_, _04018_, _03067_);
  and (_04025_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or (_04708_, _04025_, _04023_);
  and (_04027_, _04018_, _03071_);
  and (_04028_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or (_04711_, _04028_, _04027_);
  and (_04029_, _04018_, _03074_);
  and (_04031_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or (_04714_, _04031_, _04029_);
  and (_04032_, _04018_, _03077_);
  and (_04034_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or (_04717_, _04034_, _04032_);
  and (_04035_, _04018_, _03080_);
  and (_04037_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or (_04720_, _04037_, _04035_);
  and (_04038_, _04018_, _03083_);
  and (_04040_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or (_04723_, _04040_, _04038_);
  and (_04041_, _04018_, _03087_);
  and (_04043_, _04020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_04726_, _04043_, _04041_);
  and (_04044_, _03701_, _03315_);
  and (_04046_, _04044_, _03060_);
  not (_04047_, _04044_);
  and (_04048_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_04730_, _04048_, _04046_);
  and (_04050_, _04044_, _03067_);
  and (_04052_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_04733_, _04052_, _04050_);
  and (_04053_, _04044_, _03071_);
  and (_04054_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_04736_, _04054_, _04053_);
  and (_04056_, _04044_, _03074_);
  and (_04057_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_04739_, _04057_, _04056_);
  and (_04059_, _04044_, _03077_);
  and (_04060_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_04742_, _04060_, _04059_);
  and (_04062_, _04044_, _03080_);
  and (_04063_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_04745_, _04063_, _04062_);
  and (_04065_, _04044_, _03083_);
  and (_04066_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_04748_, _04066_, _04065_);
  and (_04068_, _04044_, _03087_);
  and (_04069_, _04047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_04750_, _04069_, _04068_);
  and (_04071_, _03701_, _03334_);
  and (_04072_, _04071_, _03060_);
  not (_04074_, _04071_);
  and (_04075_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_04754_, _04075_, _04072_);
  and (_04077_, _04071_, _03067_);
  and (_04078_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_04757_, _04078_, _04077_);
  and (_04080_, _04071_, _03071_);
  and (_04081_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_04760_, _04081_, _04080_);
  and (_04083_, _04071_, _03074_);
  and (_04084_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_04763_, _04084_, _04083_);
  and (_04086_, _04071_, _03077_);
  and (_04087_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_04766_, _04087_, _04086_);
  and (_04089_, _04071_, _03080_);
  and (_04090_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_04769_, _04090_, _04089_);
  and (_04092_, _04071_, _03083_);
  and (_04093_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_04772_, _04093_, _04092_);
  and (_04095_, _04071_, _03087_);
  and (_04096_, _04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_04775_, _04096_, _04095_);
  and (_04098_, _03701_, _03353_);
  and (_04099_, _04098_, _03060_);
  not (_04101_, _04098_);
  and (_04102_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or (_04779_, _04102_, _04099_);
  and (_04103_, _04098_, _03067_);
  and (_04105_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or (_04782_, _04105_, _04103_);
  and (_04106_, _04098_, _03071_);
  and (_04108_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or (_04785_, _04108_, _04106_);
  and (_04109_, _04098_, _03074_);
  and (_04111_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or (_04788_, _04111_, _04109_);
  and (_04112_, _04098_, _03077_);
  and (_04114_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or (_04791_, _04114_, _04112_);
  and (_04115_, _04098_, _03080_);
  and (_04117_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_04794_, _04117_, _04115_);
  and (_04118_, _04098_, _03083_);
  and (_04120_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or (_04797_, _04120_, _04118_);
  and (_04121_, _04098_, _03087_);
  and (_04123_, _04101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_04799_, _04123_, _04121_);
  and (_04125_, _02965_, _02964_);
  and (_04126_, _04125_, _03372_);
  and (_04127_, _04126_, _02963_);
  and (_04128_, _04127_, _03060_);
  not (_04130_, _04127_);
  and (_04131_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or (_04805_, _04131_, _04128_);
  and (_04133_, _04127_, _03067_);
  and (_04134_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  or (_04808_, _04134_, _04133_);
  and (_04136_, _04127_, _03071_);
  and (_04137_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or (_04812_, _04137_, _04136_);
  and (_04139_, _04127_, _03074_);
  and (_04140_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  or (_04815_, _04140_, _04139_);
  and (_04142_, _04127_, _03077_);
  and (_04143_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or (_04818_, _04143_, _04142_);
  and (_04145_, _04127_, _03080_);
  and (_04146_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or (_04821_, _04146_, _04145_);
  and (_04148_, _04127_, _03083_);
  and (_04149_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  or (_04824_, _04149_, _04148_);
  and (_04151_, _04127_, _03087_);
  and (_04152_, _04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  or (_04826_, _04152_, _04151_);
  and (_04154_, _04126_, _03062_);
  and (_04155_, _04154_, _03060_);
  not (_04156_, _04154_);
  and (_04158_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_04830_, _04158_, _04155_);
  and (_04159_, _04154_, _03067_);
  and (_04161_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_04834_, _04161_, _04159_);
  and (_04162_, _04154_, _03071_);
  and (_04164_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_04837_, _04164_, _04162_);
  and (_04165_, _04154_, _03074_);
  and (_04167_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_04840_, _04167_, _04165_);
  and (_04168_, _04154_, _03077_);
  and (_04170_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_04843_, _04170_, _04168_);
  and (_04171_, _04154_, _03080_);
  and (_04173_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_04846_, _04173_, _04171_);
  and (_04175_, _04154_, _03083_);
  and (_04176_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_04849_, _04176_, _04175_);
  and (_04177_, _04154_, _03087_);
  and (_04179_, _04156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_04851_, _04179_, _04177_);
  and (_04180_, _04126_, _03091_);
  and (_04182_, _04180_, _03060_);
  not (_04183_, _04180_);
  and (_04184_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_04855_, _04184_, _04182_);
  and (_04186_, _04180_, _03067_);
  and (_04187_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_04858_, _04187_, _04186_);
  and (_04189_, _04180_, _03071_);
  and (_04191_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_04861_, _04191_, _04189_);
  and (_04193_, _04180_, _03074_);
  and (_04194_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_04864_, _04194_, _04193_);
  and (_04196_, _04180_, _03077_);
  and (_04197_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_04867_, _04197_, _04196_);
  and (_04199_, _04180_, _03080_);
  and (_04201_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_04870_, _04201_, _04199_);
  and (_04202_, _04180_, _03083_);
  and (_04203_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_04873_, _04203_, _04202_);
  and (_04205_, _04180_, _03087_);
  and (_04206_, _04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_04876_, _04206_, _04205_);
  and (_04208_, _04126_, _03113_);
  and (_04209_, _04208_, _03060_);
  not (_04211_, _04208_);
  and (_04212_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or (_04879_, _04212_, _04209_);
  and (_04214_, _04208_, _03067_);
  and (_04215_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or (_04882_, _04215_, _04214_);
  and (_04217_, _04208_, _03071_);
  and (_04218_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or (_04886_, _04218_, _04217_);
  and (_04220_, _04208_, _03074_);
  and (_04221_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or (_04889_, _04221_, _04220_);
  and (_04223_, _04208_, _03077_);
  and (_04224_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or (_04892_, _04224_, _04223_);
  and (_04226_, _04208_, _03080_);
  and (_04227_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or (_04895_, _04227_, _04226_);
  and (_04229_, _04208_, _03083_);
  and (_04230_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or (_04898_, _04230_, _04229_);
  and (_04232_, _04208_, _03087_);
  and (_04233_, _04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or (_04900_, _04233_, _04232_);
  and (_04235_, _04126_, _03136_);
  and (_04236_, _04235_, _03060_);
  not (_04237_, _04235_);
  and (_04239_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or (_04904_, _04239_, _04236_);
  and (_04240_, _04235_, _03067_);
  and (_04242_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or (_04907_, _04242_, _04240_);
  and (_04243_, _04235_, _03071_);
  and (_04245_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or (_04910_, _04245_, _04243_);
  and (_04246_, _04235_, _03074_);
  and (_04248_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or (_04915_, _04248_, _04246_);
  and (_04250_, _04235_, _03077_);
  and (_04251_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or (_04918_, _04251_, _04250_);
  and (_04252_, _04235_, _03080_);
  and (_04254_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or (_04921_, _04254_, _04252_);
  and (_04255_, _04235_, _03083_);
  and (_04257_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or (_04924_, _04257_, _04255_);
  and (_04258_, _04235_, _03087_);
  and (_04260_, _04237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_04926_, _04260_, _04258_);
  and (_04261_, _04126_, _03159_);
  and (_04263_, _04261_, _03060_);
  not (_04264_, _04261_);
  and (_04265_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_04930_, _04265_, _04263_);
  and (_04267_, _04261_, _03067_);
  and (_04268_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_04933_, _04268_, _04267_);
  and (_04270_, _04261_, _03071_);
  and (_04271_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_04936_, _04271_, _04270_);
  and (_04273_, _04261_, _03074_);
  and (_04275_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_04939_, _04275_, _04273_);
  and (_04276_, _04261_, _03077_);
  and (_04277_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_04942_, _04277_, _04276_);
  and (_04279_, _04261_, _03080_);
  and (_04280_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_04945_, _04280_, _04279_);
  and (_04282_, _04261_, _03083_);
  and (_04283_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_04948_, _04283_, _04282_);
  and (_04285_, _04261_, _03087_);
  and (_04286_, _04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_04951_, _04286_, _04285_);
  and (_04288_, _04126_, _03179_);
  and (_04289_, _04288_, _03060_);
  not (_04291_, _04288_);
  and (_04292_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_04954_, _04292_, _04289_);
  and (_04295_, _04288_, _03067_);
  and (_04296_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_04957_, _04296_, _04295_);
  and (_04298_, _04288_, _03071_);
  and (_04299_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_04960_, _04299_, _04298_);
  and (_04301_, _04288_, _03074_);
  and (_04302_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_04963_, _04302_, _04301_);
  and (_04304_, _04288_, _03077_);
  and (_04305_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_04967_, _04305_, _04304_);
  and (_04307_, _04288_, _03080_);
  and (_04308_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_04970_, _04308_, _04307_);
  and (_04310_, _04288_, _03083_);
  and (_04311_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_04973_, _04311_, _04310_);
  and (_04313_, _04288_, _03087_);
  and (_04314_, _04291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_04975_, _04314_, _04313_);
  and (_04316_, _04126_, _03198_);
  and (_04317_, _04316_, _03060_);
  not (_04318_, _04316_);
  and (_04320_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or (_04979_, _04320_, _04317_);
  and (_04321_, _04316_, _03067_);
  and (_04323_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or (_04982_, _04323_, _04321_);
  and (_04325_, _04316_, _03071_);
  and (_04326_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or (_04985_, _04326_, _04325_);
  and (_04327_, _04316_, _03074_);
  and (_04329_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or (_04988_, _04329_, _04327_);
  and (_04330_, _04316_, _03077_);
  and (_04332_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or (_04991_, _04332_, _04330_);
  and (_04333_, _04316_, _03080_);
  and (_04335_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or (_04995_, _04335_, _04333_);
  and (_04336_, _04316_, _03083_);
  and (_04338_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or (_04998_, _04338_, _04336_);
  and (_04339_, _04316_, _03087_);
  and (_04341_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or (_05000_, _04341_, _04339_);
  and (_04342_, _04126_, _03218_);
  and (_04344_, _04342_, _03060_);
  not (_04345_, _04342_);
  and (_04346_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_05004_, _04346_, _04344_);
  and (_04348_, _04342_, _03067_);
  and (_04350_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_05007_, _04350_, _04348_);
  and (_04351_, _04342_, _03071_);
  and (_04352_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_05010_, _04352_, _04351_);
  and (_04354_, _04342_, _03074_);
  and (_04355_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_05013_, _04355_, _04354_);
  and (_04357_, _04342_, _03077_);
  and (_04358_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_05016_, _04358_, _04357_);
  and (_04360_, _04342_, _03080_);
  and (_04361_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_05019_, _04361_, _04360_);
  and (_04363_, _04342_, _03083_);
  and (_04364_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_05023_, _04364_, _04363_);
  and (_04366_, _04342_, _03087_);
  and (_04367_, _04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_05025_, _04367_, _04366_);
  and (_04369_, _04126_, _03237_);
  and (_04370_, _04369_, _03060_);
  not (_04372_, _04369_);
  and (_04373_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or (_05029_, _04373_, _04370_);
  and (_04375_, _04369_, _03067_);
  and (_04376_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or (_05032_, _04376_, _04375_);
  and (_04378_, _04369_, _03071_);
  and (_04379_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or (_05035_, _04379_, _04378_);
  and (_04381_, _04369_, _03074_);
  and (_04382_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or (_05038_, _04382_, _04381_);
  and (_04384_, _04369_, _03077_);
  and (_04385_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or (_05041_, _04385_, _04384_);
  and (_04387_, _04369_, _03080_);
  and (_04388_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or (_05044_, _04388_, _04387_);
  and (_04390_, _04369_, _03083_);
  and (_04391_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or (_05047_, _04391_, _04390_);
  and (_04393_, _04369_, _03087_);
  and (_04394_, _04372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or (_05050_, _04394_, _04393_);
  and (_04396_, _04126_, _03256_);
  and (_04398_, _04396_, _03060_);
  not (_04400_, _04396_);
  and (_04401_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or (_05053_, _04401_, _04398_);
  and (_04402_, _04396_, _03067_);
  and (_04403_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or (_05056_, _04403_, _04402_);
  and (_04404_, _04396_, _03071_);
  and (_04405_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or (_05059_, _04405_, _04404_);
  and (_04407_, _04396_, _03074_);
  and (_04408_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or (_05062_, _04408_, _04407_);
  and (_04410_, _04396_, _03077_);
  and (_04411_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or (_05065_, _04411_, _04410_);
  and (_04413_, _04396_, _03080_);
  and (_04414_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or (_05068_, _04414_, _04413_);
  and (_04416_, _04396_, _03083_);
  and (_04417_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or (_05071_, _04417_, _04416_);
  and (_04419_, _04396_, _03087_);
  and (_04420_, _04400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or (_05074_, _04420_, _04419_);
  and (_04422_, _04126_, _03275_);
  and (_04423_, _04422_, _03060_);
  not (_04425_, _04422_);
  and (_04426_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_05078_, _04426_, _04423_);
  and (_04428_, _04422_, _03067_);
  and (_04429_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_05081_, _04429_, _04428_);
  and (_04431_, _04422_, _03071_);
  and (_04432_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_05084_, _04432_, _04431_);
  and (_04434_, _04422_, _03074_);
  and (_04435_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_05087_, _04435_, _04434_);
  and (_04437_, _04422_, _03077_);
  and (_04438_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_05090_, _04438_, _04437_);
  and (_04440_, _04422_, _03080_);
  and (_04441_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_05093_, _04441_, _04440_);
  and (_04443_, _04422_, _03083_);
  and (_04444_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_05096_, _04444_, _04443_);
  and (_04446_, _04422_, _03087_);
  and (_04447_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_05098_, _04447_, _04446_);
  and (_04449_, _04126_, _03295_);
  and (_04450_, _04449_, _03060_);
  not (_04452_, _04449_);
  and (_04453_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_05103_, _04453_, _04450_);
  and (_04454_, _04449_, _03067_);
  and (_04456_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_05106_, _04456_, _04454_);
  and (_04457_, _04449_, _03071_);
  and (_04459_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_05109_, _04459_, _04457_);
  and (_04460_, _04449_, _03074_);
  and (_04462_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_05112_, _04462_, _04460_);
  and (_04463_, _04449_, _03077_);
  and (_04465_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_05115_, _04465_, _04463_);
  and (_04466_, _04449_, _03080_);
  and (_04468_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_05118_, _04468_, _04466_);
  and (_04469_, _04449_, _03083_);
  and (_04471_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_05121_, _04471_, _04469_);
  and (_04472_, _04449_, _03087_);
  and (_04474_, _04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_05123_, _04474_, _04472_);
  and (_04476_, _04126_, _03315_);
  and (_04477_, _04476_, _03060_);
  not (_04478_, _04476_);
  and (_04479_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or (_05127_, _04479_, _04477_);
  and (_04481_, _04476_, _03067_);
  and (_04482_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or (_05130_, _04482_, _04481_);
  and (_04484_, _04476_, _03071_);
  and (_04485_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or (_05133_, _04485_, _04484_);
  and (_04487_, _04476_, _03074_);
  and (_04488_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or (_05136_, _04488_, _04487_);
  and (_04490_, _04476_, _03077_);
  and (_04491_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or (_05139_, _04491_, _04490_);
  and (_04493_, _04476_, _03080_);
  and (_04494_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or (_05142_, _04494_, _04493_);
  and (_04496_, _04476_, _03083_);
  and (_04497_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or (_05145_, _04497_, _04496_);
  and (_04500_, _04476_, _03087_);
  and (_04502_, _04478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or (_05148_, _04502_, _04500_);
  and (_04503_, _04126_, _03334_);
  and (_04504_, _04503_, _03060_);
  not (_04506_, _04503_);
  and (_04507_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or (_05151_, _04507_, _04504_);
  and (_04509_, _04503_, _03067_);
  and (_04510_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or (_05155_, _04510_, _04509_);
  and (_04512_, _04503_, _03071_);
  and (_04513_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or (_05158_, _04513_, _04512_);
  and (_04515_, _04503_, _03074_);
  and (_04516_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or (_05161_, _04516_, _04515_);
  and (_04518_, _04503_, _03077_);
  and (_04519_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or (_05164_, _04519_, _04518_);
  and (_04521_, _04503_, _03080_);
  and (_04522_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or (_05167_, _04522_, _04521_);
  and (_04524_, _04503_, _03083_);
  and (_04525_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or (_05170_, _04525_, _04524_);
  and (_04527_, _04503_, _03087_);
  and (_04528_, _04506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or (_05172_, _04528_, _04527_);
  and (_04530_, _04126_, _03353_);
  and (_04531_, _04530_, _03060_);
  not (_04532_, _04530_);
  and (_04534_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_05176_, _04534_, _04531_);
  and (_04535_, _04530_, _03067_);
  and (_04537_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_05179_, _04537_, _04535_);
  and (_04538_, _04530_, _03071_);
  and (_04540_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_05183_, _04540_, _04538_);
  and (_04541_, _04530_, _03074_);
  and (_04543_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_05186_, _04543_, _04541_);
  and (_04544_, _04530_, _03077_);
  and (_04546_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_05189_, _04546_, _04544_);
  and (_04547_, _04530_, _03080_);
  and (_04549_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_05192_, _04549_, _04547_);
  and (_04551_, _04530_, _03083_);
  and (_04552_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_05195_, _04552_, _04551_);
  and (_04553_, _04530_, _03087_);
  and (_04555_, _04532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_05197_, _04555_, _04553_);
  and (_04556_, _25446_, _25101_);
  and (_04558_, _04556_, _02008_);
  and (_04559_, _04558_, _02966_);
  and (_04560_, _04559_, _02963_);
  and (_04562_, _04560_, _03060_);
  not (_04563_, _04560_);
  and (_04564_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_05203_, _04564_, _04562_);
  and (_04566_, _04560_, _03067_);
  and (_04567_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_05207_, _04567_, _04566_);
  and (_04569_, _04560_, _03071_);
  and (_04570_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_05210_, _04570_, _04569_);
  and (_04572_, _04560_, _03074_);
  and (_04573_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_05213_, _04573_, _04572_);
  and (_04575_, _04560_, _03077_);
  and (_04577_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_05216_, _04577_, _04575_);
  and (_04578_, _04560_, _03080_);
  and (_04579_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_05219_, _04579_, _04578_);
  and (_04581_, _04560_, _03083_);
  and (_04582_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_05222_, _04582_, _04581_);
  and (_04584_, _04560_, _03087_);
  and (_04585_, _04563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_05224_, _04585_, _04584_);
  and (_04587_, _04559_, _03062_);
  and (_04588_, _04587_, _03060_);
  not (_04590_, _04587_);
  and (_04591_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_05228_, _04591_, _04588_);
  and (_04593_, _04587_, _03067_);
  and (_04594_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_05231_, _04594_, _04593_);
  and (_04596_, _04587_, _03071_);
  and (_04597_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_05235_, _04597_, _04596_);
  and (_04599_, _04587_, _03074_);
  and (_04600_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_05238_, _04600_, _04599_);
  and (_04602_, _04587_, _03077_);
  and (_04603_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_05241_, _04603_, _04602_);
  and (_04606_, _04587_, _03080_);
  and (_04607_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or (_05244_, _04607_, _04606_);
  and (_04609_, _04587_, _03083_);
  and (_04610_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or (_05247_, _04610_, _04609_);
  and (_04612_, _04587_, _03087_);
  and (_04613_, _04590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or (_05249_, _04613_, _04612_);
  and (_04615_, _04559_, _03091_);
  and (_04616_, _04615_, _03060_);
  not (_04617_, _04615_);
  and (_04619_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or (_05253_, _04619_, _04616_);
  and (_04620_, _04615_, _03067_);
  and (_04622_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_05256_, _04622_, _04620_);
  and (_04623_, _04615_, _03071_);
  and (_04625_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or (_05259_, _04625_, _04623_);
  and (_04627_, _04615_, _03074_);
  and (_04628_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or (_05262_, _04628_, _04627_);
  and (_04629_, _04615_, _03077_);
  and (_04631_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or (_05265_, _04631_, _04629_);
  and (_04632_, _04615_, _03080_);
  and (_04634_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or (_05268_, _04634_, _04632_);
  and (_04635_, _04615_, _03083_);
  and (_04637_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or (_05271_, _04637_, _04635_);
  and (_04638_, _04615_, _03087_);
  and (_04640_, _04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or (_05274_, _04640_, _04638_);
  and (_04641_, _04559_, _03113_);
  and (_04643_, _04641_, _03060_);
  not (_04644_, _04641_);
  and (_04645_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_05277_, _04645_, _04643_);
  and (_04647_, _04641_, _03067_);
  and (_04648_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_05280_, _04648_, _04647_);
  and (_04650_, _04641_, _03071_);
  and (_04652_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_05283_, _04652_, _04650_);
  and (_04653_, _04641_, _03074_);
  and (_04654_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_05287_, _04654_, _04653_);
  and (_04656_, _04641_, _03077_);
  and (_04657_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_05290_, _04657_, _04656_);
  and (_04659_, _04641_, _03080_);
  and (_04660_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_05293_, _04660_, _04659_);
  and (_04662_, _04641_, _03083_);
  and (_04663_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_05296_, _04663_, _04662_);
  and (_04665_, _04641_, _03087_);
  and (_04666_, _04644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_05298_, _04666_, _04665_);
  and (_04668_, _04559_, _03136_);
  and (_04669_, _04668_, _03060_);
  not (_04671_, _04668_);
  and (_04672_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_05302_, _04672_, _04669_);
  and (_04674_, _04668_, _03067_);
  and (_04675_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_05305_, _04675_, _04674_);
  and (_04677_, _04668_, _03071_);
  and (_04678_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_05308_, _04678_, _04677_);
  and (_04680_, _04668_, _03074_);
  and (_04681_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_05311_, _04681_, _04680_);
  and (_04683_, _04668_, _03077_);
  and (_04684_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_05315_, _04684_, _04683_);
  and (_04686_, _04668_, _03080_);
  and (_04687_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_05318_, _04687_, _04686_);
  and (_04689_, _04668_, _03083_);
  and (_04690_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_05321_, _04690_, _04689_);
  and (_04692_, _04668_, _03087_);
  and (_04693_, _04671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_05323_, _04693_, _04692_);
  and (_04695_, _04559_, _03159_);
  and (_04696_, _04695_, _03060_);
  not (_04697_, _04695_);
  and (_04699_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_05327_, _04699_, _04696_);
  and (_04701_, _04695_, _03067_);
  and (_04702_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_05330_, _04702_, _04701_);
  and (_04703_, _04695_, _03071_);
  and (_04705_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or (_05333_, _04705_, _04703_);
  and (_04706_, _04695_, _03074_);
  and (_04709_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_05336_, _04709_, _04706_);
  and (_04710_, _04695_, _03077_);
  and (_04712_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or (_05339_, _04712_, _04710_);
  and (_04713_, _04695_, _03080_);
  and (_04715_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_05342_, _04715_, _04713_);
  and (_04716_, _04695_, _03083_);
  and (_04718_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or (_05345_, _04718_, _04716_);
  and (_04719_, _04695_, _03087_);
  and (_04721_, _04697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_05348_, _04721_, _04719_);
  and (_04722_, _04559_, _03179_);
  and (_04724_, _04722_, _03060_);
  not (_04725_, _04722_);
  and (_04727_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or (_05351_, _04727_, _04724_);
  and (_04728_, _04722_, _03067_);
  and (_04729_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_05354_, _04729_, _04728_);
  and (_04731_, _04722_, _03071_);
  and (_04732_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_05357_, _04732_, _04731_);
  and (_04734_, _04722_, _03074_);
  and (_04735_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or (_05360_, _04735_, _04734_);
  and (_04737_, _04722_, _03077_);
  and (_04738_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_05363_, _04738_, _04737_);
  and (_04740_, _04722_, _03080_);
  and (_04741_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or (_05367_, _04741_, _04740_);
  and (_04743_, _04722_, _03083_);
  and (_04744_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or (_05370_, _04744_, _04743_);
  and (_04746_, _04722_, _03087_);
  and (_04747_, _04725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or (_05372_, _04747_, _04746_);
  and (_04749_, _04559_, _03198_);
  and (_04751_, _04749_, _03060_);
  not (_04752_, _04749_);
  and (_04753_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_05376_, _04753_, _04751_);
  and (_04755_, _04749_, _03067_);
  and (_04756_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_05379_, _04756_, _04755_);
  and (_04758_, _04749_, _03071_);
  and (_04759_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_05382_, _04759_, _04758_);
  and (_04761_, _04749_, _03074_);
  and (_04762_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_05385_, _04762_, _04761_);
  and (_04764_, _04749_, _03077_);
  and (_04765_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_05388_, _04765_, _04764_);
  and (_04767_, _04749_, _03080_);
  and (_04768_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_05391_, _04768_, _04767_);
  and (_04770_, _04749_, _03083_);
  and (_04771_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_05395_, _04771_, _04770_);
  and (_04773_, _04749_, _03087_);
  and (_04774_, _04752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_05397_, _04774_, _04773_);
  and (_04776_, _04559_, _03218_);
  and (_04777_, _04776_, _03060_);
  not (_04778_, _04776_);
  and (_04780_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_05401_, _04780_, _04777_);
  and (_04781_, _04776_, _03067_);
  and (_04783_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_05404_, _04783_, _04781_);
  and (_04784_, _04776_, _03071_);
  and (_04786_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or (_05407_, _04786_, _04784_);
  and (_04787_, _04776_, _03074_);
  and (_04789_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_05410_, _04789_, _04787_);
  and (_04790_, _04776_, _03077_);
  and (_04792_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_05413_, _04792_, _04790_);
  and (_04793_, _04776_, _03080_);
  and (_04795_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_05416_, _04795_, _04793_);
  and (_04796_, _04776_, _03083_);
  and (_04798_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or (_05419_, _04798_, _04796_);
  and (_04800_, _04776_, _03087_);
  and (_04801_, _04778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or (_05422_, _04801_, _04800_);
  and (_04802_, _04559_, _03237_);
  and (_04803_, _04802_, _03060_);
  not (_04804_, _04802_);
  and (_04806_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_05426_, _04806_, _04803_);
  and (_04807_, _04802_, _03067_);
  and (_04809_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_05429_, _04809_, _04807_);
  and (_04811_, _04802_, _03071_);
  and (_04813_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_05432_, _04813_, _04811_);
  and (_04814_, _04802_, _03074_);
  and (_04816_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_05435_, _04816_, _04814_);
  and (_04817_, _04802_, _03077_);
  and (_04819_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_05438_, _04819_, _04817_);
  and (_04820_, _04802_, _03080_);
  and (_04822_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_05441_, _04822_, _04820_);
  and (_04823_, _04802_, _03083_);
  and (_04825_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_05444_, _04825_, _04823_);
  and (_04827_, _04802_, _03087_);
  and (_04828_, _04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_05446_, _04828_, _04827_);
  and (_04829_, _04559_, _03256_);
  and (_04831_, _04829_, _03060_);
  not (_04832_, _04829_);
  and (_04833_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_05450_, _04833_, _04831_);
  and (_04835_, _04829_, _03067_);
  and (_04836_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_05453_, _04836_, _04835_);
  and (_04838_, _04829_, _03071_);
  and (_04839_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_05456_, _04839_, _04838_);
  and (_04841_, _04829_, _03074_);
  and (_04842_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_05459_, _04842_, _04841_);
  and (_04844_, _04829_, _03077_);
  and (_04845_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_05462_, _04845_, _04844_);
  and (_04847_, _04829_, _03080_);
  and (_04848_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_05465_, _04848_, _04847_);
  and (_04850_, _04829_, _03083_);
  and (_04852_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_05468_, _04852_, _04850_);
  and (_04853_, _04829_, _03087_);
  and (_04854_, _04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_05471_, _04854_, _04853_);
  and (_04856_, _04559_, _03275_);
  and (_04857_, _04856_, _03060_);
  not (_04859_, _04856_);
  and (_04860_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or (_05475_, _04860_, _04857_);
  and (_04862_, _04856_, _03067_);
  and (_04863_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_05478_, _04863_, _04862_);
  and (_04865_, _04856_, _03071_);
  and (_04866_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_05481_, _04866_, _04865_);
  and (_04868_, _04856_, _03074_);
  and (_04869_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or (_05484_, _04869_, _04868_);
  and (_04871_, _04856_, _03077_);
  and (_04872_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_05487_, _04872_, _04871_);
  and (_04874_, _04856_, _03080_);
  and (_04875_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or (_05490_, _04875_, _04874_);
  and (_04877_, _04856_, _03083_);
  and (_04878_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or (_05493_, _04878_, _04877_);
  and (_04880_, _04856_, _03087_);
  and (_04881_, _04859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_05495_, _04881_, _04880_);
  and (_04883_, _04559_, _03295_);
  and (_04884_, _04883_, _03060_);
  not (_04885_, _04883_);
  and (_04887_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_05499_, _04887_, _04884_);
  and (_04888_, _04883_, _03067_);
  and (_04890_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_05503_, _04890_, _04888_);
  and (_04891_, _04883_, _03071_);
  and (_04893_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or (_05506_, _04893_, _04891_);
  and (_04894_, _04883_, _03074_);
  and (_04896_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_05509_, _04896_, _04894_);
  and (_04897_, _04883_, _03077_);
  and (_04899_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or (_05512_, _04899_, _04897_);
  and (_04901_, _04883_, _03080_);
  and (_04902_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or (_05515_, _04902_, _04901_);
  and (_04903_, _04883_, _03083_);
  and (_04905_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or (_05518_, _04905_, _04903_);
  and (_04906_, _04883_, _03087_);
  and (_04908_, _04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or (_05520_, _04908_, _04906_);
  and (_04909_, _04559_, _03315_);
  and (_04911_, _04909_, _03060_);
  not (_04912_, _04909_);
  and (_04913_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_05524_, _04913_, _04911_);
  and (_04916_, _04909_, _03067_);
  and (_04917_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_05527_, _04917_, _04916_);
  and (_04919_, _04909_, _03071_);
  and (_04920_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_05530_, _04920_, _04919_);
  and (_04922_, _04909_, _03074_);
  and (_04923_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_05533_, _04923_, _04922_);
  and (_04925_, _04909_, _03077_);
  and (_04927_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_05536_, _04927_, _04925_);
  and (_04928_, _04909_, _03080_);
  and (_04929_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_05539_, _04929_, _04928_);
  and (_04931_, _04909_, _03083_);
  and (_04932_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_05542_, _04932_, _04931_);
  and (_04934_, _04909_, _03087_);
  and (_04935_, _04912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_05545_, _04935_, _04934_);
  and (_04937_, _04559_, _03334_);
  and (_04938_, _04937_, _03060_);
  not (_04940_, _04937_);
  and (_04941_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_05548_, _04941_, _04938_);
  and (_04943_, _04937_, _03067_);
  and (_04944_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_05551_, _04944_, _04943_);
  and (_04946_, _04937_, _03071_);
  and (_04947_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_05555_, _04947_, _04946_);
  and (_04949_, _04937_, _03074_);
  and (_04950_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_05558_, _04950_, _04949_);
  and (_04952_, _04937_, _03077_);
  and (_04953_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_05561_, _04953_, _04952_);
  and (_04955_, _04937_, _03080_);
  and (_04956_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_05564_, _04956_, _04955_);
  and (_04958_, _04937_, _03083_);
  and (_04959_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_05567_, _04959_, _04958_);
  and (_04961_, _04937_, _03087_);
  and (_04962_, _04940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_05569_, _04962_, _04961_);
  and (_04964_, _04559_, _03353_);
  and (_04965_, _04964_, _03060_);
  not (_04966_, _04964_);
  and (_04968_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_05573_, _04968_, _04965_);
  and (_04969_, _04964_, _03067_);
  and (_04971_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_05576_, _04971_, _04969_);
  and (_04972_, _04964_, _03071_);
  and (_04974_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_05579_, _04974_, _04972_);
  and (_04976_, _04964_, _03074_);
  and (_04977_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_05583_, _04977_, _04976_);
  and (_04978_, _04964_, _03077_);
  and (_04980_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_05586_, _04980_, _04978_);
  and (_04981_, _04964_, _03080_);
  and (_04983_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or (_05589_, _04983_, _04981_);
  and (_04984_, _04964_, _03083_);
  and (_04986_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or (_05592_, _04986_, _04984_);
  and (_04987_, _04964_, _03087_);
  and (_04989_, _04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or (_05594_, _04989_, _04987_);
  and (_04990_, _04558_, _03373_);
  and (_04992_, _04990_, _02963_);
  and (_04993_, _04992_, _03060_);
  not (_04994_, _04992_);
  and (_04996_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or (_05598_, _04996_, _04993_);
  and (_04997_, _04992_, _03067_);
  and (_04999_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or (_05601_, _04999_, _04997_);
  and (_05001_, _04992_, _03071_);
  and (_05002_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or (_05604_, _05002_, _05001_);
  and (_05003_, _04992_, _03074_);
  and (_05005_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or (_05608_, _05005_, _05003_);
  and (_05006_, _04992_, _03077_);
  and (_05008_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or (_05611_, _05008_, _05006_);
  and (_05009_, _04992_, _03080_);
  and (_05011_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_05614_, _05011_, _05009_);
  and (_05012_, _04992_, _03083_);
  and (_05014_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or (_05617_, _05014_, _05012_);
  and (_05015_, _04992_, _03087_);
  and (_05017_, _04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_05619_, _05017_, _05015_);
  and (_05018_, _04990_, _03062_);
  and (_05020_, _05018_, _03060_);
  not (_05021_, _05018_);
  and (_05022_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_05623_, _05022_, _05020_);
  and (_05024_, _05018_, _03067_);
  and (_05026_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_05626_, _05026_, _05024_);
  and (_05027_, _05018_, _03071_);
  and (_05028_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_05629_, _05028_, _05027_);
  and (_05030_, _05018_, _03074_);
  and (_05031_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_05632_, _05031_, _05030_);
  and (_05033_, _05018_, _03077_);
  and (_05034_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_05636_, _05034_, _05033_);
  and (_05036_, _05018_, _03080_);
  and (_05037_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_05639_, _05037_, _05036_);
  and (_05039_, _05018_, _03083_);
  and (_05040_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_05642_, _05040_, _05039_);
  and (_05042_, _05018_, _03087_);
  and (_05043_, _05021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_05644_, _05043_, _05042_);
  and (_05045_, _04990_, _03091_);
  and (_05046_, _05045_, _03060_);
  not (_05048_, _05045_);
  and (_05049_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_05648_, _05049_, _05046_);
  and (_05051_, _05045_, _03067_);
  and (_05052_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_05651_, _05052_, _05051_);
  and (_05054_, _05045_, _03071_);
  and (_05055_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_05654_, _05055_, _05054_);
  and (_05057_, _05045_, _03074_);
  and (_05058_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_05657_, _05058_, _05057_);
  and (_05060_, _05045_, _03077_);
  and (_05061_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_05660_, _05061_, _05060_);
  and (_05063_, _05045_, _03080_);
  and (_05064_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_05663_, _05064_, _05063_);
  and (_05066_, _05045_, _03083_);
  and (_05067_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_05666_, _05067_, _05066_);
  and (_05069_, _05045_, _03087_);
  and (_05070_, _05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_05669_, _05070_, _05069_);
  and (_05072_, _04990_, _03113_);
  and (_05073_, _05072_, _03060_);
  not (_05075_, _05072_);
  and (_05076_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or (_05672_, _05076_, _05073_);
  and (_05077_, _05072_, _03067_);
  and (_05079_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or (_05675_, _05079_, _05077_);
  and (_05080_, _05072_, _03071_);
  and (_05082_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or (_05678_, _05082_, _05080_);
  and (_05083_, _05072_, _03074_);
  and (_05085_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or (_05681_, _05085_, _05083_);
  and (_05086_, _05072_, _03077_);
  and (_05088_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or (_05684_, _05088_, _05086_);
  and (_05089_, _05072_, _03080_);
  and (_05091_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or (_05688_, _05091_, _05089_);
  and (_05092_, _05072_, _03083_);
  and (_05094_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or (_05691_, _05094_, _05092_);
  and (_05095_, _05072_, _03087_);
  and (_05097_, _05075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_05693_, _05097_, _05095_);
  and (_05099_, _04990_, _03136_);
  and (_05100_, _05099_, _03060_);
  not (_05101_, _05099_);
  and (_05102_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or (_05697_, _05102_, _05100_);
  and (_05104_, _05099_, _03067_);
  and (_05105_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or (_05700_, _05105_, _05104_);
  and (_05107_, _05099_, _03071_);
  and (_05108_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or (_05703_, _05108_, _05107_);
  and (_05110_, _05099_, _03074_);
  and (_05111_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or (_05706_, _05111_, _05110_);
  and (_05113_, _05099_, _03077_);
  and (_05114_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or (_05709_, _05114_, _05113_);
  and (_05116_, _05099_, _03080_);
  and (_05117_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_05712_, _05117_, _05116_);
  and (_05119_, _05099_, _03083_);
  and (_05120_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or (_05716_, _05120_, _05119_);
  and (_05122_, _05099_, _03087_);
  and (_05124_, _05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or (_05718_, _05124_, _05122_);
  and (_05125_, _04990_, _03159_);
  and (_05126_, _05125_, _03060_);
  not (_05128_, _05125_);
  and (_05129_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_05722_, _05129_, _05126_);
  and (_05131_, _05125_, _03067_);
  and (_05132_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_05725_, _05132_, _05131_);
  and (_05134_, _05125_, _03071_);
  and (_05135_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_05728_, _05135_, _05134_);
  and (_05137_, _05125_, _03074_);
  and (_05138_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_05731_, _05138_, _05137_);
  and (_05140_, _05125_, _03077_);
  and (_05141_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_05734_, _05141_, _05140_);
  and (_05143_, _05125_, _03080_);
  and (_05144_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_05737_, _05144_, _05143_);
  and (_05146_, _05125_, _03083_);
  and (_05147_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_05740_, _05147_, _05146_);
  and (_05149_, _05125_, _03087_);
  and (_05150_, _05128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_05743_, _05150_, _05149_);
  and (_05152_, _04990_, _03179_);
  and (_05153_, _05152_, _03060_);
  not (_05154_, _05152_);
  and (_05156_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_05746_, _05156_, _05153_);
  and (_05157_, _05152_, _03067_);
  and (_05159_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_05749_, _05159_, _05157_);
  and (_05160_, _05152_, _03071_);
  and (_05162_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_05752_, _05162_, _05160_);
  and (_05163_, _05152_, _03074_);
  and (_05165_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_05755_, _05165_, _05163_);
  and (_05166_, _05152_, _03077_);
  and (_05168_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_05758_, _05168_, _05166_);
  and (_05169_, _05152_, _03080_);
  and (_05171_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_05761_, _05171_, _05169_);
  and (_05173_, _05152_, _03083_);
  and (_05174_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_05764_, _05174_, _05173_);
  and (_05175_, _05152_, _03087_);
  and (_05177_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_05767_, _05177_, _05175_);
  and (_05178_, _04990_, _03198_);
  and (_05180_, _05178_, _03060_);
  not (_05181_, _05178_);
  and (_05182_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or (_05771_, _05182_, _05180_);
  and (_05184_, _05178_, _03067_);
  and (_05185_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or (_05774_, _05185_, _05184_);
  and (_05187_, _05178_, _03071_);
  and (_05188_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or (_05777_, _05188_, _05187_);
  and (_05190_, _05178_, _03074_);
  and (_05191_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or (_05780_, _05191_, _05190_);
  and (_05193_, _05178_, _03077_);
  and (_05194_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or (_05783_, _05194_, _05193_);
  and (_05196_, _05178_, _03080_);
  and (_05198_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_05786_, _05198_, _05196_);
  and (_05199_, _05178_, _03083_);
  and (_05200_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or (_05789_, _05200_, _05199_);
  and (_05201_, _05178_, _03087_);
  and (_05202_, _05181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or (_05791_, _05202_, _05201_);
  and (_05204_, _04990_, _03218_);
  and (_05205_, _05204_, _03060_);
  not (_05206_, _05204_);
  and (_05208_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_05796_, _05208_, _05205_);
  and (_05209_, _05204_, _03067_);
  and (_05211_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_05799_, _05211_, _05209_);
  and (_05212_, _05204_, _03071_);
  and (_05214_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_05802_, _05214_, _05212_);
  and (_05215_, _05204_, _03074_);
  and (_05217_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_05805_, _05217_, _05215_);
  and (_05218_, _05204_, _03077_);
  and (_05220_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_05808_, _05220_, _05218_);
  and (_05221_, _05204_, _03080_);
  and (_05223_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_05811_, _05223_, _05221_);
  and (_05225_, _05204_, _03083_);
  and (_05226_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_05814_, _05226_, _05225_);
  and (_05227_, _05204_, _03087_);
  and (_05229_, _05206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_05816_, _05229_, _05227_);
  and (_05230_, _04990_, _03237_);
  and (_05232_, _05230_, _03060_);
  not (_05233_, _05230_);
  and (_05234_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or (_05820_, _05234_, _05232_);
  and (_05236_, _05230_, _03067_);
  and (_05237_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or (_05823_, _05237_, _05236_);
  and (_05239_, _05230_, _03071_);
  and (_05240_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or (_05826_, _05240_, _05239_);
  and (_05242_, _05230_, _03074_);
  and (_05243_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or (_05829_, _05243_, _05242_);
  and (_05245_, _05230_, _03077_);
  and (_05246_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or (_05832_, _05246_, _05245_);
  and (_05248_, _05230_, _03080_);
  and (_05250_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or (_05835_, _05250_, _05248_);
  and (_05251_, _05230_, _03083_);
  and (_05252_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or (_05838_, _05252_, _05251_);
  and (_05254_, _05230_, _03087_);
  and (_05255_, _05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or (_05841_, _05255_, _05254_);
  and (_05257_, _04990_, _03256_);
  and (_05258_, _05257_, _03060_);
  not (_05260_, _05257_);
  and (_05261_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or (_05844_, _05261_, _05258_);
  and (_05263_, _05257_, _03067_);
  and (_05264_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or (_05848_, _05264_, _05263_);
  and (_05266_, _05257_, _03071_);
  and (_05267_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or (_05851_, _05267_, _05266_);
  and (_05269_, _05257_, _03074_);
  and (_05270_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or (_05854_, _05270_, _05269_);
  and (_05272_, _05257_, _03077_);
  and (_05273_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or (_05857_, _05273_, _05272_);
  and (_05275_, _05257_, _03080_);
  and (_05276_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or (_05860_, _05276_, _05275_);
  and (_05278_, _05257_, _03083_);
  and (_05279_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or (_05863_, _05279_, _05278_);
  and (_05281_, _05257_, _03087_);
  and (_05282_, _05260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or (_05866_, _05282_, _05281_);
  and (_05284_, _04990_, _03275_);
  and (_05285_, _05284_, _03060_);
  not (_05286_, _05284_);
  and (_05288_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_05869_, _05288_, _05285_);
  and (_05289_, _05284_, _03067_);
  and (_05291_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_05872_, _05291_, _05289_);
  and (_05292_, _05284_, _03071_);
  and (_05294_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_05876_, _05294_, _05292_);
  and (_05295_, _05284_, _03074_);
  and (_05297_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_05879_, _05297_, _05295_);
  and (_05299_, _05284_, _03077_);
  and (_05300_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_05882_, _05300_, _05299_);
  and (_05301_, _05284_, _03080_);
  and (_05303_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_05885_, _05303_, _05301_);
  and (_05304_, _05284_, _03083_);
  and (_05306_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_05888_, _05306_, _05304_);
  and (_05307_, _05284_, _03087_);
  and (_05309_, _05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_05890_, _05309_, _05307_);
  and (_05310_, _04990_, _03295_);
  and (_05312_, _05310_, _03060_);
  not (_05313_, _05310_);
  and (_05314_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_05894_, _05314_, _05312_);
  and (_05316_, _05310_, _03067_);
  and (_05317_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_05897_, _05317_, _05316_);
  and (_05319_, _05310_, _03071_);
  and (_05320_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_05900_, _05320_, _05319_);
  and (_05322_, _05310_, _03074_);
  and (_05324_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_05904_, _05324_, _05322_);
  and (_05325_, _05310_, _03077_);
  and (_05326_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_05907_, _05326_, _05325_);
  and (_05328_, _05310_, _03080_);
  and (_05329_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_05910_, _05329_, _05328_);
  and (_05331_, _05310_, _03083_);
  and (_05332_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_05913_, _05332_, _05331_);
  and (_05334_, _05310_, _03087_);
  and (_05335_, _05313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_05915_, _05335_, _05334_);
  and (_05337_, _04990_, _03315_);
  and (_05338_, _05337_, _03060_);
  not (_05340_, _05337_);
  and (_05341_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or (_05919_, _05341_, _05338_);
  and (_05343_, _05337_, _03067_);
  and (_05344_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or (_05922_, _05344_, _05343_);
  and (_05346_, _05337_, _03071_);
  and (_05347_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or (_05925_, _05347_, _05346_);
  and (_05349_, _05337_, _03074_);
  and (_05350_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or (_05928_, _05350_, _05349_);
  and (_05352_, _05337_, _03077_);
  and (_05353_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or (_05931_, _05353_, _05352_);
  and (_05355_, _05337_, _03080_);
  and (_05356_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_05934_, _05356_, _05355_);
  and (_05358_, _05337_, _03083_);
  and (_05359_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or (_05937_, _05359_, _05358_);
  and (_05361_, _05337_, _03087_);
  and (_05362_, _05340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or (_05940_, _05362_, _05361_);
  and (_05364_, _04990_, _03334_);
  and (_05365_, _05364_, _03060_);
  not (_05366_, _05364_);
  and (_05368_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or (_05943_, _05368_, _05365_);
  and (_05369_, _05364_, _03067_);
  and (_05371_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or (_05946_, _05371_, _05369_);
  and (_05373_, _05364_, _03071_);
  and (_05374_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or (_05949_, _05374_, _05373_);
  and (_05375_, _05364_, _03074_);
  and (_05377_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or (_05952_, _05377_, _05375_);
  and (_05378_, _05364_, _03077_);
  and (_05380_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or (_05956_, _05380_, _05378_);
  and (_05381_, _05364_, _03080_);
  and (_05383_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or (_05959_, _05383_, _05381_);
  and (_05384_, _05364_, _03083_);
  and (_05386_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or (_05962_, _05386_, _05384_);
  and (_05387_, _05364_, _03087_);
  and (_05389_, _05366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_05964_, _05389_, _05387_);
  and (_05390_, _04990_, _03353_);
  and (_05392_, _05390_, _03060_);
  not (_05393_, _05390_);
  and (_05394_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_05968_, _05394_, _05392_);
  and (_05396_, _05390_, _03067_);
  and (_05398_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_05971_, _05398_, _05396_);
  and (_05399_, _05390_, _03071_);
  and (_05400_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_05974_, _05400_, _05399_);
  and (_05402_, _05390_, _03074_);
  and (_05403_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_05977_, _05403_, _05402_);
  and (_05405_, _05390_, _03077_);
  and (_05406_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_05980_, _05406_, _05405_);
  and (_05408_, _05390_, _03080_);
  and (_05409_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_05984_, _05409_, _05408_);
  and (_05411_, _05390_, _03083_);
  and (_05412_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_05987_, _05412_, _05411_);
  and (_05414_, _05390_, _03087_);
  and (_05415_, _05393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_05989_, _05415_, _05414_);
  and (_05417_, _04558_, _03699_);
  and (_05418_, _05417_, _02963_);
  and (_05420_, _05418_, _03060_);
  not (_05421_, _05418_);
  and (_05423_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_05993_, _05423_, _05420_);
  and (_05424_, _05418_, _03067_);
  and (_05425_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_05996_, _05425_, _05424_);
  and (_05427_, _05418_, _03071_);
  and (_05428_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_05999_, _05428_, _05427_);
  and (_05430_, _05418_, _03074_);
  and (_05431_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_06002_, _05431_, _05430_);
  and (_05433_, _05418_, _03077_);
  and (_05434_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_06005_, _05434_, _05433_);
  and (_05436_, _05418_, _03080_);
  and (_05437_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_06009_, _05437_, _05436_);
  and (_05439_, _05418_, _03083_);
  and (_05440_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_06012_, _05440_, _05439_);
  and (_05442_, _05418_, _03087_);
  and (_05443_, _05421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_06014_, _05443_, _05442_);
  and (_05445_, _05417_, _03062_);
  and (_05447_, _05445_, _03060_);
  not (_05448_, _05445_);
  and (_05449_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or (_06018_, _05449_, _05447_);
  and (_05451_, _05445_, _03067_);
  and (_05452_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or (_06021_, _05452_, _05451_);
  and (_05454_, _05445_, _03071_);
  and (_05455_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or (_06024_, _05455_, _05454_);
  and (_05457_, _05445_, _03074_);
  and (_05458_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or (_06027_, _05458_, _05457_);
  and (_05460_, _05445_, _03077_);
  and (_05461_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or (_06030_, _05461_, _05460_);
  and (_05463_, _05445_, _03080_);
  and (_05464_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or (_06033_, _05464_, _05463_);
  and (_05466_, _05445_, _03083_);
  and (_05467_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or (_06037_, _05467_, _05466_);
  and (_05469_, _05445_, _03087_);
  and (_05470_, _05448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_06039_, _05470_, _05469_);
  and (_05472_, _05417_, _03091_);
  and (_05473_, _05472_, _03060_);
  not (_05474_, _05472_);
  and (_05476_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or (_06043_, _05476_, _05473_);
  and (_05477_, _05472_, _03067_);
  and (_05479_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or (_06046_, _05479_, _05477_);
  and (_05480_, _05472_, _03071_);
  and (_05482_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or (_06049_, _05482_, _05480_);
  and (_05483_, _05472_, _03074_);
  and (_05485_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or (_06052_, _05485_, _05483_);
  and (_05486_, _05472_, _03077_);
  and (_05488_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or (_06055_, _05488_, _05486_);
  and (_05489_, _05472_, _03080_);
  and (_05491_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or (_06058_, _05491_, _05489_);
  and (_05492_, _05472_, _03083_);
  and (_05494_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or (_06061_, _05494_, _05492_);
  and (_05496_, _05472_, _03087_);
  and (_05497_, _05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or (_06064_, _05497_, _05496_);
  and (_05498_, _05417_, _03113_);
  and (_05500_, _05498_, _03060_);
  not (_05501_, _05498_);
  and (_05502_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_06067_, _05502_, _05500_);
  and (_05504_, _05498_, _03067_);
  and (_05505_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_06070_, _05505_, _05504_);
  and (_05507_, _05498_, _03071_);
  and (_05508_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_06073_, _05508_, _05507_);
  and (_05510_, _05498_, _03074_);
  and (_05511_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_06076_, _05511_, _05510_);
  and (_05513_, _05498_, _03077_);
  and (_05514_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_06079_, _05514_, _05513_);
  and (_05516_, _05498_, _03080_);
  and (_05517_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_06082_, _05517_, _05516_);
  and (_05519_, _05498_, _03083_);
  and (_05521_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_06085_, _05521_, _05519_);
  and (_05522_, _05498_, _03087_);
  and (_05523_, _05501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_06088_, _05523_, _05522_);
  and (_05525_, _05417_, _03136_);
  and (_05526_, _05525_, _03060_);
  not (_05528_, _05525_);
  and (_05529_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_06092_, _05529_, _05526_);
  and (_05531_, _05525_, _03067_);
  and (_05532_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_06095_, _05532_, _05531_);
  and (_05534_, _05525_, _03071_);
  and (_05535_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_06098_, _05535_, _05534_);
  and (_05537_, _05525_, _03074_);
  and (_05538_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_06101_, _05538_, _05537_);
  and (_05540_, _05525_, _03077_);
  and (_05541_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_06104_, _05541_, _05540_);
  and (_05543_, _05525_, _03080_);
  and (_05544_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_06107_, _05544_, _05543_);
  and (_05546_, _05525_, _03083_);
  and (_05547_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_06110_, _05547_, _05546_);
  and (_05549_, _05525_, _03087_);
  and (_05550_, _05528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_06112_, _05550_, _05549_);
  and (_05552_, _05417_, _03159_);
  and (_05553_, _05552_, _03060_);
  not (_05554_, _05552_);
  and (_05556_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or (_06117_, _05556_, _05553_);
  and (_05557_, _05552_, _03067_);
  and (_05559_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or (_06120_, _05559_, _05557_);
  and (_05560_, _05552_, _03071_);
  and (_05562_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or (_06123_, _05562_, _05560_);
  and (_05563_, _05552_, _03074_);
  and (_05565_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or (_06126_, _05565_, _05563_);
  and (_05566_, _05552_, _03077_);
  and (_05568_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or (_06129_, _05568_, _05566_);
  and (_05570_, _05552_, _03080_);
  and (_05571_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or (_06132_, _05571_, _05570_);
  and (_05572_, _05552_, _03083_);
  and (_05574_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or (_06135_, _05574_, _05572_);
  and (_05575_, _05552_, _03087_);
  and (_05577_, _05554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_06137_, _05577_, _05575_);
  and (_05578_, _05417_, _03179_);
  and (_05580_, _05578_, _03060_);
  not (_05581_, _05578_);
  and (_05582_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or (_06141_, _05582_, _05580_);
  and (_05584_, _05578_, _03067_);
  and (_05585_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or (_06144_, _05585_, _05584_);
  and (_05587_, _05578_, _03071_);
  and (_05588_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or (_06147_, _05588_, _05587_);
  and (_05590_, _05578_, _03074_);
  and (_05591_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or (_06150_, _05591_, _05590_);
  and (_05593_, _05578_, _03077_);
  and (_05595_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or (_06153_, _05595_, _05593_);
  and (_05596_, _05578_, _03080_);
  and (_05597_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or (_06156_, _05597_, _05596_);
  and (_05599_, _05578_, _03083_);
  and (_05600_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or (_06159_, _05600_, _05599_);
  and (_05602_, _05578_, _03087_);
  and (_05603_, _05581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or (_06162_, _05603_, _05602_);
  and (_05605_, _05417_, _03198_);
  and (_05606_, _05605_, _03060_);
  not (_05607_, _05605_);
  and (_05609_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_06165_, _05609_, _05606_);
  and (_05610_, _05605_, _03067_);
  and (_05612_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_06169_, _05612_, _05610_);
  and (_05613_, _05605_, _03071_);
  and (_05615_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_06172_, _05615_, _05613_);
  and (_05616_, _05605_, _03074_);
  and (_05618_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_06175_, _05618_, _05616_);
  and (_05620_, _05605_, _03077_);
  and (_05621_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_06178_, _05621_, _05620_);
  and (_05622_, _05605_, _03080_);
  and (_05624_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_06181_, _05624_, _05622_);
  and (_05625_, _05605_, _03083_);
  and (_05627_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_06184_, _05627_, _05625_);
  and (_05628_, _05605_, _03087_);
  and (_05630_, _05607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_06186_, _05630_, _05628_);
  and (_05631_, _05417_, _03218_);
  and (_05633_, _05631_, _03060_);
  not (_05634_, _05631_);
  and (_05635_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or (_06190_, _05635_, _05633_);
  and (_05637_, _05631_, _03067_);
  and (_05638_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or (_06193_, _05638_, _05637_);
  and (_05640_, _05631_, _03071_);
  and (_05641_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or (_06197_, _05641_, _05640_);
  and (_05643_, _05631_, _03074_);
  and (_05645_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or (_06200_, _05645_, _05643_);
  and (_05646_, _05631_, _03077_);
  and (_05647_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or (_06203_, _05647_, _05646_);
  and (_05649_, _05631_, _03080_);
  and (_05650_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or (_06206_, _05650_, _05649_);
  and (_05652_, _05631_, _03083_);
  and (_05653_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or (_06209_, _05653_, _05652_);
  and (_05655_, _05631_, _03087_);
  and (_05656_, _05634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_06211_, _05656_, _05655_);
  and (_05658_, _05417_, _03237_);
  and (_05659_, _05658_, _03060_);
  not (_05661_, _05658_);
  and (_05662_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_06215_, _05662_, _05659_);
  and (_05664_, _05658_, _03067_);
  and (_05665_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_06218_, _05665_, _05664_);
  and (_05667_, _05658_, _03071_);
  and (_05668_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_06221_, _05668_, _05667_);
  and (_05670_, _05658_, _03074_);
  and (_05671_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_06224_, _05671_, _05670_);
  and (_05673_, _05658_, _03077_);
  and (_05674_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_06227_, _05674_, _05673_);
  and (_05676_, _05658_, _03080_);
  and (_05677_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_06230_, _05677_, _05676_);
  and (_05679_, _05658_, _03083_);
  and (_05680_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_06233_, _05680_, _05679_);
  and (_05682_, _05658_, _03087_);
  and (_05683_, _05661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_06236_, _05683_, _05682_);
  and (_05685_, _05417_, _03256_);
  and (_05686_, _05685_, _03060_);
  not (_05687_, _05685_);
  and (_05689_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_06239_, _05689_, _05686_);
  and (_05690_, _05685_, _03067_);
  and (_05692_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_06242_, _05692_, _05690_);
  and (_05694_, _05685_, _03071_);
  and (_05695_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_06245_, _05695_, _05694_);
  and (_05696_, _05685_, _03074_);
  and (_05698_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_06249_, _05698_, _05696_);
  and (_05699_, _05685_, _03077_);
  and (_05701_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_06252_, _05701_, _05699_);
  and (_05702_, _05685_, _03080_);
  and (_05704_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_06255_, _05704_, _05702_);
  and (_05705_, _05685_, _03083_);
  and (_05707_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_06258_, _05707_, _05705_);
  and (_05708_, _05685_, _03087_);
  and (_05710_, _05687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_06260_, _05710_, _05708_);
  and (_05711_, _05417_, _03275_);
  and (_05713_, _05711_, _03060_);
  not (_05714_, _05711_);
  and (_05715_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or (_06264_, _05715_, _05713_);
  and (_05717_, _05711_, _03067_);
  and (_05719_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or (_06267_, _05719_, _05717_);
  and (_05720_, _05711_, _03071_);
  and (_05721_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or (_06270_, _05721_, _05720_);
  and (_05723_, _05711_, _03074_);
  and (_05724_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or (_06273_, _05724_, _05723_);
  and (_05726_, _05711_, _03077_);
  and (_05727_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or (_06277_, _05727_, _05726_);
  and (_05729_, _05711_, _03080_);
  and (_05730_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or (_06280_, _05730_, _05729_);
  and (_05732_, _05711_, _03083_);
  and (_05733_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or (_06283_, _05733_, _05732_);
  and (_05735_, _05711_, _03087_);
  and (_05736_, _05714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or (_06286_, _05736_, _05735_);
  and (_05738_, _05417_, _03295_);
  and (_05739_, _05738_, _03060_);
  not (_05741_, _05738_);
  and (_05742_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or (_06289_, _05742_, _05739_);
  and (_05744_, _05738_, _03067_);
  and (_05745_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or (_06292_, _05745_, _05744_);
  and (_05747_, _05738_, _03071_);
  and (_05748_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or (_06295_, _05748_, _05747_);
  and (_05750_, _05738_, _03074_);
  and (_05751_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or (_06298_, _05751_, _05750_);
  and (_05753_, _05738_, _03077_);
  and (_05754_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or (_06301_, _05754_, _05753_);
  and (_05756_, _05738_, _03080_);
  and (_05757_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_06305_, _05757_, _05756_);
  and (_05759_, _05738_, _03083_);
  and (_05760_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or (_06308_, _05760_, _05759_);
  and (_05762_, _05738_, _03087_);
  and (_05763_, _05741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_06310_, _05763_, _05762_);
  and (_05765_, _05417_, _03315_);
  and (_05766_, _05765_, _03060_);
  not (_05768_, _05765_);
  and (_05769_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_06314_, _05769_, _05766_);
  and (_05770_, _05765_, _03067_);
  and (_05772_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_06317_, _05772_, _05770_);
  and (_05773_, _05765_, _03071_);
  and (_05775_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_06320_, _05775_, _05773_);
  and (_05776_, _05765_, _03074_);
  and (_05778_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_06323_, _05778_, _05776_);
  and (_05779_, _05765_, _03077_);
  and (_05781_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_06326_, _05781_, _05779_);
  and (_05782_, _05765_, _03080_);
  and (_05784_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_06329_, _05784_, _05782_);
  and (_05785_, _05765_, _03083_);
  and (_05787_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_06333_, _05787_, _05785_);
  and (_05788_, _05765_, _03087_);
  and (_05790_, _05768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_06335_, _05790_, _05788_);
  and (_05792_, _05417_, _03334_);
  and (_05793_, _05792_, _03060_);
  not (_05794_, _05792_);
  and (_05795_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_06339_, _05795_, _05793_);
  and (_05797_, _05792_, _03067_);
  and (_05798_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_06342_, _05798_, _05797_);
  and (_05800_, _05792_, _03071_);
  and (_05801_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_06345_, _05801_, _05800_);
  and (_05803_, _05792_, _03074_);
  and (_05804_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_06348_, _05804_, _05803_);
  and (_05806_, _05792_, _03077_);
  and (_05807_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_06351_, _05807_, _05806_);
  and (_05809_, _05792_, _03080_);
  and (_05810_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_06354_, _05810_, _05809_);
  and (_05812_, _05792_, _03083_);
  and (_05813_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_06357_, _05813_, _05812_);
  and (_05815_, _05792_, _03087_);
  and (_05817_, _05794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_06360_, _05817_, _05815_);
  and (_05818_, _05417_, _03353_);
  and (_05819_, _05818_, _03060_);
  not (_05821_, _05818_);
  and (_05822_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or (_06363_, _05822_, _05819_);
  and (_05824_, _05818_, _03067_);
  and (_05825_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or (_06366_, _05825_, _05824_);
  and (_05827_, _05818_, _03071_);
  and (_05828_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or (_06369_, _05828_, _05827_);
  and (_05830_, _05818_, _03074_);
  and (_05831_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or (_06372_, _05831_, _05830_);
  and (_05833_, _05818_, _03077_);
  and (_05834_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or (_06375_, _05834_, _05833_);
  and (_05836_, _05818_, _03080_);
  and (_05837_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or (_06378_, _05837_, _05836_);
  and (_05839_, _05818_, _03083_);
  and (_05840_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or (_06381_, _05840_, _05839_);
  and (_05842_, _05818_, _03087_);
  and (_05843_, _05821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or (_06384_, _05843_, _05842_);
  and (_05845_, _04558_, _04125_);
  and (_05846_, _05845_, _02963_);
  and (_05847_, _05846_, _03060_);
  not (_05849_, _05846_);
  and (_05850_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or (_06389_, _05850_, _05847_);
  and (_05852_, _05846_, _03067_);
  and (_05853_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or (_06392_, _05853_, _05852_);
  and (_05855_, _05846_, _03071_);
  and (_05856_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or (_06395_, _05856_, _05855_);
  and (_05858_, _05846_, _03074_);
  and (_05859_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or (_06398_, _05859_, _05858_);
  and (_05861_, _05846_, _03077_);
  and (_05862_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or (_06401_, _05862_, _05861_);
  and (_05864_, _05846_, _03080_);
  and (_05865_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or (_06404_, _05865_, _05864_);
  and (_05867_, _05846_, _03083_);
  and (_05868_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or (_06407_, _05868_, _05867_);
  and (_05870_, _05846_, _03087_);
  and (_05871_, _05849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or (_06409_, _05871_, _05870_);
  and (_05873_, _05845_, _03062_);
  and (_05874_, _05873_, _03060_);
  not (_05875_, _05873_);
  and (_05877_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_06413_, _05877_, _05874_);
  and (_05878_, _05873_, _03067_);
  and (_05880_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_06416_, _05880_, _05878_);
  and (_05881_, _05873_, _03071_);
  and (_05883_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_06419_, _05883_, _05881_);
  and (_05884_, _05873_, _03074_);
  and (_05886_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_06422_, _05886_, _05884_);
  and (_05887_, _05873_, _03077_);
  and (_05889_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_06425_, _05889_, _05887_);
  and (_05891_, _05873_, _03080_);
  and (_05892_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_06428_, _05892_, _05891_);
  and (_05893_, _05873_, _03083_);
  and (_05895_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_06431_, _05895_, _05893_);
  and (_05896_, _05873_, _03087_);
  and (_05898_, _05875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_06434_, _05898_, _05896_);
  and (_05899_, _05845_, _03091_);
  and (_05901_, _05899_, _03060_);
  not (_05902_, _05899_);
  and (_05903_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_06438_, _05903_, _05901_);
  and (_05905_, _05899_, _03067_);
  and (_05906_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_06441_, _05906_, _05905_);
  and (_05908_, _05899_, _03071_);
  and (_05909_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_06444_, _05909_, _05908_);
  and (_05911_, _05899_, _03074_);
  and (_05912_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_06447_, _05912_, _05911_);
  and (_05914_, _05899_, _03077_);
  and (_05916_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_06450_, _05916_, _05914_);
  and (_05917_, _05899_, _03080_);
  and (_05918_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_06453_, _05918_, _05917_);
  and (_05920_, _05899_, _03083_);
  and (_05921_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_06456_, _05921_, _05920_);
  and (_05923_, _05899_, _03087_);
  and (_05924_, _05902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_06458_, _05924_, _05923_);
  and (_05926_, _05845_, _03113_);
  and (_05927_, _05926_, _03060_);
  not (_05929_, _05926_);
  and (_05930_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or (_06462_, _05930_, _05927_);
  and (_05932_, _05926_, _03067_);
  and (_05933_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or (_06466_, _05933_, _05932_);
  and (_05935_, _05926_, _03071_);
  and (_05936_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or (_06469_, _05936_, _05935_);
  and (_05938_, _05926_, _03074_);
  and (_05939_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or (_06472_, _05939_, _05938_);
  and (_05941_, _05926_, _03077_);
  and (_05942_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or (_06475_, _05942_, _05941_);
  and (_05944_, _05926_, _03080_);
  and (_05945_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or (_06478_, _05945_, _05944_);
  and (_05947_, _05926_, _03083_);
  and (_05948_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or (_06481_, _05948_, _05947_);
  and (_05950_, _05926_, _03087_);
  and (_05951_, _05929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or (_06483_, _05951_, _05950_);
  and (_05953_, _05845_, _03136_);
  and (_05954_, _05953_, _03060_);
  not (_05955_, _05953_);
  and (_05957_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or (_06487_, _05957_, _05954_);
  and (_05958_, _05953_, _03067_);
  and (_05960_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or (_06490_, _05960_, _05958_);
  and (_05961_, _05953_, _03071_);
  and (_05963_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or (_06493_, _05963_, _05961_);
  and (_05965_, _05953_, _03074_);
  and (_05966_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or (_06496_, _05966_, _05965_);
  and (_05967_, _05953_, _03077_);
  and (_05969_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or (_06499_, _05969_, _05967_);
  and (_05970_, _05953_, _03080_);
  and (_05972_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or (_06502_, _05972_, _05970_);
  and (_05973_, _05953_, _03083_);
  and (_05975_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or (_06505_, _05975_, _05973_);
  and (_05976_, _05953_, _03087_);
  and (_05978_, _05955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or (_06508_, _05978_, _05976_);
  and (_05979_, _05845_, _03159_);
  and (_05981_, _05979_, _03060_);
  not (_05982_, _05979_);
  and (_05983_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_06511_, _05983_, _05981_);
  and (_05985_, _05979_, _03067_);
  and (_05986_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_06514_, _05986_, _05985_);
  and (_05988_, _05979_, _03071_);
  and (_05990_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_06518_, _05990_, _05988_);
  and (_05991_, _05979_, _03074_);
  and (_05992_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_06521_, _05992_, _05991_);
  and (_05994_, _05979_, _03077_);
  and (_05995_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_06525_, _05995_, _05994_);
  and (_05997_, _05979_, _03080_);
  and (_05998_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_06528_, _05998_, _05997_);
  and (_06000_, _05979_, _03083_);
  and (_06001_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_06531_, _06001_, _06000_);
  and (_06003_, _05979_, _03087_);
  and (_06004_, _05982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_06533_, _06004_, _06003_);
  and (_06006_, _05845_, _03179_);
  and (_06007_, _06006_, _03060_);
  not (_06008_, _06006_);
  and (_06010_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_06537_, _06010_, _06007_);
  and (_06011_, _06006_, _03067_);
  and (_06013_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_06540_, _06013_, _06011_);
  and (_06015_, _06006_, _03071_);
  and (_06016_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_06543_, _06016_, _06015_);
  and (_06017_, _06006_, _03074_);
  and (_06019_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_06547_, _06019_, _06017_);
  and (_06020_, _06006_, _03077_);
  and (_06022_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_06550_, _06022_, _06020_);
  and (_06023_, _06006_, _03080_);
  and (_06025_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_06553_, _06025_, _06023_);
  and (_06026_, _06006_, _03083_);
  and (_06028_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_06556_, _06028_, _06026_);
  and (_06029_, _06006_, _03087_);
  and (_06031_, _06008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_06558_, _06031_, _06029_);
  and (_06032_, _05845_, _03198_);
  and (_06034_, _06032_, _03060_);
  not (_06035_, _06032_);
  and (_06036_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or (_06562_, _06036_, _06034_);
  and (_06038_, _06032_, _03067_);
  and (_06040_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or (_06565_, _06040_, _06038_);
  and (_06041_, _06032_, _03071_);
  and (_06042_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or (_06568_, _06042_, _06041_);
  and (_06044_, _06032_, _03074_);
  and (_06045_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or (_06571_, _06045_, _06044_);
  and (_06047_, _06032_, _03077_);
  and (_06048_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or (_06574_, _06048_, _06047_);
  and (_06050_, _06032_, _03080_);
  and (_06051_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or (_06577_, _06051_, _06050_);
  and (_06053_, _06032_, _03083_);
  and (_06054_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or (_06580_, _06054_, _06053_);
  and (_06056_, _06032_, _03087_);
  and (_06057_, _06035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or (_06583_, _06057_, _06056_);
  and (_06059_, _05845_, _03218_);
  and (_06060_, _06059_, _03060_);
  not (_06062_, _06059_);
  and (_06063_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_06586_, _06063_, _06060_);
  and (_06065_, _06059_, _03067_);
  and (_06066_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_06589_, _06066_, _06065_);
  and (_06068_, _06059_, _03071_);
  and (_06069_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_06592_, _06069_, _06068_);
  and (_06071_, _06059_, _03074_);
  and (_06072_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_06595_, _06072_, _06071_);
  and (_06074_, _06059_, _03077_);
  and (_06075_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_06599_, _06075_, _06074_);
  and (_06077_, _06059_, _03080_);
  and (_06078_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_06602_, _06078_, _06077_);
  and (_06080_, _06059_, _03083_);
  and (_06081_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_06605_, _06081_, _06080_);
  and (_06083_, _06059_, _03087_);
  and (_06084_, _06062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_06607_, _06084_, _06083_);
  and (_06086_, _05845_, _03237_);
  and (_06087_, _06086_, _03060_);
  not (_06089_, _06086_);
  and (_06090_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or (_06611_, _06090_, _06087_);
  and (_06091_, _06086_, _03067_);
  and (_06093_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or (_06614_, _06093_, _06091_);
  and (_06094_, _06086_, _03071_);
  and (_06096_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or (_06617_, _06096_, _06094_);
  and (_06097_, _06086_, _03074_);
  and (_06099_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or (_06620_, _06099_, _06097_);
  and (_06100_, _06086_, _03077_);
  and (_06102_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or (_06623_, _06102_, _06100_);
  and (_06103_, _06086_, _03080_);
  and (_06105_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or (_06627_, _06105_, _06103_);
  and (_06106_, _06086_, _03083_);
  and (_06108_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or (_06630_, _06108_, _06106_);
  and (_06109_, _06086_, _03087_);
  and (_06111_, _06089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or (_06632_, _06111_, _06109_);
  and (_06113_, _05845_, _03256_);
  and (_06114_, _06113_, _03060_);
  not (_06115_, _06113_);
  and (_06116_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or (_06636_, _06116_, _06114_);
  and (_06118_, _06113_, _03067_);
  and (_06119_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or (_06639_, _06119_, _06118_);
  and (_06121_, _06113_, _03071_);
  and (_06122_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or (_06642_, _06122_, _06121_);
  and (_06124_, _06113_, _03074_);
  and (_06125_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or (_06645_, _06125_, _06124_);
  and (_06127_, _06113_, _03077_);
  and (_06128_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or (_06648_, _06128_, _06127_);
  and (_06130_, _06113_, _03080_);
  and (_06131_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or (_06651_, _06131_, _06130_);
  and (_06133_, _06113_, _03083_);
  and (_06134_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or (_06654_, _06134_, _06133_);
  and (_06136_, _06113_, _03087_);
  and (_06138_, _06115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or (_06657_, _06138_, _06136_);
  and (_06139_, _05845_, _03275_);
  and (_06140_, _06139_, _03060_);
  not (_06142_, _06139_);
  and (_06143_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_06660_, _06143_, _06140_);
  and (_06145_, _06139_, _03067_);
  and (_06146_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_06663_, _06146_, _06145_);
  and (_06148_, _06139_, _03071_);
  and (_06149_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_06666_, _06149_, _06148_);
  and (_06151_, _06139_, _03074_);
  and (_06152_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_06669_, _06152_, _06151_);
  and (_06154_, _06139_, _03077_);
  and (_06155_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_06672_, _06155_, _06154_);
  and (_06157_, _06139_, _03080_);
  and (_06158_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_06675_, _06158_, _06157_);
  and (_06160_, _06139_, _03083_);
  and (_06161_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_06679_, _06161_, _06160_);
  and (_06163_, _06139_, _03087_);
  and (_06164_, _06142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_06681_, _06164_, _06163_);
  and (_06166_, _05845_, _03295_);
  and (_06167_, _06166_, _03060_);
  not (_06168_, _06166_);
  and (_06170_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_06685_, _06170_, _06167_);
  and (_06171_, _06166_, _03067_);
  and (_06173_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_06688_, _06173_, _06171_);
  and (_06174_, _06166_, _03071_);
  and (_06176_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_06691_, _06176_, _06174_);
  and (_06177_, _06166_, _03074_);
  and (_06179_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_06694_, _06179_, _06177_);
  and (_06180_, _06166_, _03077_);
  and (_06182_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_06697_, _06182_, _06180_);
  and (_06183_, _06166_, _03080_);
  and (_06185_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_06700_, _06185_, _06183_);
  and (_06187_, _06166_, _03083_);
  and (_06188_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_06703_, _06188_, _06187_);
  and (_06189_, _06166_, _03087_);
  and (_06191_, _06168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_06706_, _06191_, _06189_);
  and (_06192_, _05845_, _03315_);
  and (_06194_, _06192_, _03060_);
  not (_06195_, _06192_);
  and (_06196_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or (_06710_, _06196_, _06194_);
  and (_06198_, _06192_, _03067_);
  and (_06199_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or (_06713_, _06199_, _06198_);
  and (_06201_, _06192_, _03071_);
  and (_06202_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or (_06716_, _06202_, _06201_);
  and (_06204_, _06192_, _03074_);
  and (_06205_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or (_06719_, _06205_, _06204_);
  and (_06207_, _06192_, _03077_);
  and (_06208_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or (_06722_, _06208_, _06207_);
  and (_06210_, _06192_, _03080_);
  and (_06212_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or (_06725_, _06212_, _06210_);
  and (_06213_, _06192_, _03083_);
  and (_06214_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or (_06728_, _06214_, _06213_);
  and (_06216_, _06192_, _03087_);
  and (_06217_, _06195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or (_06730_, _06217_, _06216_);
  and (_06219_, _05845_, _03334_);
  and (_06220_, _06219_, _03060_);
  not (_06222_, _06219_);
  and (_06223_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or (_06735_, _06223_, _06220_);
  and (_06225_, _06219_, _03067_);
  and (_06226_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or (_06738_, _06226_, _06225_);
  and (_06228_, _06219_, _03071_);
  and (_06229_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or (_06741_, _06229_, _06228_);
  and (_06231_, _06219_, _03074_);
  and (_06232_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or (_06744_, _06232_, _06231_);
  and (_06234_, _06219_, _03077_);
  and (_06235_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or (_06747_, _06235_, _06234_);
  and (_06237_, _06219_, _03080_);
  and (_06238_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or (_06750_, _06238_, _06237_);
  and (_06240_, _06219_, _03083_);
  and (_06241_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or (_06753_, _06241_, _06240_);
  and (_06243_, _06219_, _03087_);
  and (_06244_, _06222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or (_06755_, _06244_, _06243_);
  and (_06246_, _05845_, _03353_);
  and (_06247_, _06246_, _03060_);
  not (_06248_, _06246_);
  and (_06250_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_06759_, _06250_, _06247_);
  and (_06251_, _06246_, _03067_);
  and (_06253_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_06762_, _06253_, _06251_);
  and (_06254_, _06246_, _03071_);
  and (_06256_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_06765_, _06256_, _06254_);
  and (_06257_, _06246_, _03074_);
  and (_06259_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_06768_, _06259_, _06257_);
  and (_06261_, _06246_, _03077_);
  and (_06262_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_06771_, _06262_, _06261_);
  and (_06263_, _06246_, _03080_);
  and (_06265_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_06774_, _06265_, _06263_);
  and (_06266_, _06246_, _03083_);
  and (_06268_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_06777_, _06268_, _06266_);
  and (_06269_, _06246_, _03087_);
  and (_06271_, _06248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_06780_, _06271_, _06269_);
  and (_06272_, _02137_, _26459_);
  and (_06274_, _06272_, _02966_);
  and (_06275_, _06274_, _02963_);
  and (_06276_, _06275_, _03060_);
  not (_06278_, _06275_);
  and (_06279_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_06787_, _06279_, _06276_);
  and (_06281_, _06275_, _03067_);
  and (_06282_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_06790_, _06282_, _06281_);
  and (_06284_, _06275_, _03071_);
  and (_06285_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_06793_, _06285_, _06284_);
  and (_06287_, _06275_, _03074_);
  and (_06288_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_06796_, _06288_, _06287_);
  and (_06290_, _06275_, _03077_);
  and (_06291_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_06799_, _06291_, _06290_);
  and (_06293_, _06275_, _03080_);
  and (_06294_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_06802_, _06294_, _06293_);
  and (_06296_, _06275_, _03083_);
  and (_06297_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_06805_, _06297_, _06296_);
  and (_06299_, _06275_, _03087_);
  and (_06300_, _06278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_06808_, _06300_, _06299_);
  and (_06302_, _06274_, _03062_);
  and (_06303_, _06302_, _03060_);
  not (_06304_, _06302_);
  and (_06306_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  or (_06812_, _06306_, _06303_);
  and (_06307_, _06302_, _03067_);
  and (_06309_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or (_06815_, _06309_, _06307_);
  and (_06311_, _06302_, _03071_);
  and (_06312_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or (_06818_, _06312_, _06311_);
  and (_06313_, _06302_, _03074_);
  and (_06315_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  or (_06821_, _06315_, _06313_);
  and (_06316_, _06302_, _03077_);
  and (_06318_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or (_06824_, _06318_, _06316_);
  and (_06319_, _06302_, _03080_);
  and (_06321_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or (_06827_, _06321_, _06319_);
  and (_06322_, _06302_, _03083_);
  and (_06324_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or (_06830_, _06324_, _06322_);
  and (_06325_, _06302_, _03087_);
  and (_06327_, _06304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or (_06832_, _06327_, _06325_);
  and (_06328_, _06274_, _03091_);
  and (_06330_, _06328_, _03060_);
  not (_06331_, _06328_);
  and (_06332_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or (_06836_, _06332_, _06330_);
  and (_06334_, _06328_, _03067_);
  and (_06336_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or (_06840_, _06336_, _06334_);
  and (_06337_, _06328_, _03071_);
  and (_06338_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or (_06843_, _06338_, _06337_);
  and (_06340_, _06328_, _03074_);
  and (_06341_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or (_06846_, _06341_, _06340_);
  and (_06343_, _06328_, _03077_);
  and (_06344_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or (_06849_, _06344_, _06343_);
  and (_06346_, _06328_, _03080_);
  and (_06347_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  or (_06852_, _06347_, _06346_);
  and (_06349_, _06328_, _03083_);
  and (_06350_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or (_06855_, _06350_, _06349_);
  and (_06352_, _06328_, _03087_);
  and (_06353_, _06331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or (_06857_, _06353_, _06352_);
  and (_06355_, _06274_, _03113_);
  and (_06356_, _06355_, _03060_);
  not (_06358_, _06355_);
  and (_06359_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_06861_, _06359_, _06356_);
  and (_06361_, _06355_, _03067_);
  and (_06362_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_06864_, _06362_, _06361_);
  and (_06364_, _06355_, _03071_);
  and (_06365_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_06867_, _06365_, _06364_);
  and (_06367_, _06355_, _03074_);
  and (_06368_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_06870_, _06368_, _06367_);
  and (_06370_, _06355_, _03077_);
  and (_06371_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_06873_, _06371_, _06370_);
  and (_06373_, _06355_, _03080_);
  and (_06374_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_06876_, _06374_, _06373_);
  and (_06376_, _06355_, _03083_);
  and (_06377_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_06879_, _06377_, _06376_);
  and (_06379_, _06355_, _03087_);
  and (_06380_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_06882_, _06380_, _06379_);
  and (_06382_, _06274_, _03136_);
  and (_06383_, _06382_, _03060_);
  not (_06385_, _06382_);
  and (_06386_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_06885_, _06386_, _06383_);
  and (_06387_, _06382_, _03067_);
  and (_06388_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_06888_, _06388_, _06387_);
  and (_06390_, _06382_, _03071_);
  and (_06391_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_06892_, _06391_, _06390_);
  and (_06393_, _06382_, _03074_);
  and (_06394_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_06895_, _06394_, _06393_);
  and (_06396_, _06382_, _03077_);
  and (_06397_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_06898_, _06397_, _06396_);
  and (_06399_, _06382_, _03080_);
  and (_06400_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_06901_, _06400_, _06399_);
  and (_06402_, _06382_, _03083_);
  and (_06403_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_06904_, _06403_, _06402_);
  and (_06405_, _06382_, _03087_);
  and (_06406_, _06385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_06906_, _06406_, _06405_);
  and (_06408_, _06274_, _03159_);
  and (_06410_, _06408_, _03060_);
  not (_06411_, _06408_);
  and (_06412_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  or (_06910_, _06412_, _06410_);
  and (_06414_, _06408_, _03067_);
  and (_06415_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or (_06913_, _06415_, _06414_);
  and (_06417_, _06408_, _03071_);
  and (_06418_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or (_06916_, _06418_, _06417_);
  and (_06420_, _06408_, _03074_);
  and (_06421_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or (_06920_, _06421_, _06420_);
  and (_06423_, _06408_, _03077_);
  and (_06424_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or (_06923_, _06424_, _06423_);
  and (_06426_, _06408_, _03080_);
  and (_06427_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or (_06926_, _06427_, _06426_);
  and (_06429_, _06408_, _03083_);
  and (_06430_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or (_06929_, _06430_, _06429_);
  and (_06432_, _06408_, _03087_);
  and (_06433_, _06411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or (_06931_, _06433_, _06432_);
  and (_06435_, _06274_, _03179_);
  and (_06436_, _06435_, _03060_);
  not (_06437_, _06435_);
  and (_06439_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or (_06935_, _06439_, _06436_);
  and (_06440_, _06435_, _03067_);
  and (_06442_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or (_06938_, _06442_, _06440_);
  and (_06443_, _06435_, _03071_);
  and (_06445_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or (_06941_, _06445_, _06443_);
  and (_06446_, _06435_, _03074_);
  and (_06448_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  or (_06944_, _06448_, _06446_);
  and (_06449_, _06435_, _03077_);
  and (_06451_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or (_06947_, _06451_, _06449_);
  and (_06452_, _06435_, _03080_);
  and (_06454_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  or (_06950_, _06454_, _06452_);
  and (_06455_, _06435_, _03083_);
  and (_06457_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or (_06953_, _06457_, _06455_);
  and (_06459_, _06435_, _03087_);
  and (_06460_, _06437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or (_06956_, _06460_, _06459_);
  and (_06461_, _06274_, _03198_);
  and (_06463_, _06461_, _03060_);
  not (_06464_, _06461_);
  and (_06465_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_06959_, _06465_, _06463_);
  and (_06467_, _06461_, _03067_);
  and (_06468_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_06962_, _06468_, _06467_);
  and (_06470_, _06461_, _03071_);
  and (_06471_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_06965_, _06471_, _06470_);
  and (_06473_, _06461_, _03074_);
  and (_06474_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_06968_, _06474_, _06473_);
  and (_06476_, _06461_, _03077_);
  and (_06477_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_06972_, _06477_, _06476_);
  and (_06479_, _06461_, _03080_);
  and (_06480_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_06975_, _06480_, _06479_);
  and (_06482_, _06461_, _03083_);
  and (_06484_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_06978_, _06484_, _06482_);
  and (_06485_, _06461_, _03087_);
  and (_06486_, _06464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_06980_, _06486_, _06485_);
  and (_06488_, _06274_, _03218_);
  and (_06489_, _06488_, _03060_);
  not (_06491_, _06488_);
  and (_06492_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  or (_06984_, _06492_, _06489_);
  and (_06494_, _06488_, _03067_);
  and (_06495_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or (_06987_, _06495_, _06494_);
  and (_06497_, _06488_, _03071_);
  and (_06498_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or (_06990_, _06498_, _06497_);
  and (_06500_, _06488_, _03074_);
  and (_06501_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  or (_06993_, _06501_, _06500_);
  and (_06503_, _06488_, _03077_);
  and (_06504_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or (_06996_, _06504_, _06503_);
  and (_06506_, _06488_, _03080_);
  and (_06507_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or (_07000_, _06507_, _06506_);
  and (_06509_, _06488_, _03083_);
  and (_06510_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or (_07003_, _06510_, _06509_);
  and (_06512_, _06488_, _03087_);
  and (_06513_, _06491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or (_07005_, _06513_, _06512_);
  and (_06515_, _06274_, _03237_);
  and (_06516_, _06515_, _03060_);
  not (_06517_, _06515_);
  and (_06519_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_07009_, _06519_, _06516_);
  and (_06520_, _06515_, _03067_);
  and (_06522_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_07012_, _06522_, _06520_);
  and (_06523_, _06515_, _03071_);
  and (_06526_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_07015_, _06526_, _06523_);
  and (_06527_, _06515_, _03074_);
  and (_06529_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_07018_, _06529_, _06527_);
  and (_06530_, _06515_, _03077_);
  and (_06532_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_07021_, _06532_, _06530_);
  and (_06534_, _06515_, _03080_);
  and (_06535_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_07024_, _06535_, _06534_);
  and (_06536_, _06515_, _03083_);
  and (_06538_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_07027_, _06538_, _06536_);
  and (_06539_, _06515_, _03087_);
  and (_06541_, _06517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_07030_, _06541_, _06539_);
  and (_06542_, _06274_, _03256_);
  and (_06544_, _06542_, _03060_);
  not (_06545_, _06542_);
  and (_06546_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_07033_, _06546_, _06544_);
  and (_06548_, _06542_, _03067_);
  and (_06549_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_07036_, _06549_, _06548_);
  and (_06551_, _06542_, _03071_);
  and (_06552_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_07039_, _06552_, _06551_);
  and (_06554_, _06542_, _03074_);
  and (_06555_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_07042_, _06555_, _06554_);
  and (_06557_, _06542_, _03077_);
  and (_06559_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_07045_, _06559_, _06557_);
  and (_06560_, _06542_, _03080_);
  and (_06561_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_07048_, _06561_, _06560_);
  and (_06563_, _06542_, _03083_);
  and (_06564_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_07052_, _06564_, _06563_);
  and (_06566_, _06542_, _03087_);
  and (_06567_, _06545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_07054_, _06567_, _06566_);
  and (_06569_, _06274_, _03275_);
  and (_06570_, _06569_, _03060_);
  not (_06572_, _06569_);
  and (_06573_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or (_07058_, _06573_, _06570_);
  and (_06575_, _06569_, _03067_);
  and (_06576_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or (_07061_, _06576_, _06575_);
  and (_06578_, _06569_, _03071_);
  and (_06579_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or (_07064_, _06579_, _06578_);
  and (_06581_, _06569_, _03074_);
  and (_06582_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  or (_07067_, _06582_, _06581_);
  and (_06584_, _06569_, _03077_);
  and (_06585_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or (_07070_, _06585_, _06584_);
  and (_06587_, _06569_, _03080_);
  and (_06588_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or (_07073_, _06588_, _06587_);
  and (_06590_, _06569_, _03083_);
  and (_06591_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or (_07076_, _06591_, _06590_);
  and (_06593_, _06569_, _03087_);
  and (_06594_, _06572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or (_07079_, _06594_, _06593_);
  and (_06596_, _06274_, _03295_);
  and (_06597_, _06596_, _03060_);
  not (_06598_, _06596_);
  and (_06600_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  or (_07083_, _06600_, _06597_);
  and (_06601_, _06596_, _03067_);
  and (_06603_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or (_07086_, _06603_, _06601_);
  and (_06604_, _06596_, _03071_);
  and (_06606_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or (_07089_, _06606_, _06604_);
  and (_06608_, _06596_, _03074_);
  and (_06609_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or (_07092_, _06609_, _06608_);
  and (_06610_, _06596_, _03077_);
  and (_06612_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or (_07095_, _06612_, _06610_);
  and (_06613_, _06596_, _03080_);
  and (_06615_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  or (_07098_, _06615_, _06613_);
  and (_06616_, _06596_, _03083_);
  and (_06618_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or (_07101_, _06618_, _06616_);
  and (_06619_, _06596_, _03087_);
  and (_06621_, _06598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or (_07103_, _06621_, _06619_);
  and (_06622_, _06274_, _03315_);
  and (_06624_, _06622_, _03060_);
  not (_06625_, _06622_);
  and (_06626_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_07107_, _06626_, _06624_);
  and (_06628_, _06622_, _03067_);
  and (_06629_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_07110_, _06629_, _06628_);
  and (_06631_, _06622_, _03071_);
  and (_06633_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_07113_, _06633_, _06631_);
  and (_06634_, _06622_, _03074_);
  and (_06635_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_07116_, _06635_, _06634_);
  and (_06637_, _06622_, _03077_);
  and (_06638_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_07119_, _06638_, _06637_);
  and (_06640_, _06622_, _03080_);
  and (_06641_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_07122_, _06641_, _06640_);
  and (_06643_, _06622_, _03083_);
  and (_06644_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_07125_, _06644_, _06643_);
  and (_06646_, _06622_, _03087_);
  and (_06647_, _06625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_07128_, _06647_, _06646_);
  and (_06649_, _06274_, _03334_);
  and (_06650_, _06649_, _03060_);
  not (_06652_, _06649_);
  and (_06653_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_07132_, _06653_, _06650_);
  and (_06655_, _06649_, _03067_);
  and (_06656_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_07135_, _06656_, _06655_);
  and (_06658_, _06649_, _03071_);
  and (_06659_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_07138_, _06659_, _06658_);
  and (_06661_, _06649_, _03074_);
  and (_06662_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_07141_, _06662_, _06661_);
  and (_06664_, _06649_, _03077_);
  and (_06665_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_07144_, _06665_, _06664_);
  and (_06667_, _06649_, _03080_);
  and (_06668_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_07147_, _06668_, _06667_);
  and (_06670_, _06649_, _03083_);
  and (_06671_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_07150_, _06671_, _06670_);
  and (_06673_, _06649_, _03087_);
  and (_06674_, _06652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_07153_, _06674_, _06673_);
  and (_06676_, _06274_, _03353_);
  and (_06677_, _06676_, _03060_);
  not (_06678_, _06676_);
  and (_06680_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  or (_07156_, _06680_, _06677_);
  and (_06682_, _06676_, _03067_);
  and (_06683_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or (_07160_, _06683_, _06682_);
  and (_06684_, _06676_, _03071_);
  and (_06686_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or (_07163_, _06686_, _06684_);
  and (_06687_, _06676_, _03074_);
  and (_06689_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or (_07166_, _06689_, _06687_);
  and (_06690_, _06676_, _03077_);
  and (_06692_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or (_07169_, _06692_, _06690_);
  and (_06693_, _06676_, _03080_);
  and (_06695_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  or (_07172_, _06695_, _06693_);
  and (_06696_, _06676_, _03083_);
  and (_06698_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or (_07175_, _06698_, _06696_);
  and (_06699_, _06676_, _03087_);
  and (_06701_, _06678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or (_07177_, _06701_, _06699_);
  and (_06702_, _03373_, _26459_);
  and (_06704_, _06702_, _02963_);
  and (_06705_, _06704_, _03060_);
  not (_06707_, _06704_);
  and (_06708_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or (_07182_, _06708_, _06705_);
  and (_06709_, _06704_, _03067_);
  and (_06711_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  or (_07185_, _06711_, _06709_);
  and (_06712_, _06704_, _03071_);
  and (_06714_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  or (_07188_, _06714_, _06712_);
  and (_06715_, _06704_, _03074_);
  and (_06717_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  or (_07191_, _06717_, _06715_);
  and (_06718_, _06704_, _03077_);
  and (_06720_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  or (_07194_, _06720_, _06718_);
  and (_06721_, _06704_, _03080_);
  and (_06723_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or (_07197_, _06723_, _06721_);
  and (_06724_, _06704_, _03083_);
  and (_06726_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  or (_07200_, _06726_, _06724_);
  and (_06727_, _06704_, _03087_);
  and (_06729_, _06707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or (_07203_, _06729_, _06727_);
  and (_06731_, _06702_, _03062_);
  and (_06732_, _06731_, _03060_);
  not (_06733_, _06731_);
  and (_06734_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_07206_, _06734_, _06732_);
  and (_06736_, _06731_, _03067_);
  and (_06737_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_07209_, _06737_, _06736_);
  and (_06739_, _06731_, _03071_);
  and (_06740_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_07213_, _06740_, _06739_);
  and (_06742_, _06731_, _03074_);
  and (_06743_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_07216_, _06743_, _06742_);
  and (_06745_, _06731_, _03077_);
  and (_06746_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_07219_, _06746_, _06745_);
  and (_06748_, _06731_, _03080_);
  and (_06749_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_07222_, _06749_, _06748_);
  and (_06751_, _06731_, _03083_);
  and (_06752_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_07225_, _06752_, _06751_);
  and (_06754_, _06731_, _03087_);
  and (_06756_, _06733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_07227_, _06756_, _06754_);
  and (_06757_, _06702_, _03091_);
  and (_06758_, _06757_, _03060_);
  not (_06760_, _06757_);
  and (_06761_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_07231_, _06761_, _06758_);
  and (_06763_, _06757_, _03067_);
  and (_06764_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_07234_, _06764_, _06763_);
  and (_06766_, _06757_, _03071_);
  and (_06767_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_07237_, _06767_, _06766_);
  and (_06769_, _06757_, _03074_);
  and (_06770_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_07241_, _06770_, _06769_);
  and (_06772_, _06757_, _03077_);
  and (_06773_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_07244_, _06773_, _06772_);
  and (_06775_, _06757_, _03080_);
  and (_06776_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_07247_, _06776_, _06775_);
  and (_06778_, _06757_, _03083_);
  and (_06779_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_07250_, _06779_, _06778_);
  and (_06781_, _06757_, _03087_);
  and (_06782_, _06760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_07252_, _06782_, _06781_);
  and (_06783_, _06702_, _03113_);
  and (_06784_, _06783_, _03060_);
  not (_06785_, _06783_);
  and (_06786_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or (_07256_, _06786_, _06784_);
  and (_06788_, _06783_, _03067_);
  and (_06789_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  or (_07259_, _06789_, _06788_);
  and (_06791_, _06783_, _03071_);
  and (_06792_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  or (_07262_, _06792_, _06791_);
  and (_06794_, _06783_, _03074_);
  and (_06795_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  or (_07265_, _06795_, _06794_);
  and (_06797_, _06783_, _03077_);
  and (_06798_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or (_07268_, _06798_, _06797_);
  and (_06800_, _06783_, _03080_);
  and (_06801_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or (_07271_, _06801_, _06800_);
  and (_06803_, _06783_, _03083_);
  and (_06804_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or (_07274_, _06804_, _06803_);
  and (_06806_, _06783_, _03087_);
  and (_06807_, _06785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  or (_07277_, _06807_, _06806_);
  and (_06809_, _06702_, _03136_);
  and (_06810_, _06809_, _03060_);
  not (_06811_, _06809_);
  and (_06813_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  or (_07280_, _06813_, _06810_);
  and (_06814_, _06809_, _03067_);
  and (_06816_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or (_07283_, _06816_, _06814_);
  and (_06817_, _06809_, _03071_);
  and (_06819_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or (_07286_, _06819_, _06817_);
  and (_06820_, _06809_, _03074_);
  and (_06822_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or (_07289_, _06822_, _06820_);
  and (_06823_, _06809_, _03077_);
  and (_06825_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  or (_07293_, _06825_, _06823_);
  and (_06826_, _06809_, _03080_);
  and (_06828_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or (_07296_, _06828_, _06826_);
  and (_06829_, _06809_, _03083_);
  and (_06831_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  or (_07299_, _06831_, _06829_);
  and (_06833_, _06809_, _03087_);
  and (_06834_, _06811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or (_07301_, _06834_, _06833_);
  and (_06835_, _06702_, _03159_);
  and (_06837_, _06835_, _03060_);
  not (_06838_, _06835_);
  and (_06839_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_07305_, _06839_, _06837_);
  and (_06841_, _06835_, _03067_);
  and (_06842_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_07308_, _06842_, _06841_);
  and (_06844_, _06835_, _03071_);
  and (_06845_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_07311_, _06845_, _06844_);
  and (_06847_, _06835_, _03074_);
  and (_06848_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_07314_, _06848_, _06847_);
  and (_06850_, _06835_, _03077_);
  and (_06851_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_07317_, _06851_, _06850_);
  and (_06853_, _06835_, _03080_);
  and (_06854_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_07321_, _06854_, _06853_);
  and (_06856_, _06835_, _03083_);
  and (_06858_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_07324_, _06858_, _06856_);
  and (_06859_, _06835_, _03087_);
  and (_06860_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_07326_, _06860_, _06859_);
  and (_06862_, _06702_, _03179_);
  and (_06863_, _06862_, _03060_);
  not (_06865_, _06862_);
  and (_06866_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_07330_, _06866_, _06863_);
  and (_06868_, _06862_, _03067_);
  and (_06869_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_07333_, _06869_, _06868_);
  and (_06871_, _06862_, _03071_);
  and (_06872_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_07336_, _06872_, _06871_);
  and (_06874_, _06862_, _03074_);
  and (_06875_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_07339_, _06875_, _06874_);
  and (_06877_, _06862_, _03077_);
  and (_06878_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_07342_, _06878_, _06877_);
  and (_06880_, _06862_, _03080_);
  and (_06881_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_07345_, _06881_, _06880_);
  and (_06883_, _06862_, _03083_);
  and (_06884_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_07348_, _06884_, _06883_);
  and (_06886_, _06862_, _03087_);
  and (_06887_, _06865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_07351_, _06887_, _06886_);
  and (_06889_, _06702_, _03198_);
  and (_06890_, _06889_, _03060_);
  not (_06891_, _06889_);
  and (_06893_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or (_07354_, _06893_, _06890_);
  and (_06894_, _06889_, _03067_);
  and (_06896_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or (_07357_, _06896_, _06894_);
  and (_06897_, _06889_, _03071_);
  and (_06899_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or (_07360_, _06899_, _06897_);
  and (_06900_, _06889_, _03074_);
  and (_06902_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  or (_07363_, _06902_, _06900_);
  and (_06903_, _06889_, _03077_);
  and (_06905_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  or (_07366_, _06905_, _06903_);
  and (_06907_, _06889_, _03080_);
  and (_06908_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  or (_07369_, _06908_, _06907_);
  and (_06909_, _06889_, _03083_);
  and (_06911_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or (_07373_, _06911_, _06909_);
  and (_06912_, _06889_, _03087_);
  and (_06914_, _06891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or (_07375_, _06914_, _06912_);
  and (_06915_, _06702_, _03218_);
  and (_06917_, _06915_, _03060_);
  not (_06918_, _06915_);
  and (_06919_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_07379_, _06919_, _06917_);
  and (_06921_, _06915_, _03067_);
  and (_06922_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_07382_, _06922_, _06921_);
  and (_06924_, _06915_, _03071_);
  and (_06925_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_07385_, _06925_, _06924_);
  and (_06927_, _06915_, _03074_);
  and (_06928_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_07388_, _06928_, _06927_);
  and (_06930_, _06915_, _03077_);
  and (_06932_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_07391_, _06932_, _06930_);
  and (_06933_, _06915_, _03080_);
  and (_06934_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_07394_, _06934_, _06933_);
  and (_06936_, _06915_, _03083_);
  and (_06937_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_07397_, _06937_, _06936_);
  and (_06939_, _06915_, _03087_);
  and (_06940_, _06918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_07400_, _06940_, _06939_);
  and (_06942_, _06702_, _03237_);
  and (_06943_, _06942_, _03060_);
  not (_06945_, _06942_);
  and (_06946_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  or (_07404_, _06946_, _06943_);
  and (_06948_, _06942_, _03067_);
  and (_06949_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  or (_07407_, _06949_, _06948_);
  and (_06951_, _06942_, _03071_);
  and (_06952_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  or (_07410_, _06952_, _06951_);
  and (_06954_, _06942_, _03074_);
  and (_06955_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  or (_07413_, _06955_, _06954_);
  and (_06957_, _06942_, _03077_);
  and (_06958_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or (_07416_, _06958_, _06957_);
  and (_06960_, _06942_, _03080_);
  and (_06961_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  or (_07419_, _06961_, _06960_);
  and (_06963_, _06942_, _03083_);
  and (_06964_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  or (_07422_, _06964_, _06963_);
  and (_06966_, _06942_, _03087_);
  and (_06967_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or (_07424_, _06967_, _06966_);
  and (_06969_, _06702_, _03256_);
  and (_06970_, _06969_, _03060_);
  not (_06971_, _06969_);
  and (_06973_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or (_07428_, _06973_, _06970_);
  and (_06974_, _06969_, _03067_);
  and (_06976_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or (_07431_, _06976_, _06974_);
  and (_06977_, _06969_, _03071_);
  and (_06979_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or (_07434_, _06979_, _06977_);
  and (_06981_, _06969_, _03074_);
  and (_06982_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or (_07437_, _06982_, _06981_);
  and (_06983_, _06969_, _03077_);
  and (_06985_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  or (_07440_, _06985_, _06983_);
  and (_06986_, _06969_, _03080_);
  and (_06988_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or (_07443_, _06988_, _06986_);
  and (_06989_, _06969_, _03083_);
  and (_06991_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or (_07446_, _06991_, _06989_);
  and (_06992_, _06969_, _03087_);
  and (_06994_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  or (_07449_, _06994_, _06992_);
  and (_06995_, _06702_, _03275_);
  and (_06997_, _06995_, _03060_);
  not (_06998_, _06995_);
  and (_06999_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_07453_, _06999_, _06997_);
  and (_07001_, _06995_, _03067_);
  and (_07002_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_07456_, _07002_, _07001_);
  and (_07004_, _06995_, _03071_);
  and (_07006_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_07459_, _07006_, _07004_);
  and (_07007_, _06995_, _03074_);
  and (_07008_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_07462_, _07008_, _07007_);
  and (_07010_, _06995_, _03077_);
  and (_07011_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_07465_, _07011_, _07010_);
  and (_07013_, _06995_, _03080_);
  and (_07014_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_07468_, _07014_, _07013_);
  and (_07016_, _06995_, _03083_);
  and (_07017_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_07471_, _07017_, _07016_);
  and (_07019_, _06995_, _03087_);
  and (_07020_, _06998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_07473_, _07020_, _07019_);
  and (_07022_, _06702_, _03295_);
  and (_07023_, _07022_, _03060_);
  not (_07025_, _07022_);
  and (_07026_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_07477_, _07026_, _07023_);
  and (_07028_, _07022_, _03067_);
  and (_07029_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_07481_, _07029_, _07028_);
  and (_07031_, _07022_, _03071_);
  and (_07032_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_07484_, _07032_, _07031_);
  and (_07034_, _07022_, _03074_);
  and (_07035_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_07487_, _07035_, _07034_);
  and (_07037_, _07022_, _03077_);
  and (_07038_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_07490_, _07038_, _07037_);
  and (_07040_, _07022_, _03080_);
  and (_07041_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_07493_, _07041_, _07040_);
  and (_07043_, _07022_, _03083_);
  and (_07044_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_07496_, _07044_, _07043_);
  and (_07046_, _07022_, _03087_);
  and (_07047_, _07025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_07498_, _07047_, _07046_);
  and (_07049_, _06702_, _03315_);
  and (_07050_, _07049_, _03060_);
  not (_07051_, _07049_);
  and (_07053_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or (_07502_, _07053_, _07050_);
  and (_07055_, _07049_, _03067_);
  and (_07056_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  or (_07505_, _07056_, _07055_);
  and (_07057_, _07049_, _03071_);
  and (_07059_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or (_07508_, _07059_, _07057_);
  and (_07060_, _07049_, _03074_);
  and (_07062_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or (_07511_, _07062_, _07060_);
  and (_07063_, _07049_, _03077_);
  and (_07065_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or (_07514_, _07065_, _07063_);
  and (_07066_, _07049_, _03080_);
  and (_07068_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  or (_07517_, _07068_, _07066_);
  and (_07069_, _07049_, _03083_);
  and (_07071_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  or (_07520_, _07071_, _07069_);
  and (_07072_, _07049_, _03087_);
  and (_07074_, _07051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  or (_07523_, _07074_, _07072_);
  and (_07075_, _06702_, _03334_);
  and (_07077_, _07075_, _03060_);
  not (_07078_, _07075_);
  and (_07080_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  or (_07526_, _07080_, _07077_);
  and (_07081_, _07075_, _03067_);
  and (_07082_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or (_07529_, _07082_, _07081_);
  and (_07084_, _07075_, _03071_);
  and (_07085_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  or (_07533_, _07085_, _07084_);
  and (_07087_, _07075_, _03074_);
  and (_07088_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  or (_07536_, _07088_, _07087_);
  and (_07090_, _07075_, _03077_);
  and (_07091_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  or (_07539_, _07091_, _07090_);
  and (_07093_, _07075_, _03080_);
  and (_07094_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or (_07542_, _07094_, _07093_);
  and (_07096_, _07075_, _03083_);
  and (_07097_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or (_07545_, _07097_, _07096_);
  and (_07099_, _07075_, _03087_);
  and (_07100_, _07078_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or (_07547_, _07100_, _07099_);
  and (_07102_, _06702_, _03353_);
  and (_07104_, _07102_, _03060_);
  not (_07105_, _07102_);
  and (_07106_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_07551_, _07106_, _07104_);
  and (_07108_, _07102_, _03067_);
  and (_07109_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_07554_, _07109_, _07108_);
  and (_07111_, _07102_, _03071_);
  and (_07112_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_07557_, _07112_, _07111_);
  and (_07114_, _07102_, _03074_);
  and (_07115_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_07561_, _07115_, _07114_);
  and (_07117_, _07102_, _03077_);
  and (_07118_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_07564_, _07118_, _07117_);
  and (_07120_, _07102_, _03080_);
  and (_07121_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_07567_, _07121_, _07120_);
  and (_07123_, _07102_, _03083_);
  and (_07124_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_07570_, _07124_, _07123_);
  and (_07126_, _07102_, _03087_);
  and (_07127_, _07105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_07572_, _07127_, _07126_);
  and (_07129_, _03699_, _26459_);
  and (_07130_, _07129_, _02963_);
  and (_07131_, _07130_, _03060_);
  not (_07133_, _07130_);
  and (_07134_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_07577_, _07134_, _07131_);
  and (_07136_, _07130_, _03067_);
  and (_07137_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_07580_, _07137_, _07136_);
  and (_07139_, _07130_, _03071_);
  and (_07140_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_07583_, _07140_, _07139_);
  and (_07142_, _07130_, _03074_);
  and (_07143_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_07586_, _07143_, _07142_);
  and (_07145_, _07130_, _03077_);
  and (_07146_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_07589_, _07146_, _07145_);
  and (_07148_, _07130_, _03080_);
  and (_07149_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_07592_, _07149_, _07148_);
  and (_07151_, _07130_, _03083_);
  and (_07152_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_07595_, _07152_, _07151_);
  and (_07154_, _07130_, _03087_);
  and (_07155_, _07133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_07598_, _07155_, _07154_);
  and (_07157_, _07129_, _03062_);
  and (_07158_, _07157_, _03060_);
  not (_07159_, _07157_);
  and (_07161_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  or (_07601_, _07161_, _07158_);
  and (_07162_, _07157_, _03067_);
  and (_07164_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  or (_07604_, _07164_, _07162_);
  and (_07165_, _07157_, _03071_);
  and (_07167_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  or (_07607_, _07167_, _07165_);
  and (_07168_, _07157_, _03074_);
  and (_07170_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  or (_07610_, _07170_, _07168_);
  and (_07171_, _07157_, _03077_);
  and (_07173_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  or (_07614_, _07173_, _07171_);
  and (_07174_, _07157_, _03080_);
  and (_07176_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  or (_07617_, _07176_, _07174_);
  and (_07178_, _07157_, _03083_);
  and (_07179_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  or (_07620_, _07179_, _07178_);
  and (_07180_, _07157_, _03087_);
  and (_07181_, _07159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  or (_07622_, _07181_, _07180_);
  and (_07183_, _07129_, _03091_);
  and (_07184_, _07183_, _03060_);
  not (_07186_, _07183_);
  and (_07187_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  or (_07626_, _07187_, _07184_);
  and (_07189_, _07183_, _03067_);
  and (_07190_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  or (_07629_, _07190_, _07189_);
  and (_07192_, _07183_, _03071_);
  and (_07193_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  or (_07632_, _07193_, _07192_);
  and (_07195_, _07183_, _03074_);
  and (_07196_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  or (_07635_, _07196_, _07195_);
  and (_07198_, _07183_, _03077_);
  and (_07199_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  or (_07638_, _07199_, _07198_);
  and (_07201_, _07183_, _03080_);
  and (_07202_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  or (_07642_, _07202_, _07201_);
  and (_07204_, _07183_, _03083_);
  and (_07205_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  or (_07645_, _07205_, _07204_);
  and (_07207_, _07183_, _03087_);
  and (_07208_, _07186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  or (_07647_, _07208_, _07207_);
  and (_07210_, _07129_, _03113_);
  and (_07211_, _07210_, _03060_);
  not (_07212_, _07210_);
  and (_07214_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_07651_, _07214_, _07211_);
  and (_07215_, _07210_, _03067_);
  and (_07217_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_07654_, _07217_, _07215_);
  and (_07218_, _07210_, _03071_);
  and (_07220_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_07657_, _07220_, _07218_);
  and (_07221_, _07210_, _03074_);
  and (_07223_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_07660_, _07223_, _07221_);
  and (_07224_, _07210_, _03077_);
  and (_07226_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_07663_, _07226_, _07224_);
  and (_07228_, _07210_, _03080_);
  and (_07229_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_07666_, _07229_, _07228_);
  and (_07230_, _07210_, _03083_);
  and (_07232_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_07669_, _07232_, _07230_);
  and (_07233_, _07210_, _03087_);
  and (_07235_, _07212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_07672_, _07235_, _07233_);
  and (_07236_, _07129_, _03136_);
  and (_07238_, _07236_, _03060_);
  not (_07239_, _07236_);
  and (_07240_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_07675_, _07240_, _07238_);
  and (_07242_, _07236_, _03067_);
  and (_07243_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_07678_, _07243_, _07242_);
  and (_07245_, _07236_, _03071_);
  and (_07246_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_07681_, _07246_, _07245_);
  and (_07248_, _07236_, _03074_);
  and (_07249_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_07684_, _07249_, _07248_);
  and (_07251_, _07236_, _03077_);
  and (_07253_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_07687_, _07253_, _07251_);
  and (_07254_, _07236_, _03080_);
  and (_07255_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_07690_, _07255_, _07254_);
  and (_07257_, _07236_, _03083_);
  and (_07258_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_07694_, _07258_, _07257_);
  and (_07260_, _07236_, _03087_);
  and (_07261_, _07239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_07696_, _07261_, _07260_);
  and (_07263_, _07129_, _03159_);
  and (_07264_, _07263_, _03060_);
  not (_07266_, _07263_);
  and (_07267_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  or (_07700_, _07267_, _07264_);
  and (_07269_, _07263_, _03067_);
  and (_07270_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  or (_07703_, _07270_, _07269_);
  and (_07272_, _07263_, _03071_);
  and (_07273_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  or (_07706_, _07273_, _07272_);
  and (_07275_, _07263_, _03074_);
  and (_07276_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  or (_07709_, _07276_, _07275_);
  and (_07278_, _07263_, _03077_);
  and (_07279_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  or (_07712_, _07279_, _07278_);
  and (_07281_, _07263_, _03080_);
  and (_07282_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  or (_07715_, _07282_, _07281_);
  and (_07284_, _07263_, _03083_);
  and (_07285_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  or (_07718_, _07285_, _07284_);
  and (_07287_, _07263_, _03087_);
  and (_07288_, _07266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  or (_07721_, _07288_, _07287_);
  and (_07290_, _07129_, _03179_);
  and (_07291_, _07290_, _03060_);
  not (_07292_, _07290_);
  and (_07294_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  or (_07725_, _07294_, _07291_);
  and (_07295_, _07290_, _03067_);
  and (_07297_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  or (_07728_, _07297_, _07295_);
  and (_07298_, _07290_, _03071_);
  and (_07300_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  or (_07731_, _07300_, _07298_);
  and (_07302_, _07290_, _03074_);
  and (_07303_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  or (_07734_, _07303_, _07302_);
  and (_07304_, _07290_, _03077_);
  and (_07306_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  or (_07737_, _07306_, _07304_);
  and (_07307_, _07290_, _03080_);
  and (_07309_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  or (_07740_, _07309_, _07307_);
  and (_07310_, _07290_, _03083_);
  and (_07312_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  or (_07743_, _07312_, _07310_);
  and (_07313_, _07290_, _03087_);
  and (_07315_, _07292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  or (_07745_, _07315_, _07313_);
  and (_07316_, _07129_, _03198_);
  and (_07318_, _07316_, _03060_);
  not (_07319_, _07316_);
  and (_07320_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_07749_, _07320_, _07318_);
  and (_07322_, _07316_, _03067_);
  and (_07323_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_07752_, _07323_, _07322_);
  and (_07325_, _07316_, _03071_);
  and (_07327_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_07755_, _07327_, _07325_);
  and (_07328_, _07316_, _03074_);
  and (_07329_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_07758_, _07329_, _07328_);
  and (_07331_, _07316_, _03077_);
  and (_07332_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_07761_, _07332_, _07331_);
  and (_07334_, _07316_, _03080_);
  and (_07335_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_07764_, _07335_, _07334_);
  and (_07337_, _07316_, _03083_);
  and (_07338_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_07767_, _07338_, _07337_);
  and (_07340_, _07316_, _03087_);
  and (_07341_, _07319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_07770_, _07341_, _07340_);
  and (_07343_, _07129_, _03218_);
  and (_07344_, _07343_, _03060_);
  not (_07346_, _07343_);
  and (_07347_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  or (_07774_, _07347_, _07344_);
  and (_07349_, _07343_, _03067_);
  and (_07350_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  or (_07777_, _07350_, _07349_);
  and (_07352_, _07343_, _03071_);
  and (_07353_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  or (_07780_, _07353_, _07352_);
  and (_07355_, _07343_, _03074_);
  and (_07356_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  or (_07783_, _07356_, _07355_);
  and (_07358_, _07343_, _03077_);
  and (_07359_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  or (_07786_, _07359_, _07358_);
  and (_07361_, _07343_, _03080_);
  and (_07362_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  or (_07789_, _07362_, _07361_);
  and (_07364_, _07343_, _03083_);
  and (_07365_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  or (_07792_, _07365_, _07364_);
  and (_07367_, _07343_, _03087_);
  and (_07368_, _07346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  or (_07794_, _07368_, _07367_);
  and (_07370_, _07129_, _03237_);
  and (_07371_, _07370_, _03060_);
  not (_07372_, _07370_);
  and (_07374_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_07798_, _07374_, _07371_);
  and (_07376_, _07370_, _03067_);
  and (_07377_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_07802_, _07377_, _07376_);
  and (_07378_, _07370_, _03071_);
  and (_07380_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_07805_, _07380_, _07378_);
  and (_07381_, _07370_, _03074_);
  and (_07383_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_07808_, _07383_, _07381_);
  and (_07384_, _07370_, _03077_);
  and (_07386_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_07811_, _07386_, _07384_);
  and (_07387_, _07370_, _03080_);
  and (_07389_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_07814_, _07389_, _07387_);
  and (_07390_, _07370_, _03083_);
  and (_07392_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_07817_, _07392_, _07390_);
  and (_07393_, _07370_, _03087_);
  and (_07395_, _07372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_07819_, _07395_, _07393_);
  and (_07396_, _07129_, _03256_);
  and (_07398_, _07396_, _03060_);
  not (_07399_, _07396_);
  and (_07401_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_07823_, _07401_, _07398_);
  and (_07402_, _07396_, _03067_);
  and (_07403_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_07826_, _07403_, _07402_);
  and (_07405_, _07396_, _03071_);
  and (_07406_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_07829_, _07406_, _07405_);
  and (_07408_, _07396_, _03074_);
  and (_07409_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_07832_, _07409_, _07408_);
  and (_07411_, _07396_, _03077_);
  and (_07412_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_07835_, _07412_, _07411_);
  and (_07414_, _07396_, _03080_);
  and (_07415_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_07838_, _07415_, _07414_);
  and (_07417_, _07396_, _03083_);
  and (_07418_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_07841_, _07418_, _07417_);
  and (_07420_, _07396_, _03087_);
  and (_07421_, _07399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_07844_, _07421_, _07420_);
  and (_07423_, _07129_, _03275_);
  and (_07425_, _07423_, _03060_);
  not (_07426_, _07423_);
  and (_07427_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  or (_07847_, _07427_, _07425_);
  and (_07429_, _07423_, _03067_);
  and (_07430_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  or (_07850_, _07430_, _07429_);
  and (_07432_, _07423_, _03071_);
  and (_07433_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  or (_07854_, _07433_, _07432_);
  and (_07435_, _07423_, _03074_);
  and (_07436_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  or (_07857_, _07436_, _07435_);
  and (_07438_, _07423_, _03077_);
  and (_07439_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  or (_07860_, _07439_, _07438_);
  and (_07441_, _07423_, _03080_);
  and (_07442_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  or (_07863_, _07442_, _07441_);
  and (_07444_, _07423_, _03083_);
  and (_07445_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  or (_07866_, _07445_, _07444_);
  and (_07447_, _07423_, _03087_);
  and (_07448_, _07426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  or (_07868_, _07448_, _07447_);
  and (_07450_, _07129_, _03295_);
  and (_07451_, _07450_, _03060_);
  not (_07452_, _07450_);
  and (_07454_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  or (_07872_, _07454_, _07451_);
  and (_07455_, _07450_, _03067_);
  and (_07457_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  or (_07875_, _07457_, _07455_);
  and (_07458_, _07450_, _03071_);
  and (_07460_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  or (_07878_, _07460_, _07458_);
  and (_07461_, _07450_, _03074_);
  and (_07463_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  or (_07882_, _07463_, _07461_);
  and (_07464_, _07450_, _03077_);
  and (_07466_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  or (_07885_, _07466_, _07464_);
  and (_07467_, _07450_, _03080_);
  and (_07469_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  or (_07888_, _07469_, _07467_);
  and (_07470_, _07450_, _03083_);
  and (_07472_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  or (_07891_, _07472_, _07470_);
  and (_07474_, _07450_, _03087_);
  and (_07475_, _07452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  or (_07893_, _07475_, _07474_);
  and (_07476_, _07129_, _03315_);
  and (_07478_, _07476_, _03060_);
  not (_07479_, _07476_);
  and (_07480_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_07897_, _07480_, _07478_);
  and (_07482_, _07476_, _03067_);
  and (_07483_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_07900_, _07483_, _07482_);
  and (_07485_, _07476_, _03071_);
  and (_07486_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_07903_, _07486_, _07485_);
  and (_07488_, _07476_, _03074_);
  and (_07489_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_07906_, _07489_, _07488_);
  and (_07491_, _07476_, _03077_);
  and (_07492_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_07909_, _07492_, _07491_);
  and (_07494_, _07476_, _03080_);
  and (_07495_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_07912_, _07495_, _07494_);
  and (_07497_, _07476_, _03083_);
  and (_07499_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_07915_, _07499_, _07497_);
  and (_07500_, _07476_, _03087_);
  and (_07501_, _07479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_07918_, _07501_, _07500_);
  and (_07503_, _07129_, _03334_);
  and (_07504_, _07503_, _03060_);
  not (_07506_, _07503_);
  and (_07507_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_07921_, _07507_, _07504_);
  and (_07509_, _07503_, _03067_);
  and (_07510_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_07924_, _07510_, _07509_);
  and (_07512_, _07503_, _03071_);
  and (_07513_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_07927_, _07513_, _07512_);
  and (_07515_, _07503_, _03074_);
  and (_07516_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_07930_, _07516_, _07515_);
  and (_07518_, _07503_, _03077_);
  and (_07519_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_07934_, _07519_, _07518_);
  and (_07521_, _07503_, _03080_);
  and (_07522_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_07937_, _07522_, _07521_);
  and (_07524_, _07503_, _03083_);
  and (_07525_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_07940_, _07525_, _07524_);
  and (_07527_, _07503_, _03087_);
  and (_07528_, _07506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_07942_, _07528_, _07527_);
  and (_07530_, _07129_, _03353_);
  and (_07531_, _07530_, _03060_);
  not (_07532_, _07530_);
  and (_07534_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  or (_07946_, _07534_, _07531_);
  and (_07535_, _07530_, _03067_);
  and (_07537_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  or (_07949_, _07537_, _07535_);
  and (_07538_, _07530_, _03071_);
  and (_07540_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  or (_07952_, _07540_, _07538_);
  and (_07541_, _07530_, _03074_);
  and (_07543_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  or (_07955_, _07543_, _07541_);
  and (_07544_, _07530_, _03077_);
  and (_07546_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  or (_07958_, _07546_, _07544_);
  and (_07548_, _07530_, _03080_);
  and (_07549_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  or (_07962_, _07549_, _07548_);
  and (_07550_, _07530_, _03083_);
  and (_07552_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  or (_07965_, _07552_, _07550_);
  and (_07553_, _07530_, _03087_);
  and (_07555_, _07532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  or (_07967_, _07555_, _07553_);
  and (_07556_, _04125_, _26459_);
  and (_07558_, _07556_, _02963_);
  and (_07559_, _07558_, _03060_);
  not (_07560_, _07558_);
  and (_07562_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or (_07971_, _07562_, _07559_);
  and (_07563_, _07558_, _03067_);
  and (_07565_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or (_07974_, _07565_, _07563_);
  and (_07566_, _07558_, _03071_);
  and (_07568_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or (_07977_, _07568_, _07566_);
  and (_07569_, _07558_, _03074_);
  and (_07571_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or (_07980_, _07571_, _07569_);
  and (_07573_, _07558_, _03077_);
  and (_07574_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or (_07983_, _07574_, _07573_);
  and (_07575_, _07558_, _03080_);
  and (_07576_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or (_07987_, _07576_, _07575_);
  and (_07578_, _07558_, _03083_);
  and (_07579_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or (_07991_, _07579_, _07578_);
  and (_07581_, _07558_, _03087_);
  and (_07582_, _07560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or (_07993_, _07582_, _07581_);
  and (_07584_, _07556_, _03062_);
  and (_07585_, _07584_, _03060_);
  not (_07587_, _07584_);
  and (_07588_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_07997_, _07588_, _07585_);
  and (_07590_, _07584_, _03067_);
  and (_07591_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_08000_, _07591_, _07590_);
  and (_07593_, _07584_, _03071_);
  and (_07594_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_08003_, _07594_, _07593_);
  and (_07596_, _07584_, _03074_);
  and (_07597_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_08006_, _07597_, _07596_);
  and (_07599_, _07584_, _03077_);
  and (_07600_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_08009_, _07600_, _07599_);
  and (_07602_, _07584_, _03080_);
  and (_07603_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_08012_, _07603_, _07602_);
  and (_07605_, _07584_, _03083_);
  and (_07606_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_08015_, _07606_, _07605_);
  and (_07608_, _07584_, _03087_);
  and (_07609_, _07587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_08018_, _07609_, _07608_);
  and (_07611_, _07556_, _03091_);
  and (_07612_, _07611_, _03060_);
  not (_07613_, _07611_);
  and (_07615_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_08021_, _07615_, _07612_);
  and (_07616_, _07611_, _03067_);
  and (_07618_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_08024_, _07618_, _07616_);
  and (_07619_, _07611_, _03071_);
  and (_07621_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_08027_, _07621_, _07619_);
  and (_07623_, _07611_, _03074_);
  and (_07624_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_08030_, _07624_, _07623_);
  and (_07625_, _07611_, _03077_);
  and (_07627_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_08033_, _07627_, _07625_);
  and (_07628_, _07611_, _03080_);
  and (_07630_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_08036_, _07630_, _07628_);
  and (_07631_, _07611_, _03083_);
  and (_07633_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_08039_, _07633_, _07631_);
  and (_07634_, _07611_, _03087_);
  and (_07636_, _07613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_08042_, _07636_, _07634_);
  and (_07637_, _07556_, _03113_);
  and (_07639_, _07637_, _03060_);
  not (_07640_, _07637_);
  and (_07641_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or (_08046_, _07641_, _07639_);
  and (_07643_, _07637_, _03067_);
  and (_07644_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or (_08049_, _07644_, _07643_);
  and (_07646_, _07637_, _03071_);
  and (_07648_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or (_08052_, _07648_, _07646_);
  and (_07649_, _07637_, _03074_);
  and (_07650_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or (_08055_, _07650_, _07649_);
  and (_07652_, _07637_, _03077_);
  and (_07653_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or (_08058_, _07653_, _07652_);
  and (_07655_, _07637_, _03080_);
  and (_07656_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or (_08061_, _07656_, _07655_);
  and (_07658_, _07637_, _03083_);
  and (_07659_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or (_08064_, _07659_, _07658_);
  and (_07661_, _07637_, _03087_);
  and (_07662_, _07640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or (_08066_, _07662_, _07661_);
  and (_07664_, _07556_, _03136_);
  and (_07665_, _07664_, _03060_);
  not (_07667_, _07664_);
  and (_07668_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or (_08071_, _07668_, _07665_);
  and (_07670_, _07664_, _03067_);
  and (_07671_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or (_08074_, _07671_, _07670_);
  and (_07673_, _07664_, _03071_);
  and (_07674_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or (_08077_, _07674_, _07673_);
  and (_07676_, _07664_, _03074_);
  and (_07677_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or (_08080_, _07677_, _07676_);
  and (_07679_, _07664_, _03077_);
  and (_07680_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or (_08083_, _07680_, _07679_);
  and (_07682_, _07664_, _03080_);
  and (_07683_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or (_08086_, _07683_, _07682_);
  and (_07685_, _07664_, _03083_);
  and (_07686_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or (_08089_, _07686_, _07685_);
  and (_07688_, _07664_, _03087_);
  and (_07689_, _07667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or (_08091_, _07689_, _07688_);
  and (_07691_, _07556_, _03159_);
  and (_07692_, _07691_, _03060_);
  not (_07693_, _07691_);
  and (_07695_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_08095_, _07695_, _07692_);
  and (_07697_, _07691_, _03067_);
  and (_07698_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_08098_, _07698_, _07697_);
  and (_07699_, _07691_, _03071_);
  and (_07701_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_08101_, _07701_, _07699_);
  and (_07702_, _07691_, _03074_);
  and (_07704_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_08104_, _07704_, _07702_);
  and (_07705_, _07691_, _03077_);
  and (_07707_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_08107_, _07707_, _07705_);
  and (_07708_, _07691_, _03080_);
  and (_07710_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_08110_, _07710_, _07708_);
  and (_07711_, _07691_, _03083_);
  and (_07713_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_08113_, _07713_, _07711_);
  and (_07714_, _07691_, _03087_);
  and (_07716_, _07693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_08116_, _07716_, _07714_);
  and (_07717_, _07556_, _03179_);
  and (_07719_, _07717_, _03060_);
  not (_07720_, _07717_);
  and (_07722_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_08119_, _07722_, _07719_);
  and (_07723_, _07717_, _03067_);
  and (_07724_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_08123_, _07724_, _07723_);
  and (_07726_, _07717_, _03071_);
  and (_07727_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_08126_, _07727_, _07726_);
  and (_07729_, _07717_, _03074_);
  and (_07730_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_08129_, _07730_, _07729_);
  and (_07732_, _07717_, _03077_);
  and (_07733_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_08132_, _07733_, _07732_);
  and (_07735_, _07717_, _03080_);
  and (_07736_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_08135_, _07736_, _07735_);
  and (_07738_, _07717_, _03083_);
  and (_07739_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_08138_, _07739_, _07738_);
  and (_07741_, _07717_, _03087_);
  and (_07742_, _07720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_08140_, _07742_, _07741_);
  and (_07744_, _07556_, _03198_);
  and (_07746_, _07744_, _03060_);
  not (_07747_, _07744_);
  and (_07748_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or (_08144_, _07748_, _07746_);
  and (_07750_, _07744_, _03067_);
  and (_07751_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or (_08147_, _07751_, _07750_);
  and (_07753_, _07744_, _03071_);
  and (_07754_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or (_08151_, _07754_, _07753_);
  and (_07756_, _07744_, _03074_);
  and (_07757_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or (_08154_, _07757_, _07756_);
  and (_07759_, _07744_, _03077_);
  and (_07760_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or (_08157_, _07760_, _07759_);
  and (_07762_, _07744_, _03080_);
  and (_07763_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or (_08160_, _07763_, _07762_);
  and (_07765_, _07744_, _03083_);
  and (_07766_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or (_08163_, _07766_, _07765_);
  and (_07768_, _07744_, _03087_);
  and (_07769_, _07747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or (_08165_, _07769_, _07768_);
  and (_07771_, _07556_, _03218_);
  and (_07772_, _07771_, _03060_);
  not (_07773_, _07771_);
  and (_07775_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_08169_, _07775_, _07772_);
  and (_07776_, _07771_, _03067_);
  and (_07778_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_08172_, _07778_, _07776_);
  and (_07779_, _07771_, _03071_);
  and (_07781_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_08175_, _07781_, _07779_);
  and (_07782_, _07771_, _03074_);
  and (_07784_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_08178_, _07784_, _07782_);
  and (_07785_, _07771_, _03077_);
  and (_07787_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_08181_, _07787_, _07785_);
  and (_07788_, _07771_, _03080_);
  and (_07790_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_08184_, _07790_, _07788_);
  and (_07791_, _07771_, _03083_);
  and (_07793_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_08187_, _07793_, _07791_);
  and (_07795_, _07771_, _03087_);
  and (_07796_, _07773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_08190_, _07796_, _07795_);
  and (_07797_, _07556_, _03237_);
  and (_07799_, _07797_, _03060_);
  not (_07800_, _07797_);
  and (_07801_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or (_08193_, _07801_, _07799_);
  and (_07803_, _07797_, _03067_);
  and (_07804_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or (_08196_, _07804_, _07803_);
  and (_07806_, _07797_, _03071_);
  and (_07807_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or (_08199_, _07807_, _07806_);
  and (_07809_, _07797_, _03074_);
  and (_07810_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or (_08203_, _07810_, _07809_);
  and (_07812_, _07797_, _03077_);
  and (_07813_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or (_08206_, _07813_, _07812_);
  and (_07815_, _07797_, _03080_);
  and (_07816_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or (_08209_, _07816_, _07815_);
  and (_07818_, _07797_, _03083_);
  and (_07820_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or (_08212_, _07820_, _07818_);
  and (_07821_, _07797_, _03087_);
  and (_07822_, _07800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or (_08214_, _07822_, _07821_);
  and (_07824_, _07556_, _03256_);
  and (_07825_, _07824_, _03060_);
  not (_07827_, _07824_);
  and (_07828_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or (_08218_, _07828_, _07825_);
  and (_07830_, _07824_, _03067_);
  and (_07831_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or (_08221_, _07831_, _07830_);
  and (_07833_, _07824_, _03071_);
  and (_07834_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or (_08224_, _07834_, _07833_);
  and (_07836_, _07824_, _03074_);
  and (_07837_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or (_08227_, _07837_, _07836_);
  and (_07839_, _07824_, _03077_);
  and (_07840_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or (_08231_, _07840_, _07839_);
  and (_07842_, _07824_, _03080_);
  and (_07843_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or (_08234_, _07843_, _07842_);
  and (_07845_, _07824_, _03083_);
  and (_07846_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or (_08237_, _07846_, _07845_);
  and (_07848_, _07824_, _03087_);
  and (_07849_, _07827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or (_08239_, _07849_, _07848_);
  and (_07851_, _07556_, _03275_);
  and (_07852_, _07851_, _03060_);
  not (_07853_, _07851_);
  and (_07855_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_08243_, _07855_, _07852_);
  and (_07856_, _07851_, _03067_);
  and (_07858_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_08246_, _07858_, _07856_);
  and (_07859_, _07851_, _03071_);
  and (_07861_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_08249_, _07861_, _07859_);
  and (_07862_, _07851_, _03074_);
  and (_07864_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_08252_, _07864_, _07862_);
  and (_07865_, _07851_, _03077_);
  and (_07867_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_08255_, _07867_, _07865_);
  and (_07869_, _07851_, _03080_);
  and (_07870_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_08258_, _07870_, _07869_);
  and (_07871_, _07851_, _03083_);
  and (_07873_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_08261_, _07873_, _07871_);
  and (_07874_, _07851_, _03087_);
  and (_07876_, _07853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_08264_, _07876_, _07874_);
  and (_07877_, _07556_, _03295_);
  and (_07879_, _07877_, _03060_);
  not (_07880_, _07877_);
  and (_07881_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_08267_, _07881_, _07879_);
  and (_07883_, _07877_, _03067_);
  and (_07884_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_08270_, _07884_, _07883_);
  and (_07886_, _07877_, _03071_);
  and (_07887_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_08273_, _07887_, _07886_);
  and (_07889_, _07877_, _03074_);
  and (_07890_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_08276_, _07890_, _07889_);
  and (_07892_, _07877_, _03077_);
  and (_07894_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_08279_, _07894_, _07892_);
  and (_07895_, _07877_, _03080_);
  and (_07896_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_08283_, _07896_, _07895_);
  and (_07898_, _07877_, _03083_);
  and (_07899_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_08286_, _07899_, _07898_);
  and (_07901_, _07877_, _03087_);
  and (_07902_, _07880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_08288_, _07902_, _07901_);
  and (_07904_, _07556_, _03315_);
  and (_07905_, _07904_, _03060_);
  not (_07907_, _07904_);
  and (_07908_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or (_08292_, _07908_, _07905_);
  and (_07910_, _07904_, _03067_);
  and (_07911_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or (_08295_, _07911_, _07910_);
  and (_07913_, _07904_, _03071_);
  and (_07914_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or (_08298_, _07914_, _07913_);
  and (_07916_, _07904_, _03074_);
  and (_07917_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or (_08301_, _07917_, _07916_);
  and (_07919_, _07904_, _03077_);
  and (_07920_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or (_08304_, _07920_, _07919_);
  and (_07922_, _07904_, _03080_);
  and (_07923_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or (_08307_, _07923_, _07922_);
  and (_07925_, _07904_, _03083_);
  and (_07926_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or (_08311_, _07926_, _07925_);
  and (_07928_, _07904_, _03087_);
  and (_07929_, _07907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or (_08313_, _07929_, _07928_);
  and (_07931_, _07556_, _03334_);
  and (_07932_, _07931_, _03060_);
  not (_07933_, _07931_);
  and (_07935_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or (_08317_, _07935_, _07932_);
  and (_07936_, _07931_, _03067_);
  and (_07938_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or (_08320_, _07938_, _07936_);
  and (_07939_, _07931_, _03071_);
  and (_07941_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or (_08323_, _07941_, _07939_);
  and (_07943_, _07931_, _03074_);
  and (_07944_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or (_08326_, _07944_, _07943_);
  and (_07945_, _07931_, _03077_);
  and (_07947_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or (_08329_, _07947_, _07945_);
  and (_07948_, _07931_, _03080_);
  and (_07950_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or (_08332_, _07950_, _07948_);
  and (_07951_, _07931_, _03083_);
  and (_07953_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or (_08335_, _07953_, _07951_);
  and (_07954_, _07931_, _03087_);
  and (_07956_, _07933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or (_08338_, _07956_, _07954_);
  and (_07957_, _07556_, _03353_);
  and (_07959_, _07957_, _03060_);
  not (_07960_, _07957_);
  and (_07961_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_08341_, _07961_, _07959_);
  and (_07963_, _07957_, _03067_);
  and (_07964_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_08344_, _07964_, _07963_);
  and (_07966_, _07957_, _03071_);
  and (_07968_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_08347_, _07968_, _07966_);
  and (_07969_, _07957_, _03074_);
  and (_07970_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_08350_, _07970_, _07969_);
  and (_07972_, _07957_, _03077_);
  and (_07973_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_08353_, _07973_, _07972_);
  and (_07975_, _07957_, _03080_);
  and (_07976_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_08356_, _07976_, _07975_);
  and (_07978_, _07957_, _03083_);
  and (_07979_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_08359_, _07979_, _07978_);
  and (_07981_, _07957_, _03087_);
  and (_07982_, _07960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_08362_, _07982_, _07981_);
  and (_07984_, _02137_, _26939_);
  and (_07985_, _07984_, _02966_);
  and (_07986_, _07985_, _02963_);
  and (_07988_, _07986_, _03060_);
  not (_07989_, _07986_);
  and (_07990_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_08367_, _07990_, _07988_);
  and (_07992_, _07986_, _03067_);
  and (_07994_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_08370_, _07994_, _07992_);
  and (_07995_, _07986_, _03071_);
  and (_07996_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_08373_, _07996_, _07995_);
  and (_07998_, _07986_, _03074_);
  and (_07999_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_08376_, _07999_, _07998_);
  and (_08001_, _07986_, _03077_);
  and (_08002_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_08379_, _08002_, _08001_);
  and (_08004_, _07986_, _03080_);
  and (_08005_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_08382_, _08005_, _08004_);
  and (_08007_, _07986_, _03083_);
  and (_08008_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_08385_, _08008_, _08007_);
  and (_08010_, _07986_, _03087_);
  and (_08011_, _07989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_08388_, _08011_, _08010_);
  and (_08013_, _07985_, _03062_);
  and (_08014_, _08013_, _03060_);
  not (_08016_, _08013_);
  and (_08017_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or (_08392_, _08017_, _08014_);
  and (_08019_, _08013_, _03067_);
  and (_08020_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or (_08395_, _08020_, _08019_);
  and (_08022_, _08013_, _03071_);
  and (_08023_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or (_08398_, _08023_, _08022_);
  and (_08025_, _08013_, _03074_);
  and (_08026_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or (_08401_, _08026_, _08025_);
  and (_08028_, _08013_, _03077_);
  and (_08029_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or (_08404_, _08029_, _08028_);
  and (_08031_, _08013_, _03080_);
  and (_08032_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_08407_, _08032_, _08031_);
  and (_08034_, _08013_, _03083_);
  and (_08035_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or (_08410_, _08035_, _08034_);
  and (_08037_, _08013_, _03087_);
  and (_08038_, _08016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or (_08412_, _08038_, _08037_);
  and (_08040_, _07985_, _03091_);
  and (_08041_, _08040_, _03060_);
  not (_08043_, _08040_);
  and (_08044_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_08417_, _08044_, _08041_);
  and (_08045_, _08040_, _03067_);
  and (_08047_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or (_08420_, _08047_, _08045_);
  and (_08048_, _08040_, _03071_);
  and (_08050_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or (_08423_, _08050_, _08048_);
  and (_08051_, _08040_, _03074_);
  and (_08053_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or (_08426_, _08053_, _08051_);
  and (_08054_, _08040_, _03077_);
  and (_08056_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or (_08429_, _08056_, _08054_);
  and (_08057_, _08040_, _03080_);
  and (_08059_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_08432_, _08059_, _08057_);
  and (_08060_, _08040_, _03083_);
  and (_08062_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or (_08435_, _08062_, _08060_);
  and (_08063_, _08040_, _03087_);
  and (_08065_, _08043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or (_08437_, _08065_, _08063_);
  and (_08067_, _07985_, _03113_);
  and (_08068_, _08067_, _03060_);
  not (_08069_, _08067_);
  and (_08070_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_08441_, _08070_, _08068_);
  and (_08072_, _08067_, _03067_);
  and (_08073_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_08445_, _08073_, _08072_);
  and (_08075_, _08067_, _03071_);
  and (_08076_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_08448_, _08076_, _08075_);
  and (_08078_, _08067_, _03074_);
  and (_08079_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_08451_, _08079_, _08078_);
  and (_08081_, _08067_, _03077_);
  and (_08082_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_08454_, _08082_, _08081_);
  and (_08084_, _08067_, _03080_);
  and (_08085_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_08457_, _08085_, _08084_);
  and (_08087_, _08067_, _03083_);
  and (_08088_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_08460_, _08088_, _08087_);
  and (_08090_, _08067_, _03087_);
  and (_08092_, _08069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_08462_, _08092_, _08090_);
  and (_08093_, _07985_, _03136_);
  and (_08094_, _08093_, _03060_);
  not (_08096_, _08093_);
  and (_08097_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_08466_, _08097_, _08094_);
  and (_08099_, _08093_, _03067_);
  and (_08100_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_08469_, _08100_, _08099_);
  and (_08102_, _08093_, _03071_);
  and (_08103_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_08472_, _08103_, _08102_);
  and (_08105_, _08093_, _03074_);
  and (_08106_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_08475_, _08106_, _08105_);
  and (_08108_, _08093_, _03077_);
  and (_08109_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_08478_, _08109_, _08108_);
  and (_08111_, _08093_, _03080_);
  and (_08112_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_08481_, _08112_, _08111_);
  and (_08114_, _08093_, _03083_);
  and (_08115_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_08484_, _08115_, _08114_);
  and (_08117_, _08093_, _03087_);
  and (_08118_, _08096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_08487_, _08118_, _08117_);
  and (_08120_, _07985_, _03159_);
  and (_08121_, _08120_, _03060_);
  not (_08122_, _08120_);
  and (_08124_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or (_08490_, _08124_, _08121_);
  and (_08125_, _08120_, _03067_);
  and (_08127_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or (_08493_, _08127_, _08125_);
  and (_08128_, _08120_, _03071_);
  and (_08130_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or (_08497_, _08130_, _08128_);
  and (_08131_, _08120_, _03074_);
  and (_08133_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or (_08500_, _08133_, _08131_);
  and (_08134_, _08120_, _03077_);
  and (_08136_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or (_08503_, _08136_, _08134_);
  and (_08137_, _08120_, _03080_);
  and (_08139_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_08506_, _08139_, _08137_);
  and (_08141_, _08120_, _03083_);
  and (_08142_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or (_08509_, _08142_, _08141_);
  and (_08143_, _08120_, _03087_);
  and (_08145_, _08122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or (_08511_, _08145_, _08143_);
  and (_08146_, _07985_, _03179_);
  and (_08148_, _08146_, _03060_);
  not (_08149_, _08146_);
  and (_08150_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_08515_, _08150_, _08148_);
  and (_08152_, _08146_, _03067_);
  and (_08153_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or (_08518_, _08153_, _08152_);
  and (_08155_, _08146_, _03071_);
  and (_08156_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or (_08521_, _08156_, _08155_);
  and (_08158_, _08146_, _03074_);
  and (_08159_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or (_08525_, _08159_, _08158_);
  and (_08161_, _08146_, _03077_);
  and (_08162_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or (_08528_, _08162_, _08161_);
  and (_08164_, _08146_, _03080_);
  and (_08166_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_08531_, _08166_, _08164_);
  and (_08167_, _08146_, _03083_);
  and (_08168_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or (_08534_, _08168_, _08167_);
  and (_08170_, _08146_, _03087_);
  and (_08171_, _08149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or (_08536_, _08171_, _08170_);
  and (_08173_, _07985_, _03198_);
  and (_08174_, _08173_, _03060_);
  not (_08176_, _08173_);
  and (_08177_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_08540_, _08177_, _08174_);
  and (_08179_, _08173_, _03067_);
  and (_08180_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_08543_, _08180_, _08179_);
  and (_08182_, _08173_, _03071_);
  and (_08183_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_08546_, _08183_, _08182_);
  and (_08185_, _08173_, _03074_);
  and (_08186_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_08549_, _08186_, _08185_);
  and (_08188_, _08173_, _03077_);
  and (_08189_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_08552_, _08189_, _08188_);
  and (_08191_, _08173_, _03080_);
  and (_08192_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_08555_, _08192_, _08191_);
  and (_08194_, _08173_, _03083_);
  and (_08195_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_08558_, _08195_, _08194_);
  and (_08197_, _08173_, _03087_);
  and (_08198_, _08176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_08561_, _08198_, _08197_);
  and (_08200_, _07985_, _03218_);
  and (_08201_, _08200_, _03060_);
  not (_08202_, _08200_);
  and (_08204_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_08564_, _08204_, _08201_);
  and (_08205_, _08200_, _03067_);
  and (_08207_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or (_08567_, _08207_, _08205_);
  and (_08208_, _08200_, _03071_);
  and (_08210_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or (_08570_, _08210_, _08208_);
  and (_08211_, _08200_, _03074_);
  and (_08213_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or (_08573_, _08213_, _08211_);
  and (_08215_, _08200_, _03077_);
  and (_08216_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or (_08577_, _08216_, _08215_);
  and (_08217_, _08200_, _03080_);
  and (_08219_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_08580_, _08219_, _08217_);
  and (_08220_, _08200_, _03083_);
  and (_08222_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or (_08583_, _08222_, _08220_);
  and (_08223_, _08200_, _03087_);
  and (_08225_, _08202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_08585_, _08225_, _08223_);
  and (_08226_, _07985_, _03237_);
  and (_08228_, _08226_, _03060_);
  not (_08229_, _08226_);
  and (_08230_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_08589_, _08230_, _08228_);
  and (_08232_, _08226_, _03067_);
  and (_08233_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_08592_, _08233_, _08232_);
  and (_08235_, _08226_, _03071_);
  and (_08236_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_08595_, _08236_, _08235_);
  and (_08238_, _08226_, _03074_);
  and (_08240_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_08598_, _08240_, _08238_);
  and (_08241_, _08226_, _03077_);
  and (_08242_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_08601_, _08242_, _08241_);
  and (_08244_, _08226_, _03080_);
  and (_08245_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_08605_, _08245_, _08244_);
  and (_08247_, _08226_, _03083_);
  and (_08248_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_08608_, _08248_, _08247_);
  and (_08250_, _08226_, _03087_);
  and (_08251_, _08229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_08610_, _08251_, _08250_);
  and (_08253_, _07985_, _03256_);
  and (_08254_, _08253_, _03060_);
  not (_08256_, _08253_);
  and (_08257_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_08614_, _08257_, _08254_);
  and (_08259_, _08253_, _03067_);
  and (_08260_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_08617_, _08260_, _08259_);
  and (_08262_, _08253_, _03071_);
  and (_08263_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_08620_, _08263_, _08262_);
  and (_08265_, _08253_, _03074_);
  and (_08266_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_08623_, _08266_, _08265_);
  and (_08268_, _08253_, _03077_);
  and (_08269_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_08626_, _08269_, _08268_);
  and (_08271_, _08253_, _03080_);
  and (_08272_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_08629_, _08272_, _08271_);
  and (_08274_, _08253_, _03083_);
  and (_08275_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_08632_, _08275_, _08274_);
  and (_08277_, _08253_, _03087_);
  and (_08278_, _08256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_08635_, _08278_, _08277_);
  and (_08280_, _07985_, _03275_);
  and (_08281_, _08280_, _03060_);
  not (_08282_, _08280_);
  and (_08284_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or (_08638_, _08284_, _08281_);
  and (_08285_, _08280_, _03067_);
  and (_08287_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or (_08641_, _08287_, _08285_);
  and (_08289_, _08280_, _03071_);
  and (_08290_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or (_08644_, _08290_, _08289_);
  and (_08291_, _08280_, _03074_);
  and (_08293_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or (_08647_, _08293_, _08291_);
  and (_08294_, _08280_, _03077_);
  and (_08296_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or (_08650_, _08296_, _08294_);
  and (_08297_, _08280_, _03080_);
  and (_08299_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_08653_, _08299_, _08297_);
  and (_08300_, _08280_, _03083_);
  and (_08302_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or (_08657_, _08302_, _08300_);
  and (_08303_, _08280_, _03087_);
  and (_08305_, _08282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or (_08659_, _08305_, _08303_);
  and (_08306_, _07985_, _03295_);
  and (_08308_, _08306_, _03060_);
  not (_08309_, _08306_);
  and (_08310_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_08663_, _08310_, _08308_);
  and (_08312_, _08306_, _03067_);
  and (_08314_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or (_08666_, _08314_, _08312_);
  and (_08315_, _08306_, _03071_);
  and (_08316_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or (_08669_, _08316_, _08315_);
  and (_08318_, _08306_, _03074_);
  and (_08319_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or (_08672_, _08319_, _08318_);
  and (_08321_, _08306_, _03077_);
  and (_08322_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or (_08675_, _08322_, _08321_);
  and (_08324_, _08306_, _03080_);
  and (_08325_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_08678_, _08325_, _08324_);
  and (_08327_, _08306_, _03083_);
  and (_08328_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or (_08681_, _08328_, _08327_);
  and (_08330_, _08306_, _03087_);
  and (_08331_, _08309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or (_08684_, _08331_, _08330_);
  and (_08333_, _07985_, _03315_);
  and (_08334_, _08333_, _03060_);
  not (_08336_, _08333_);
  and (_08337_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_08688_, _08337_, _08334_);
  and (_08339_, _08333_, _03067_);
  and (_08340_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_08691_, _08340_, _08339_);
  and (_08342_, _08333_, _03071_);
  and (_08343_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_08694_, _08343_, _08342_);
  and (_08345_, _08333_, _03074_);
  and (_08346_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_08697_, _08346_, _08345_);
  and (_08348_, _08333_, _03077_);
  and (_08349_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_08700_, _08349_, _08348_);
  and (_08351_, _08333_, _03080_);
  and (_08352_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_08703_, _08352_, _08351_);
  and (_08354_, _08333_, _03083_);
  and (_08355_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_08706_, _08355_, _08354_);
  and (_08357_, _08333_, _03087_);
  and (_08358_, _08336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_08708_, _08358_, _08357_);
  and (_08360_, _07985_, _03334_);
  and (_08361_, _08360_, _03060_);
  not (_08363_, _08360_);
  and (_08364_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_08712_, _08364_, _08361_);
  and (_08365_, _08360_, _03067_);
  and (_08366_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_08715_, _08366_, _08365_);
  and (_08368_, _08360_, _03071_);
  and (_08369_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_08718_, _08369_, _08368_);
  and (_08371_, _08360_, _03074_);
  and (_08372_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_08721_, _08372_, _08371_);
  and (_08374_, _08360_, _03077_);
  and (_08375_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_08724_, _08375_, _08374_);
  and (_08377_, _08360_, _03080_);
  and (_08378_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_08727_, _08378_, _08377_);
  and (_08380_, _08360_, _03083_);
  and (_08381_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_08730_, _08381_, _08380_);
  and (_08383_, _08360_, _03087_);
  and (_08384_, _08363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_08733_, _08384_, _08383_);
  and (_08386_, _07985_, _03353_);
  and (_08387_, _08386_, _03060_);
  not (_08389_, _08386_);
  and (_08390_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_08737_, _08390_, _08387_);
  and (_08391_, _08386_, _03067_);
  and (_08393_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or (_08740_, _08393_, _08391_);
  and (_08394_, _08386_, _03071_);
  and (_08396_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or (_08743_, _08396_, _08394_);
  and (_08397_, _08386_, _03074_);
  and (_08399_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or (_08746_, _08399_, _08397_);
  and (_08400_, _08386_, _03077_);
  and (_08402_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or (_08749_, _08402_, _08400_);
  and (_08403_, _08386_, _03080_);
  and (_08405_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_08752_, _08405_, _08403_);
  and (_08406_, _08386_, _03083_);
  and (_08408_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or (_08755_, _08408_, _08406_);
  and (_08409_, _08386_, _03087_);
  and (_08411_, _08389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or (_08757_, _08411_, _08409_);
  and (_08413_, _03373_, _26939_);
  and (_08414_, _08413_, _02963_);
  and (_08415_, _08414_, _03060_);
  not (_08416_, _08414_);
  and (_08418_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  or (_08762_, _08418_, _08415_);
  and (_08419_, _08414_, _03067_);
  and (_08421_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  or (_08765_, _08421_, _08419_);
  and (_08422_, _08414_, _03071_);
  and (_08424_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  or (_08768_, _08424_, _08422_);
  and (_08425_, _08414_, _03074_);
  and (_08427_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  or (_08771_, _08427_, _08425_);
  and (_08428_, _08414_, _03077_);
  and (_08430_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  or (_08774_, _08430_, _08428_);
  and (_08431_, _08414_, _03080_);
  and (_08433_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  or (_08777_, _08433_, _08431_);
  and (_08434_, _08414_, _03083_);
  and (_08436_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  or (_08780_, _08436_, _08434_);
  and (_08438_, _08414_, _03087_);
  and (_08439_, _08416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  or (_08783_, _08439_, _08438_);
  and (_08440_, _08413_, _03062_);
  and (_08442_, _08440_, _03060_);
  not (_08443_, _08440_);
  and (_08444_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_08786_, _08444_, _08442_);
  and (_08446_, _08440_, _03067_);
  and (_08447_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_08790_, _08447_, _08446_);
  and (_08449_, _08440_, _03071_);
  and (_08450_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_08793_, _08450_, _08449_);
  and (_08452_, _08440_, _03074_);
  and (_08453_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_08796_, _08453_, _08452_);
  and (_08455_, _08440_, _03077_);
  and (_08456_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_08799_, _08456_, _08455_);
  and (_08458_, _08440_, _03080_);
  and (_08459_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_08802_, _08459_, _08458_);
  and (_08461_, _08440_, _03083_);
  and (_08463_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_08805_, _08463_, _08461_);
  and (_08464_, _08440_, _03087_);
  and (_08465_, _08443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_08807_, _08465_, _08464_);
  and (_08467_, _08413_, _03091_);
  and (_08468_, _08467_, _03060_);
  not (_08470_, _08467_);
  and (_08471_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_08811_, _08471_, _08468_);
  and (_08473_, _08467_, _03067_);
  and (_08474_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_08814_, _08474_, _08473_);
  and (_08476_, _08467_, _03071_);
  and (_08477_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_08818_, _08477_, _08476_);
  and (_08479_, _08467_, _03074_);
  and (_08480_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_08821_, _08480_, _08479_);
  and (_08482_, _08467_, _03077_);
  and (_08483_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_08824_, _08483_, _08482_);
  and (_08485_, _08467_, _03080_);
  and (_08486_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_08827_, _08486_, _08485_);
  and (_08488_, _08467_, _03083_);
  and (_08489_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_08830_, _08489_, _08488_);
  and (_08491_, _08467_, _03087_);
  and (_08492_, _08470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_08832_, _08492_, _08491_);
  and (_08494_, _08413_, _03113_);
  and (_08495_, _08494_, _03060_);
  not (_08496_, _08494_);
  and (_08498_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  or (_08836_, _08498_, _08495_);
  and (_08499_, _08494_, _03067_);
  and (_08501_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  or (_08839_, _08501_, _08499_);
  and (_08502_, _08494_, _03071_);
  and (_08504_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  or (_08843_, _08504_, _08502_);
  and (_08505_, _08494_, _03074_);
  and (_08507_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  or (_08847_, _08507_, _08505_);
  and (_08508_, _08494_, _03077_);
  and (_08510_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  or (_08850_, _08510_, _08508_);
  and (_08512_, _08494_, _03080_);
  and (_08513_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  or (_08854_, _08513_, _08512_);
  and (_08514_, _08494_, _03083_);
  and (_08516_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  or (_08857_, _08516_, _08514_);
  and (_08517_, _08494_, _03087_);
  and (_08519_, _08496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  or (_08859_, _08519_, _08517_);
  and (_08520_, _08413_, _03136_);
  and (_08522_, _08520_, _03060_);
  not (_08523_, _08520_);
  and (_08524_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  or (_08863_, _08524_, _08522_);
  and (_08526_, _08520_, _03067_);
  and (_08527_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  or (_08867_, _08527_, _08526_);
  and (_08529_, _08520_, _03071_);
  and (_08530_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  or (_08870_, _08530_, _08529_);
  and (_08532_, _08520_, _03074_);
  and (_08533_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  or (_08873_, _08533_, _08532_);
  and (_08535_, _08520_, _03077_);
  and (_08537_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  or (_08877_, _08537_, _08535_);
  and (_08538_, _08520_, _03080_);
  and (_08539_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or (_08880_, _08539_, _08538_);
  and (_08541_, _08520_, _03083_);
  and (_08542_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  or (_08883_, _08542_, _08541_);
  and (_08544_, _08520_, _03087_);
  and (_08545_, _08523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or (_08886_, _08545_, _08544_);
  and (_08547_, _08413_, _03159_);
  and (_08548_, _08547_, _03060_);
  not (_08550_, _08547_);
  and (_08551_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_08890_, _08551_, _08548_);
  and (_08553_, _08547_, _03067_);
  and (_08554_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_08893_, _08554_, _08553_);
  and (_08556_, _08547_, _03071_);
  and (_08557_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_08896_, _08557_, _08556_);
  and (_08559_, _08547_, _03074_);
  and (_08560_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_08900_, _08560_, _08559_);
  and (_08562_, _08547_, _03077_);
  and (_08563_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_08904_, _08563_, _08562_);
  and (_08565_, _08547_, _03080_);
  and (_08566_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_08907_, _08566_, _08565_);
  and (_08568_, _08547_, _03083_);
  and (_08569_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_08911_, _08569_, _08568_);
  and (_08571_, _08547_, _03087_);
  and (_08572_, _08550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_08913_, _08572_, _08571_);
  and (_08574_, _08413_, _03179_);
  and (_08575_, _08574_, _03060_);
  not (_08576_, _08574_);
  and (_08578_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_08917_, _08578_, _08575_);
  and (_08579_, _08574_, _03067_);
  and (_08581_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_08920_, _08581_, _08579_);
  and (_08582_, _08574_, _03071_);
  and (_08584_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_08923_, _08584_, _08582_);
  and (_08586_, _08574_, _03074_);
  and (_08587_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_08926_, _08587_, _08586_);
  and (_08588_, _08574_, _03077_);
  and (_08590_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_08929_, _08590_, _08588_);
  and (_08591_, _08574_, _03080_);
  and (_08593_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_08933_, _08593_, _08591_);
  and (_08594_, _08574_, _03083_);
  and (_08596_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_08936_, _08596_, _08594_);
  and (_08597_, _08574_, _03087_);
  and (_08599_, _08576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_08938_, _08599_, _08597_);
  and (_08600_, _08413_, _03198_);
  and (_08602_, _08600_, _03060_);
  not (_08603_, _08600_);
  and (_08604_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  or (_08942_, _08604_, _08602_);
  and (_08606_, _08600_, _03067_);
  and (_08607_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  or (_08945_, _08607_, _08606_);
  and (_08609_, _08600_, _03071_);
  and (_08611_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  or (_08948_, _08611_, _08609_);
  and (_08612_, _08600_, _03074_);
  and (_08613_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  or (_08951_, _08613_, _08612_);
  and (_08615_, _08600_, _03077_);
  and (_08616_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  or (_08954_, _08616_, _08615_);
  and (_08618_, _08600_, _03080_);
  and (_08619_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  or (_08957_, _08619_, _08618_);
  and (_08621_, _08600_, _03083_);
  and (_08622_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  or (_08960_, _08622_, _08621_);
  and (_08624_, _08600_, _03087_);
  and (_08625_, _08603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  or (_08963_, _08625_, _08624_);
  and (_08627_, _08413_, _03218_);
  and (_08628_, _08627_, _03060_);
  not (_08630_, _08627_);
  and (_08631_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_08966_, _08631_, _08628_);
  and (_08633_, _08627_, _03067_);
  and (_08634_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_08969_, _08634_, _08633_);
  and (_08636_, _08627_, _03071_);
  and (_08637_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_08972_, _08637_, _08636_);
  and (_08639_, _08627_, _03074_);
  and (_08640_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_08975_, _08640_, _08639_);
  and (_08642_, _08627_, _03077_);
  and (_08643_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_08978_, _08643_, _08642_);
  and (_08645_, _08627_, _03080_);
  and (_08646_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_08981_, _08646_, _08645_);
  and (_08648_, _08627_, _03083_);
  and (_08649_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_08985_, _08649_, _08648_);
  and (_08651_, _08627_, _03087_);
  and (_08652_, _08630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_08987_, _08652_, _08651_);
  and (_08654_, _08413_, _03237_);
  and (_08655_, _08654_, _03060_);
  not (_08656_, _08654_);
  and (_08658_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  or (_08991_, _08658_, _08655_);
  and (_08660_, _08654_, _03067_);
  and (_08661_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  or (_08994_, _08661_, _08660_);
  and (_08662_, _08654_, _03071_);
  and (_08664_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  or (_08997_, _08664_, _08662_);
  and (_08665_, _08654_, _03074_);
  and (_08667_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  or (_09000_, _08667_, _08665_);
  and (_08668_, _08654_, _03077_);
  and (_08670_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  or (_09003_, _08670_, _08668_);
  and (_08671_, _08654_, _03080_);
  and (_08673_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or (_09006_, _08673_, _08671_);
  and (_08674_, _08654_, _03083_);
  and (_08676_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  or (_09009_, _08676_, _08674_);
  and (_08677_, _08654_, _03087_);
  and (_08679_, _08656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  or (_09012_, _08679_, _08677_);
  and (_08680_, _08413_, _03256_);
  and (_08682_, _08680_, _03060_);
  not (_08683_, _08680_);
  and (_08685_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  or (_09016_, _08685_, _08682_);
  and (_08686_, _08680_, _03067_);
  and (_08687_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  or (_09019_, _08687_, _08686_);
  and (_08689_, _08680_, _03071_);
  and (_08690_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  or (_09022_, _08690_, _08689_);
  and (_08692_, _08680_, _03074_);
  and (_08693_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  or (_09025_, _08693_, _08692_);
  and (_08695_, _08680_, _03077_);
  and (_08696_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  or (_09028_, _08696_, _08695_);
  and (_08698_, _08680_, _03080_);
  and (_08699_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  or (_09031_, _08699_, _08698_);
  and (_08701_, _08680_, _03083_);
  and (_08702_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  or (_09034_, _08702_, _08701_);
  and (_08704_, _08680_, _03087_);
  and (_08705_, _08683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  or (_09036_, _08705_, _08704_);
  and (_08707_, _08413_, _03275_);
  and (_08709_, _08707_, _03060_);
  not (_08710_, _08707_);
  and (_08711_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_09040_, _08711_, _08709_);
  and (_08713_, _08707_, _03067_);
  and (_08714_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_09043_, _08714_, _08713_);
  and (_08716_, _08707_, _03071_);
  and (_08717_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_09046_, _08717_, _08716_);
  and (_08719_, _08707_, _03074_);
  and (_08720_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_09049_, _08720_, _08719_);
  and (_08722_, _08707_, _03077_);
  and (_08723_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_09052_, _08723_, _08722_);
  and (_08725_, _08707_, _03080_);
  and (_08726_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_09055_, _08726_, _08725_);
  and (_08728_, _08707_, _03083_);
  and (_08729_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_09058_, _08729_, _08728_);
  and (_08731_, _08707_, _03087_);
  and (_08732_, _08710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_09061_, _08732_, _08731_);
  and (_08734_, _08413_, _03295_);
  and (_08735_, _08734_, _03060_);
  not (_08736_, _08734_);
  and (_08738_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_09065_, _08738_, _08735_);
  and (_08739_, _08734_, _03067_);
  and (_08741_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_09068_, _08741_, _08739_);
  and (_08742_, _08734_, _03071_);
  and (_08744_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_09071_, _08744_, _08742_);
  and (_08745_, _08734_, _03074_);
  and (_08747_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_09074_, _08747_, _08745_);
  and (_08748_, _08734_, _03077_);
  and (_08750_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_09077_, _08750_, _08748_);
  and (_08751_, _08734_, _03080_);
  and (_08753_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_09080_, _08753_, _08751_);
  and (_08754_, _08734_, _03083_);
  and (_08756_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_09083_, _08756_, _08754_);
  and (_08758_, _08734_, _03087_);
  and (_08759_, _08736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_09085_, _08759_, _08758_);
  and (_08760_, _08413_, _03315_);
  and (_08761_, _08760_, _03060_);
  not (_08763_, _08760_);
  and (_08764_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  or (_09089_, _08764_, _08761_);
  and (_08766_, _08760_, _03067_);
  and (_08767_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  or (_09093_, _08767_, _08766_);
  and (_08769_, _08760_, _03071_);
  and (_08770_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  or (_09096_, _08770_, _08769_);
  and (_08772_, _08760_, _03074_);
  and (_08773_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  or (_09099_, _08773_, _08772_);
  and (_08775_, _08760_, _03077_);
  and (_08776_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  or (_09102_, _08776_, _08775_);
  and (_08778_, _08760_, _03080_);
  and (_08779_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or (_09105_, _08779_, _08778_);
  and (_08781_, _08760_, _03083_);
  and (_08782_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  or (_09108_, _08782_, _08781_);
  and (_08784_, _08760_, _03087_);
  and (_08785_, _08763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  or (_09110_, _08785_, _08784_);
  and (_08787_, _08413_, _03334_);
  and (_08788_, _08787_, _03060_);
  not (_08789_, _08787_);
  and (_08791_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  or (_09114_, _08791_, _08788_);
  and (_08792_, _08787_, _03067_);
  and (_08794_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  or (_09117_, _08794_, _08792_);
  and (_08795_, _08787_, _03071_);
  and (_08797_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  or (_09120_, _08797_, _08795_);
  and (_08798_, _08787_, _03074_);
  and (_08800_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  or (_09123_, _08800_, _08798_);
  and (_08801_, _08787_, _03077_);
  and (_08803_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  or (_09126_, _08803_, _08801_);
  and (_08804_, _08787_, _03080_);
  and (_08806_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  or (_09129_, _08806_, _08804_);
  and (_08808_, _08787_, _03083_);
  and (_08809_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  or (_09132_, _08809_, _08808_);
  and (_08810_, _08787_, _03087_);
  and (_08812_, _08789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  or (_09135_, _08812_, _08810_);
  and (_08813_, _08413_, _03353_);
  and (_08815_, _08813_, _03060_);
  not (_08816_, _08813_);
  and (_08817_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_09138_, _08817_, _08815_);
  and (_08819_, _08813_, _03067_);
  and (_08820_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_09141_, _08820_, _08819_);
  and (_08822_, _08813_, _03071_);
  and (_08823_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_09145_, _08823_, _08822_);
  and (_08825_, _08813_, _03074_);
  and (_08826_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_09148_, _08826_, _08825_);
  and (_08828_, _08813_, _03077_);
  and (_08829_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_09151_, _08829_, _08828_);
  and (_08831_, _08813_, _03080_);
  and (_08833_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_09154_, _08833_, _08831_);
  and (_08834_, _08813_, _03083_);
  and (_08835_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_09157_, _08835_, _08834_);
  and (_08837_, _08813_, _03087_);
  and (_08838_, _08816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_09159_, _08838_, _08837_);
  and (_08840_, _03699_, _26939_);
  and (_08842_, _08840_, _02963_);
  and (_08844_, _08842_, _03060_);
  not (_08845_, _08842_);
  and (_08846_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_09164_, _08846_, _08844_);
  and (_08848_, _08842_, _03067_);
  and (_08849_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_09167_, _08849_, _08848_);
  and (_08851_, _08842_, _03071_);
  and (_08852_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_09170_, _08852_, _08851_);
  and (_08855_, _08842_, _03074_);
  and (_08856_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_09173_, _08856_, _08855_);
  and (_08858_, _08842_, _03077_);
  and (_08860_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_09176_, _08860_, _08858_);
  and (_08861_, _08842_, _03080_);
  and (_08862_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_09179_, _08862_, _08861_);
  and (_08865_, _08842_, _03083_);
  and (_08866_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_09182_, _08866_, _08865_);
  and (_08868_, _08842_, _03087_);
  and (_08869_, _08845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_09185_, _08869_, _08868_);
  and (_08871_, _08840_, _03062_);
  and (_08872_, _08871_, _03060_);
  not (_08874_, _08871_);
  and (_08875_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or (_09188_, _08875_, _08872_);
  and (_08878_, _08871_, _03067_);
  and (_08879_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or (_09191_, _08879_, _08878_);
  and (_08881_, _08871_, _03071_);
  and (_08882_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or (_09194_, _08882_, _08881_);
  and (_08884_, _08871_, _03074_);
  and (_08885_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or (_09198_, _08885_, _08884_);
  and (_08888_, _08871_, _03077_);
  and (_08889_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or (_09201_, _08889_, _08888_);
  and (_08891_, _08871_, _03080_);
  and (_08892_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or (_09204_, _08892_, _08891_);
  and (_08894_, _08871_, _03083_);
  and (_08895_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or (_09207_, _08895_, _08894_);
  and (_08897_, _08871_, _03087_);
  and (_08899_, _08874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or (_09209_, _08899_, _08897_);
  and (_08901_, _08840_, _03091_);
  and (_08902_, _08901_, _03060_);
  not (_08903_, _08901_);
  and (_08905_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or (_09213_, _08905_, _08902_);
  and (_08906_, _08901_, _03067_);
  and (_08908_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or (_09216_, _08908_, _08906_);
  and (_08910_, _08901_, _03071_);
  and (_08912_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or (_09219_, _08912_, _08910_);
  and (_08914_, _08901_, _03074_);
  and (_08915_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or (_09222_, _08915_, _08914_);
  and (_08916_, _08901_, _03077_);
  and (_08918_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or (_09226_, _08918_, _08916_);
  and (_08919_, _08901_, _03080_);
  and (_08921_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or (_09229_, _08921_, _08919_);
  and (_08922_, _08901_, _03083_);
  and (_08924_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or (_09232_, _08924_, _08922_);
  and (_08925_, _08901_, _03087_);
  and (_08927_, _08903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or (_09234_, _08927_, _08925_);
  and (_08928_, _08840_, _03113_);
  and (_08930_, _08928_, _03060_);
  not (_08931_, _08928_);
  and (_08932_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_09238_, _08932_, _08930_);
  and (_08934_, _08928_, _03067_);
  and (_08935_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_09241_, _08935_, _08934_);
  and (_08937_, _08928_, _03071_);
  and (_08939_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_09244_, _08939_, _08937_);
  and (_08940_, _08928_, _03074_);
  and (_08941_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_09247_, _08941_, _08940_);
  and (_08943_, _08928_, _03077_);
  and (_08944_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_09250_, _08944_, _08943_);
  and (_08946_, _08928_, _03080_);
  and (_08947_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_09253_, _08947_, _08946_);
  and (_08949_, _08928_, _03083_);
  and (_08950_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_09256_, _08950_, _08949_);
  and (_08952_, _08928_, _03087_);
  and (_08953_, _08931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_09259_, _08953_, _08952_);
  and (_08955_, _08840_, _03136_);
  and (_08956_, _08955_, _03060_);
  not (_08958_, _08955_);
  and (_08959_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_09262_, _08959_, _08956_);
  and (_08961_, _08955_, _03067_);
  and (_08962_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_09265_, _08962_, _08961_);
  and (_08964_, _08955_, _03071_);
  and (_08965_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_09268_, _08965_, _08964_);
  and (_08967_, _08955_, _03074_);
  and (_08968_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_09271_, _08968_, _08967_);
  and (_08970_, _08955_, _03077_);
  and (_08971_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_09274_, _08971_, _08970_);
  and (_08973_, _08955_, _03080_);
  and (_08974_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_09278_, _08974_, _08973_);
  and (_08976_, _08955_, _03083_);
  and (_08977_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_09281_, _08977_, _08976_);
  and (_08979_, _08955_, _03087_);
  and (_08980_, _08958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_09284_, _08980_, _08979_);
  and (_08982_, _08840_, _03159_);
  and (_08983_, _08982_, _03060_);
  not (_08984_, _08982_);
  and (_08986_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or (_09287_, _08986_, _08983_);
  and (_08988_, _08982_, _03067_);
  and (_08989_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or (_09290_, _08989_, _08988_);
  and (_08990_, _08982_, _03071_);
  and (_08992_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or (_09293_, _08992_, _08990_);
  and (_08993_, _08982_, _03074_);
  and (_08995_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or (_09296_, _08995_, _08993_);
  and (_08996_, _08982_, _03077_);
  and (_08998_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or (_09299_, _08998_, _08996_);
  and (_08999_, _08982_, _03080_);
  and (_09001_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or (_09302_, _09001_, _08999_);
  and (_09002_, _08982_, _03083_);
  and (_09004_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or (_09306_, _09004_, _09002_);
  and (_09005_, _08982_, _03087_);
  and (_09007_, _08984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or (_09308_, _09007_, _09005_);
  and (_09008_, _08840_, _03179_);
  and (_09010_, _09008_, _03060_);
  not (_09011_, _09008_);
  and (_09013_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or (_09312_, _09013_, _09010_);
  and (_09014_, _09008_, _03067_);
  and (_09015_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or (_09315_, _09015_, _09014_);
  and (_09017_, _09008_, _03071_);
  and (_09018_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or (_09318_, _09018_, _09017_);
  and (_09020_, _09008_, _03074_);
  and (_09021_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or (_09321_, _09021_, _09020_);
  and (_09023_, _09008_, _03077_);
  and (_09024_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or (_09324_, _09024_, _09023_);
  and (_09026_, _09008_, _03080_);
  and (_09027_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or (_09327_, _09027_, _09026_);
  and (_09029_, _09008_, _03083_);
  and (_09030_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or (_09330_, _09030_, _09029_);
  and (_09032_, _09008_, _03087_);
  and (_09033_, _09011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or (_09333_, _09033_, _09032_);
  and (_09035_, _08840_, _03198_);
  and (_09037_, _09035_, _03060_);
  not (_09038_, _09035_);
  and (_09039_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_09337_, _09039_, _09037_);
  and (_09041_, _09035_, _03067_);
  and (_09042_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_09340_, _09042_, _09041_);
  and (_09044_, _09035_, _03071_);
  and (_09045_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_09343_, _09045_, _09044_);
  and (_09047_, _09035_, _03074_);
  and (_09048_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_09346_, _09048_, _09047_);
  and (_09050_, _09035_, _03077_);
  and (_09051_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_09349_, _09051_, _09050_);
  and (_09053_, _09035_, _03080_);
  and (_09054_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_09352_, _09054_, _09053_);
  and (_09056_, _09035_, _03083_);
  and (_09057_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_09355_, _09057_, _09056_);
  and (_09059_, _09035_, _03087_);
  and (_09060_, _09038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_09357_, _09060_, _09059_);
  and (_09062_, _08840_, _03218_);
  and (_09063_, _09062_, _03060_);
  not (_09064_, _09062_);
  and (_09066_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or (_09361_, _09066_, _09063_);
  and (_09067_, _09062_, _03067_);
  and (_09069_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or (_09364_, _09069_, _09067_);
  and (_09070_, _09062_, _03071_);
  and (_09072_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or (_09367_, _09072_, _09070_);
  and (_09073_, _09062_, _03074_);
  and (_09075_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or (_09370_, _09075_, _09073_);
  and (_09076_, _09062_, _03077_);
  and (_09078_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or (_09373_, _09078_, _09076_);
  and (_09079_, _09062_, _03080_);
  and (_09081_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or (_09376_, _09081_, _09079_);
  and (_09082_, _09062_, _03083_);
  and (_09084_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or (_09379_, _09084_, _09082_);
  and (_09086_, _09062_, _03087_);
  and (_09087_, _09064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or (_09382_, _09087_, _09086_);
  and (_09088_, _08840_, _03237_);
  and (_09090_, _09088_, _03060_);
  not (_09091_, _09088_);
  and (_09092_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_09386_, _09092_, _09090_);
  and (_09094_, _09088_, _03067_);
  and (_09095_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_09389_, _09095_, _09094_);
  and (_09097_, _09088_, _03071_);
  and (_09098_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_09392_, _09098_, _09097_);
  and (_09100_, _09088_, _03074_);
  and (_09101_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_09395_, _09101_, _09100_);
  and (_09103_, _09088_, _03077_);
  and (_09104_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_09398_, _09104_, _09103_);
  and (_09106_, _09088_, _03080_);
  and (_09107_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_09401_, _09107_, _09106_);
  and (_09109_, _09088_, _03083_);
  and (_09111_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_09404_, _09111_, _09109_);
  and (_09112_, _09088_, _03087_);
  and (_09113_, _09091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_09406_, _09113_, _09112_);
  and (_09115_, _08840_, _03256_);
  and (_09116_, _09115_, _03060_);
  not (_09118_, _09115_);
  and (_09119_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_09410_, _09119_, _09116_);
  and (_09121_, _09115_, _03067_);
  and (_09122_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_09414_, _09122_, _09121_);
  and (_09124_, _09115_, _03071_);
  and (_09125_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_09417_, _09125_, _09124_);
  and (_09127_, _09115_, _03074_);
  and (_09128_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_09420_, _09128_, _09127_);
  and (_09130_, _09115_, _03077_);
  and (_09131_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_09423_, _09131_, _09130_);
  and (_09133_, _09115_, _03080_);
  and (_09134_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_09426_, _09134_, _09133_);
  and (_09136_, _09115_, _03083_);
  and (_09137_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_09429_, _09137_, _09136_);
  and (_09139_, _09115_, _03087_);
  and (_09140_, _09118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_09431_, _09140_, _09139_);
  and (_09142_, _08840_, _03275_);
  and (_09143_, _09142_, _03060_);
  not (_09144_, _09142_);
  and (_09146_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or (_09435_, _09146_, _09143_);
  and (_09147_, _09142_, _03067_);
  and (_09149_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or (_09438_, _09149_, _09147_);
  and (_09150_, _09142_, _03071_);
  and (_09152_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or (_09441_, _09152_, _09150_);
  and (_09153_, _09142_, _03074_);
  and (_09155_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or (_09444_, _09155_, _09153_);
  and (_09156_, _09142_, _03077_);
  and (_09158_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or (_09447_, _09158_, _09156_);
  and (_09160_, _09142_, _03080_);
  and (_09161_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or (_09450_, _09161_, _09160_);
  and (_09162_, _09142_, _03083_);
  and (_09163_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or (_09453_, _09163_, _09162_);
  and (_09165_, _09142_, _03087_);
  and (_09166_, _09144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or (_09456_, _09166_, _09165_);
  and (_09168_, _08840_, _03295_);
  and (_09169_, _09168_, _03060_);
  not (_09171_, _09168_);
  and (_09172_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or (_09459_, _09172_, _09169_);
  and (_09174_, _09168_, _03067_);
  and (_09175_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or (_09462_, _09175_, _09174_);
  and (_09177_, _09168_, _03071_);
  and (_09178_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or (_09466_, _09178_, _09177_);
  and (_09180_, _09168_, _03074_);
  and (_09181_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or (_09469_, _09181_, _09180_);
  and (_09183_, _09168_, _03077_);
  and (_09184_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or (_09472_, _09184_, _09183_);
  and (_09186_, _09168_, _03080_);
  and (_09187_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or (_09476_, _09187_, _09186_);
  and (_09189_, _09168_, _03083_);
  and (_09190_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or (_09479_, _09190_, _09189_);
  and (_09192_, _09168_, _03087_);
  and (_09193_, _09171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or (_09481_, _09193_, _09192_);
  and (_09195_, _08840_, _03315_);
  and (_09196_, _09195_, _03060_);
  not (_09197_, _09195_);
  and (_09199_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_09485_, _09199_, _09196_);
  and (_09200_, _09195_, _03067_);
  and (_09202_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_09488_, _09202_, _09200_);
  and (_09203_, _09195_, _03071_);
  and (_09205_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_09491_, _09205_, _09203_);
  and (_09206_, _09195_, _03074_);
  and (_09208_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_09495_, _09208_, _09206_);
  and (_09210_, _09195_, _03077_);
  and (_09211_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_09499_, _09211_, _09210_);
  and (_09212_, _09195_, _03080_);
  and (_09214_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_09502_, _09214_, _09212_);
  and (_09215_, _09195_, _03083_);
  and (_09217_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_09505_, _09217_, _09215_);
  and (_09218_, _09195_, _03087_);
  and (_09220_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_09507_, _09220_, _09218_);
  and (_09221_, _08840_, _03334_);
  and (_09223_, _09221_, _03060_);
  not (_09224_, _09221_);
  and (_09225_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_09511_, _09225_, _09223_);
  and (_09227_, _09221_, _03067_);
  and (_09228_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_09514_, _09228_, _09227_);
  and (_09230_, _09221_, _03071_);
  and (_09231_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_09517_, _09231_, _09230_);
  and (_09233_, _09221_, _03074_);
  and (_09235_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_09520_, _09235_, _09233_);
  and (_09236_, _09221_, _03077_);
  and (_09237_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_09523_, _09237_, _09236_);
  and (_09239_, _09221_, _03080_);
  and (_09240_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_09526_, _09240_, _09239_);
  and (_09242_, _09221_, _03083_);
  and (_09243_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_09529_, _09243_, _09242_);
  and (_09245_, _09221_, _03087_);
  and (_09246_, _09224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_09532_, _09246_, _09245_);
  and (_09248_, _08840_, _03353_);
  and (_09249_, _09248_, _03060_);
  not (_09251_, _09248_);
  and (_09252_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or (_09535_, _09252_, _09249_);
  and (_09254_, _09248_, _03067_);
  and (_09255_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or (_09538_, _09255_, _09254_);
  and (_09257_, _09248_, _03071_);
  and (_09258_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or (_09541_, _09258_, _09257_);
  and (_09260_, _09248_, _03074_);
  and (_09261_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or (_09544_, _09261_, _09260_);
  and (_09263_, _09248_, _03077_);
  and (_09264_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or (_09548_, _09264_, _09263_);
  and (_09266_, _09248_, _03080_);
  and (_09267_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or (_09551_, _09267_, _09266_);
  and (_09269_, _09248_, _03083_);
  and (_09270_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or (_09554_, _09270_, _09269_);
  and (_09272_, _09248_, _03087_);
  and (_09273_, _09251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or (_09556_, _09273_, _09272_);
  and (_09275_, _04125_, _26939_);
  and (_09276_, _09275_, _02963_);
  not (_09277_, _09276_);
  and (_09279_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_09280_, _09276_, _03060_);
  or (_09561_, _09280_, _09279_);
  and (_09282_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_09283_, _09276_, _03067_);
  or (_09564_, _09283_, _09282_);
  and (_09285_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_09286_, _09276_, _03071_);
  or (_09567_, _09286_, _09285_);
  and (_09288_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_09289_, _09276_, _03074_);
  or (_09570_, _09289_, _09288_);
  and (_09291_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_09292_, _09276_, _03077_);
  or (_09573_, _09292_, _09291_);
  and (_09294_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_09295_, _09276_, _03080_);
  or (_09576_, _09295_, _09294_);
  and (_09297_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_09298_, _09276_, _03083_);
  or (_09579_, _09298_, _09297_);
  and (_09300_, _09277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_09301_, _09276_, _03087_);
  or (_09582_, _09301_, _09300_);
  and (_09303_, _09275_, _03062_);
  not (_09304_, _09303_);
  and (_09305_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  and (_09307_, _09303_, _03060_);
  or (_09585_, _09307_, _09305_);
  and (_09309_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  and (_09310_, _09303_, _03067_);
  or (_09588_, _09310_, _09309_);
  and (_09311_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  and (_09313_, _09303_, _03071_);
  or (_09591_, _09313_, _09311_);
  and (_09314_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  and (_09316_, _09303_, _03074_);
  or (_09594_, _09316_, _09314_);
  and (_09317_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  and (_09319_, _09303_, _03077_);
  or (_09597_, _09319_, _09317_);
  and (_09320_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  and (_09322_, _09303_, _03080_);
  or (_09601_, _09322_, _09320_);
  and (_09323_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  and (_09325_, _09303_, _03083_);
  or (_09604_, _09325_, _09323_);
  and (_09326_, _09304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  and (_09328_, _09303_, _03087_);
  or (_09606_, _09328_, _09326_);
  and (_09329_, _09275_, _03091_);
  not (_09331_, _09329_);
  and (_09332_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  and (_09334_, _09329_, _03060_);
  or (_09610_, _09334_, _09332_);
  and (_09335_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  and (_09336_, _09329_, _03067_);
  or (_09613_, _09336_, _09335_);
  and (_09338_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  and (_09339_, _09329_, _03071_);
  or (_09616_, _09339_, _09338_);
  and (_09341_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  and (_09342_, _09329_, _03074_);
  or (_09619_, _09342_, _09341_);
  and (_09344_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and (_09345_, _09329_, _03077_);
  or (_09622_, _09345_, _09344_);
  and (_09347_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  and (_09348_, _09329_, _03080_);
  or (_09625_, _09348_, _09347_);
  and (_09350_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  and (_09351_, _09329_, _03083_);
  or (_09629_, _09351_, _09350_);
  and (_09353_, _09331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and (_09354_, _09329_, _03087_);
  or (_09631_, _09354_, _09353_);
  and (_09356_, _09275_, _03113_);
  not (_09358_, _09356_);
  and (_09359_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_09360_, _09356_, _03060_);
  or (_09635_, _09360_, _09359_);
  and (_09362_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_09363_, _09356_, _03067_);
  or (_09638_, _09363_, _09362_);
  and (_09365_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_09366_, _09356_, _03071_);
  or (_09641_, _09366_, _09365_);
  and (_09368_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_09369_, _09356_, _03074_);
  or (_09644_, _09369_, _09368_);
  and (_09371_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_09372_, _09356_, _03077_);
  or (_09647_, _09372_, _09371_);
  and (_09374_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_09375_, _09356_, _03080_);
  or (_09650_, _09375_, _09374_);
  and (_09377_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_09378_, _09356_, _03083_);
  or (_09653_, _09378_, _09377_);
  and (_09380_, _09358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_09381_, _09356_, _03087_);
  or (_09656_, _09381_, _09380_);
  and (_09383_, _09275_, _03136_);
  not (_09384_, _09383_);
  and (_09385_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_09387_, _09383_, _03060_);
  or (_09659_, _09387_, _09385_);
  and (_09388_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_09390_, _09383_, _03067_);
  or (_09662_, _09390_, _09388_);
  and (_09391_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_09393_, _09383_, _03071_);
  or (_09665_, _09393_, _09391_);
  and (_09394_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_09396_, _09383_, _03074_);
  or (_09668_, _09396_, _09394_);
  and (_09397_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_09399_, _09383_, _03077_);
  or (_09671_, _09399_, _09397_);
  and (_09400_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_09402_, _09383_, _03080_);
  or (_09674_, _09402_, _09400_);
  and (_09403_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_09405_, _09383_, _03083_);
  or (_09677_, _09405_, _09403_);
  and (_09407_, _09384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_09408_, _09383_, _03087_);
  or (_09680_, _09408_, _09407_);
  and (_09409_, _09275_, _03159_);
  not (_09411_, _09409_);
  and (_09412_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  and (_09413_, _09409_, _03060_);
  or (_09684_, _09413_, _09412_);
  and (_09415_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and (_09416_, _09409_, _03067_);
  or (_09687_, _09416_, _09415_);
  and (_09418_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  and (_09419_, _09409_, _03071_);
  or (_09690_, _09419_, _09418_);
  and (_09421_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and (_09422_, _09409_, _03074_);
  or (_09693_, _09422_, _09421_);
  and (_09424_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and (_09425_, _09409_, _03077_);
  or (_09696_, _09425_, _09424_);
  and (_09427_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and (_09428_, _09409_, _03080_);
  or (_09699_, _09428_, _09427_);
  and (_09430_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and (_09432_, _09409_, _03083_);
  or (_09702_, _09432_, _09430_);
  and (_09433_, _09411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and (_09434_, _09409_, _03087_);
  or (_09704_, _09434_, _09433_);
  and (_09436_, _09275_, _03179_);
  not (_09437_, _09436_);
  and (_09439_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  and (_09440_, _09436_, _03060_);
  or (_09709_, _09440_, _09439_);
  and (_09442_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  and (_09443_, _09436_, _03067_);
  or (_09713_, _09443_, _09442_);
  and (_09445_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and (_09446_, _09436_, _03071_);
  or (_09717_, _09446_, _09445_);
  and (_09448_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  and (_09449_, _09436_, _03074_);
  or (_09721_, _09449_, _09448_);
  and (_09451_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  and (_09452_, _09436_, _03077_);
  or (_09725_, _09452_, _09451_);
  and (_09454_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  and (_09455_, _09436_, _03080_);
  or (_09729_, _09455_, _09454_);
  and (_09457_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  and (_09458_, _09436_, _03083_);
  or (_09733_, _09458_, _09457_);
  and (_09460_, _09437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  and (_09461_, _09436_, _03087_);
  or (_09736_, _09461_, _09460_);
  and (_09463_, _09275_, _03198_);
  not (_09464_, _09463_);
  and (_09465_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_09467_, _09463_, _03060_);
  or (_09741_, _09467_, _09465_);
  and (_09468_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_09470_, _09463_, _03067_);
  or (_09745_, _09470_, _09468_);
  and (_09471_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_09473_, _09463_, _03071_);
  or (_09749_, _09473_, _09471_);
  and (_09475_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_09477_, _09463_, _03074_);
  or (_09753_, _09477_, _09475_);
  and (_09478_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_09480_, _09463_, _03077_);
  or (_09757_, _09480_, _09478_);
  and (_09482_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_09483_, _09463_, _03080_);
  or (_09761_, _09483_, _09482_);
  and (_09484_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_09486_, _09463_, _03083_);
  or (_09765_, _09486_, _09484_);
  and (_09487_, _09464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_09489_, _09463_, _03087_);
  or (_09768_, _09489_, _09487_);
  and (_09490_, _09275_, _03218_);
  not (_09492_, _09490_);
  and (_09493_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  and (_09494_, _09490_, _03060_);
  or (_09773_, _09494_, _09493_);
  and (_09497_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  and (_09498_, _09490_, _03067_);
  or (_09777_, _09498_, _09497_);
  and (_09500_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  and (_09501_, _09490_, _03071_);
  or (_09781_, _09501_, _09500_);
  and (_09503_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  and (_09504_, _09490_, _03074_);
  or (_09785_, _09504_, _09503_);
  and (_09506_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  and (_09508_, _09490_, _03077_);
  or (_09789_, _09508_, _09506_);
  and (_09509_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  and (_09510_, _09490_, _03080_);
  or (_09793_, _09510_, _09509_);
  and (_09512_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  and (_09513_, _09490_, _03083_);
  or (_09797_, _09513_, _09512_);
  and (_09515_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  and (_09516_, _09490_, _03087_);
  or (_09800_, _09516_, _09515_);
  and (_09518_, _09275_, _03237_);
  not (_09519_, _09518_);
  and (_09521_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_09522_, _09518_, _03060_);
  or (_09805_, _09522_, _09521_);
  and (_09524_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_09525_, _09518_, _03067_);
  or (_09809_, _09525_, _09524_);
  and (_09527_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_09528_, _09518_, _03071_);
  or (_09813_, _09528_, _09527_);
  and (_09530_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_09531_, _09518_, _03074_);
  or (_09817_, _09531_, _09530_);
  and (_09533_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_09534_, _09518_, _03077_);
  or (_09821_, _09534_, _09533_);
  and (_09536_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_09537_, _09518_, _03080_);
  or (_09825_, _09537_, _09536_);
  and (_09539_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_09540_, _09518_, _03083_);
  or (_09829_, _09540_, _09539_);
  and (_09542_, _09519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_09543_, _09518_, _03087_);
  or (_09832_, _09543_, _09542_);
  and (_09545_, _09275_, _03256_);
  not (_09546_, _09545_);
  and (_09547_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_09549_, _09545_, _03060_);
  or (_09837_, _09549_, _09547_);
  and (_09550_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_09552_, _09545_, _03067_);
  or (_09841_, _09552_, _09550_);
  and (_09553_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_09555_, _09545_, _03071_);
  or (_09845_, _09555_, _09553_);
  and (_09557_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_09558_, _09545_, _03074_);
  or (_09849_, _09558_, _09557_);
  and (_09559_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_09560_, _09545_, _03077_);
  or (_09853_, _09560_, _09559_);
  and (_09562_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_09563_, _09545_, _03080_);
  or (_09857_, _09563_, _09562_);
  and (_09565_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_09566_, _09545_, _03083_);
  or (_09861_, _09566_, _09565_);
  and (_09568_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_09569_, _09545_, _03087_);
  or (_09864_, _09569_, _09568_);
  and (_09571_, _09275_, _03275_);
  not (_09572_, _09571_);
  and (_09574_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  and (_09575_, _09571_, _03060_);
  or (_09869_, _09575_, _09574_);
  and (_09577_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  and (_09578_, _09571_, _03067_);
  or (_09873_, _09578_, _09577_);
  and (_09580_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  and (_09581_, _09571_, _03071_);
  or (_09877_, _09581_, _09580_);
  and (_09583_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and (_09584_, _09571_, _03074_);
  or (_09881_, _09584_, _09583_);
  and (_09586_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and (_09587_, _09571_, _03077_);
  or (_09885_, _09587_, _09586_);
  and (_09589_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  and (_09590_, _09571_, _03080_);
  or (_09889_, _09590_, _09589_);
  and (_09592_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  and (_09593_, _09571_, _03083_);
  or (_09893_, _09593_, _09592_);
  and (_09595_, _09572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  and (_09596_, _09571_, _03087_);
  or (_09896_, _09596_, _09595_);
  and (_09598_, _09275_, _03295_);
  not (_09599_, _09598_);
  and (_09600_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and (_09602_, _09598_, _03060_);
  or (_09901_, _09602_, _09600_);
  and (_09603_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  and (_09605_, _09598_, _03067_);
  or (_09905_, _09605_, _09603_);
  and (_09607_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  and (_09608_, _09598_, _03071_);
  or (_09909_, _09608_, _09607_);
  and (_09609_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  and (_09611_, _09598_, _03074_);
  or (_09913_, _09611_, _09609_);
  and (_09612_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  and (_09614_, _09598_, _03077_);
  or (_09917_, _09614_, _09612_);
  and (_09615_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  and (_09617_, _09598_, _03080_);
  or (_09921_, _09617_, _09615_);
  and (_09618_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  and (_09620_, _09598_, _03083_);
  or (_09925_, _09620_, _09618_);
  and (_09621_, _09599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  and (_09623_, _09598_, _03087_);
  or (_09928_, _09623_, _09621_);
  and (_09624_, _09275_, _03315_);
  not (_09626_, _09624_);
  and (_09627_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_09628_, _09624_, _03060_);
  or (_09933_, _09628_, _09627_);
  and (_09630_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_09632_, _09624_, _03067_);
  or (_09937_, _09632_, _09630_);
  and (_09633_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_09634_, _09624_, _03071_);
  or (_09941_, _09634_, _09633_);
  and (_09636_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_09637_, _09624_, _03074_);
  or (_09945_, _09637_, _09636_);
  and (_09639_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_09640_, _09624_, _03077_);
  or (_09949_, _09640_, _09639_);
  and (_09642_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_09643_, _09624_, _03080_);
  or (_09953_, _09643_, _09642_);
  and (_09645_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_09646_, _09624_, _03083_);
  or (_09957_, _09646_, _09645_);
  and (_09648_, _09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_09649_, _09624_, _03087_);
  or (_09960_, _09649_, _09648_);
  and (_09651_, _09275_, _03334_);
  not (_09652_, _09651_);
  and (_09654_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_09655_, _09651_, _03060_);
  or (_09965_, _09655_, _09654_);
  and (_09657_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_09658_, _09651_, _03067_);
  or (_09969_, _09658_, _09657_);
  and (_09660_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_09661_, _09651_, _03071_);
  or (_09973_, _09661_, _09660_);
  and (_09663_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_09664_, _09651_, _03074_);
  or (_09977_, _09664_, _09663_);
  and (_09666_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_09667_, _09651_, _03077_);
  or (_09981_, _09667_, _09666_);
  and (_09669_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_09670_, _09651_, _03080_);
  or (_09985_, _09670_, _09669_);
  and (_09672_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_09673_, _09651_, _03083_);
  or (_09989_, _09673_, _09672_);
  and (_09675_, _09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_09676_, _09651_, _03087_);
  or (_09992_, _09676_, _09675_);
  and (_09678_, _09275_, _03353_);
  not (_09679_, _09678_);
  and (_09681_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  and (_09682_, _09678_, _03060_);
  or (_09997_, _09682_, _09681_);
  and (_09683_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  and (_09685_, _09678_, _03067_);
  or (_10001_, _09685_, _09683_);
  and (_09686_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  and (_09688_, _09678_, _03071_);
  or (_10005_, _09688_, _09686_);
  and (_09689_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  and (_09691_, _09678_, _03074_);
  or (_10009_, _09691_, _09689_);
  and (_09692_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  and (_09694_, _09678_, _03077_);
  or (_10013_, _09694_, _09692_);
  and (_09695_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  and (_09697_, _09678_, _03080_);
  or (_10017_, _09697_, _09695_);
  and (_09698_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  and (_09700_, _09678_, _03083_);
  or (_10021_, _09700_, _09698_);
  and (_09701_, _09679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  and (_09703_, _09678_, _03087_);
  or (_10024_, _09703_, _09701_);
  and (_09705_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_09706_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_09707_, _09706_, _09705_);
  and (_09708_, _09707_, _01954_);
  and (_09710_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and (_09711_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_09712_, _09711_, _09710_);
  and (_09714_, _09712_, _02150_);
  or (_09715_, _09714_, _09708_);
  or (_09716_, _09715_, _02144_);
  and (_09718_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_09719_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_09720_, _09719_, _09718_);
  and (_09722_, _09720_, _01954_);
  and (_09723_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_09724_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_09726_, _09724_, _09723_);
  and (_09727_, _09726_, _02150_);
  or (_09728_, _09727_, _09722_);
  or (_09730_, _09728_, _02131_);
  and (_09731_, _09730_, _02157_);
  and (_09732_, _09731_, _09716_);
  or (_09734_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_09735_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and (_09737_, _09735_, _09734_);
  and (_09738_, _09737_, _01954_);
  or (_09739_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_09740_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_09742_, _09740_, _09739_);
  and (_09743_, _09742_, _02150_);
  or (_09744_, _09743_, _09738_);
  or (_09746_, _09744_, _02144_);
  or (_09747_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_09748_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_09750_, _09748_, _09747_);
  and (_09751_, _09750_, _01954_);
  or (_09752_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_09754_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and (_09755_, _09754_, _09752_);
  and (_09756_, _09755_, _02150_);
  or (_09758_, _09756_, _09751_);
  or (_09759_, _09758_, _02131_);
  and (_09760_, _09759_, _02077_);
  and (_09762_, _09760_, _09746_);
  or (_09763_, _09762_, _09732_);
  and (_09764_, _09763_, _02065_);
  and (_09766_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_09767_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_09769_, _09767_, _09766_);
  and (_09770_, _09769_, _01954_);
  and (_09771_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and (_09772_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_09774_, _09772_, _09771_);
  and (_09775_, _09774_, _02150_);
  or (_09776_, _09775_, _09770_);
  or (_09778_, _09776_, _02144_);
  and (_09779_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_09780_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_09782_, _09780_, _09779_);
  and (_09783_, _09782_, _01954_);
  and (_09784_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and (_09786_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_09787_, _09786_, _09784_);
  and (_09788_, _09787_, _02150_);
  or (_09790_, _09788_, _09783_);
  or (_09791_, _09790_, _02131_);
  and (_09792_, _09791_, _02157_);
  and (_09794_, _09792_, _09778_);
  or (_09795_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_09796_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and (_09798_, _09796_, _02150_);
  and (_09799_, _09798_, _09795_);
  or (_09801_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_09802_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_09803_, _09802_, _01954_);
  and (_09804_, _09803_, _09801_);
  or (_09806_, _09804_, _09799_);
  or (_09807_, _09806_, _02144_);
  or (_09808_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_09810_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_09811_, _09810_, _02150_);
  and (_09812_, _09811_, _09808_);
  or (_09814_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_09815_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_09816_, _09815_, _01954_);
  and (_09818_, _09816_, _09814_);
  or (_09819_, _09818_, _09812_);
  or (_09820_, _09819_, _02131_);
  and (_09822_, _09820_, _02077_);
  and (_09823_, _09822_, _09807_);
  or (_09824_, _09823_, _09794_);
  and (_09826_, _09824_, _02194_);
  or (_09827_, _09826_, _09764_);
  and (_09828_, _09827_, _02143_);
  and (_09830_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_09831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_09833_, _09831_, _09830_);
  and (_09834_, _09833_, _01954_);
  and (_09835_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_09836_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_09838_, _09836_, _09835_);
  and (_09839_, _09838_, _02150_);
  or (_09840_, _09839_, _09834_);
  and (_09842_, _09840_, _02131_);
  and (_09843_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_09844_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_09846_, _09844_, _09843_);
  and (_09847_, _09846_, _01954_);
  and (_09848_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_09850_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_09851_, _09850_, _09848_);
  and (_09852_, _09851_, _02150_);
  or (_09854_, _09852_, _09847_);
  and (_09855_, _09854_, _02144_);
  or (_09856_, _09855_, _09842_);
  and (_09858_, _09856_, _02157_);
  or (_09859_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_09860_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_09862_, _09860_, _02150_);
  and (_09863_, _09862_, _09859_);
  or (_09865_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_09866_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_09867_, _09866_, _01954_);
  and (_09868_, _09867_, _09865_);
  or (_09870_, _09868_, _09863_);
  and (_09871_, _09870_, _02131_);
  or (_09872_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_09874_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_09875_, _09874_, _02150_);
  and (_09876_, _09875_, _09872_);
  or (_09878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_09879_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_09880_, _09879_, _01954_);
  and (_09882_, _09880_, _09878_);
  or (_09883_, _09882_, _09876_);
  and (_09884_, _09883_, _02144_);
  or (_09886_, _09884_, _09871_);
  and (_09887_, _09886_, _02077_);
  or (_09888_, _09887_, _09858_);
  and (_09890_, _09888_, _02194_);
  and (_09891_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_09892_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_09894_, _09892_, _09891_);
  and (_09895_, _09894_, _01954_);
  and (_09897_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and (_09898_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_09899_, _09898_, _09897_);
  and (_09900_, _09899_, _02150_);
  or (_09902_, _09900_, _09895_);
  and (_09903_, _09902_, _02131_);
  and (_09904_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_09906_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_09907_, _09906_, _09904_);
  and (_09908_, _09907_, _01954_);
  and (_09910_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_09911_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_09912_, _09911_, _09910_);
  and (_09914_, _09912_, _02150_);
  or (_09915_, _09914_, _09908_);
  and (_09916_, _09915_, _02144_);
  or (_09918_, _09916_, _09903_);
  and (_09919_, _09918_, _02157_);
  or (_09920_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_09922_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_09923_, _09922_, _09920_);
  and (_09924_, _09923_, _01954_);
  or (_09926_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_09927_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_09929_, _09927_, _09926_);
  and (_09930_, _09929_, _02150_);
  or (_09931_, _09930_, _09924_);
  and (_09932_, _09931_, _02131_);
  or (_09934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_09935_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_09936_, _09935_, _09934_);
  and (_09938_, _09936_, _01954_);
  or (_09939_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_09940_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_09942_, _09940_, _09939_);
  and (_09943_, _09942_, _02150_);
  or (_09944_, _09943_, _09938_);
  and (_09946_, _09944_, _02144_);
  or (_09947_, _09946_, _09932_);
  and (_09948_, _09947_, _02077_);
  or (_09950_, _09948_, _09919_);
  and (_09951_, _09950_, _02065_);
  or (_09952_, _09951_, _09890_);
  and (_09954_, _09952_, _02005_);
  or (_09955_, _09954_, _09828_);
  or (_09956_, _09955_, _02054_);
  and (_09958_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_09959_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_09961_, _09959_, _09958_);
  and (_09962_, _09961_, _01954_);
  and (_09963_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_09964_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_09966_, _09964_, _09963_);
  and (_09967_, _09966_, _02150_);
  or (_09968_, _09967_, _09962_);
  or (_09970_, _09968_, _02144_);
  and (_09971_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_09972_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_09974_, _09972_, _09971_);
  and (_09975_, _09974_, _01954_);
  and (_09976_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_09978_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_09979_, _09978_, _09976_);
  and (_09980_, _09979_, _02150_);
  or (_09982_, _09980_, _09975_);
  or (_09983_, _09982_, _02131_);
  and (_09984_, _09983_, _02157_);
  and (_09986_, _09984_, _09970_);
  or (_09987_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_09988_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and (_09990_, _09988_, _02150_);
  and (_09991_, _09990_, _09987_);
  or (_09993_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_09994_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_09995_, _09994_, _01954_);
  and (_09996_, _09995_, _09993_);
  or (_09998_, _09996_, _09991_);
  or (_09999_, _09998_, _02144_);
  or (_10000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_10002_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_10003_, _10002_, _02150_);
  and (_10004_, _10003_, _10000_);
  or (_10006_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_10007_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_10008_, _10007_, _01954_);
  and (_10010_, _10008_, _10006_);
  or (_10011_, _10010_, _10004_);
  or (_10012_, _10011_, _02131_);
  and (_10014_, _10012_, _02077_);
  and (_10015_, _10014_, _09999_);
  or (_10016_, _10015_, _09986_);
  and (_10018_, _10016_, _02194_);
  and (_10019_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_10020_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_10022_, _10020_, _10019_);
  and (_10023_, _10022_, _01954_);
  and (_10025_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_10026_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_10027_, _10026_, _10025_);
  and (_10028_, _10027_, _02150_);
  or (_10029_, _10028_, _10023_);
  or (_10030_, _10029_, _02144_);
  and (_10031_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_10032_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_10033_, _10032_, _10031_);
  and (_10035_, _10033_, _01954_);
  and (_10036_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_10037_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_10039_, _10037_, _10036_);
  and (_10040_, _10039_, _02150_);
  or (_10041_, _10040_, _10035_);
  or (_10043_, _10041_, _02131_);
  and (_10044_, _10043_, _02157_);
  and (_10045_, _10044_, _10030_);
  or (_10047_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_10048_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_10049_, _10048_, _10047_);
  and (_10051_, _10049_, _01954_);
  or (_10052_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_10053_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_10055_, _10053_, _10052_);
  and (_10056_, _10055_, _02150_);
  or (_10057_, _10056_, _10051_);
  or (_10059_, _10057_, _02144_);
  or (_10060_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_10061_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_10062_, _10061_, _10060_);
  and (_10063_, _10062_, _01954_);
  or (_10064_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_10065_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_10066_, _10065_, _10064_);
  and (_10067_, _10066_, _02150_);
  or (_10068_, _10067_, _10063_);
  or (_10069_, _10068_, _02131_);
  and (_10070_, _10069_, _02077_);
  and (_10071_, _10070_, _10059_);
  or (_10072_, _10071_, _10045_);
  and (_10073_, _10072_, _02065_);
  or (_10074_, _10073_, _10018_);
  and (_10075_, _10074_, _02143_);
  or (_10076_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_10077_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_10078_, _10077_, _10076_);
  and (_10079_, _10078_, _01954_);
  or (_10080_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_10081_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_10082_, _10081_, _10080_);
  and (_10083_, _10082_, _02150_);
  or (_10084_, _10083_, _10079_);
  and (_10085_, _10084_, _02144_);
  or (_10086_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_10087_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_10088_, _10087_, _10086_);
  and (_10089_, _10088_, _01954_);
  or (_10090_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_10091_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_10092_, _10091_, _10090_);
  and (_10093_, _10092_, _02150_);
  or (_10094_, _10093_, _10089_);
  and (_10095_, _10094_, _02131_);
  or (_10096_, _10095_, _10085_);
  and (_10097_, _10096_, _02077_);
  and (_10098_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_10099_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_10100_, _10099_, _10098_);
  and (_10101_, _10100_, _01954_);
  and (_10102_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_10103_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_10104_, _10103_, _10102_);
  and (_10105_, _10104_, _02150_);
  or (_10106_, _10105_, _10101_);
  and (_10107_, _10106_, _02144_);
  and (_10108_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_10109_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_10110_, _10109_, _10108_);
  and (_10111_, _10110_, _01954_);
  and (_10112_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_10113_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_10114_, _10113_, _10112_);
  and (_10115_, _10114_, _02150_);
  or (_10116_, _10115_, _10111_);
  and (_10117_, _10116_, _02131_);
  or (_10118_, _10117_, _10107_);
  and (_10119_, _10118_, _02157_);
  or (_10120_, _10119_, _10097_);
  and (_10121_, _10120_, _02065_);
  or (_10122_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_10123_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and (_10124_, _10123_, _02150_);
  and (_10125_, _10124_, _10122_);
  or (_10126_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_10127_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and (_10128_, _10127_, _01954_);
  and (_10129_, _10128_, _10126_);
  or (_10130_, _10129_, _10125_);
  and (_10131_, _10130_, _02144_);
  or (_10132_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_10133_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and (_10134_, _10133_, _02150_);
  and (_10135_, _10134_, _10132_);
  or (_10136_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_10137_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and (_10138_, _10137_, _01954_);
  and (_10139_, _10138_, _10136_);
  or (_10140_, _10139_, _10135_);
  and (_10141_, _10140_, _02131_);
  or (_10142_, _10141_, _10131_);
  and (_10143_, _10142_, _02077_);
  and (_10144_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and (_10145_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_10146_, _10145_, _10144_);
  and (_10147_, _10146_, _01954_);
  and (_10148_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and (_10149_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_10150_, _10149_, _10148_);
  and (_10151_, _10150_, _02150_);
  or (_10152_, _10151_, _10147_);
  and (_10153_, _10152_, _02144_);
  and (_10154_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and (_10155_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_10156_, _10155_, _10154_);
  and (_10157_, _10156_, _01954_);
  and (_10158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_10159_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_10160_, _10159_, _10158_);
  and (_10161_, _10160_, _02150_);
  or (_10162_, _10161_, _10157_);
  and (_10163_, _10162_, _02131_);
  or (_10164_, _10163_, _10153_);
  and (_10165_, _10164_, _02157_);
  or (_10166_, _10165_, _10143_);
  and (_10167_, _10166_, _02194_);
  or (_10168_, _10167_, _10121_);
  and (_10169_, _10168_, _02005_);
  or (_10170_, _10169_, _10075_);
  or (_10171_, _10170_, _02374_);
  and (_10172_, _10171_, _09956_);
  or (_10173_, _10172_, _02142_);
  and (_10174_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_10175_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_10176_, _10175_, _10174_);
  and (_10177_, _10176_, _01954_);
  and (_10178_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_10179_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_10180_, _10179_, _10178_);
  and (_10181_, _10180_, _02150_);
  or (_10182_, _10181_, _10177_);
  and (_10183_, _10182_, _02131_);
  and (_10184_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_10185_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_10186_, _10185_, _10184_);
  and (_10187_, _10186_, _01954_);
  and (_10188_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_10189_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_10190_, _10189_, _10188_);
  and (_10191_, _10190_, _02150_);
  or (_10192_, _10191_, _10187_);
  and (_10193_, _10192_, _02144_);
  or (_10194_, _10193_, _10183_);
  and (_10195_, _10194_, _02157_);
  or (_10196_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_10197_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_10198_, _10197_, _02150_);
  and (_10199_, _10198_, _10196_);
  or (_10200_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_10201_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_10202_, _10201_, _01954_);
  and (_10203_, _10202_, _10200_);
  or (_10204_, _10203_, _10199_);
  and (_10205_, _10204_, _02131_);
  or (_10206_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_10207_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_10208_, _10207_, _02150_);
  and (_10209_, _10208_, _10206_);
  or (_10210_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_10211_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_10212_, _10211_, _01954_);
  and (_10213_, _10212_, _10210_);
  or (_10214_, _10213_, _10209_);
  and (_10215_, _10214_, _02144_);
  or (_10216_, _10215_, _10205_);
  and (_10217_, _10216_, _02077_);
  or (_10218_, _10217_, _10195_);
  and (_10219_, _10218_, _02194_);
  and (_10220_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_10221_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_10222_, _10221_, _10220_);
  and (_10223_, _10222_, _01954_);
  and (_10224_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_10225_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_10226_, _10225_, _10224_);
  and (_10227_, _10226_, _02150_);
  or (_10228_, _10227_, _10223_);
  and (_10229_, _10228_, _02131_);
  and (_10230_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_10231_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_10232_, _10231_, _10230_);
  and (_10233_, _10232_, _01954_);
  and (_10234_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_10235_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_10236_, _10235_, _10234_);
  and (_10237_, _10236_, _02150_);
  or (_10238_, _10237_, _10233_);
  and (_10239_, _10238_, _02144_);
  or (_10240_, _10239_, _10229_);
  and (_10241_, _10240_, _02157_);
  or (_10242_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_10243_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_10244_, _10243_, _10242_);
  and (_10245_, _10244_, _01954_);
  or (_10246_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_10247_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_10248_, _10247_, _10246_);
  and (_10249_, _10248_, _02150_);
  or (_10250_, _10249_, _10245_);
  and (_10251_, _10250_, _02131_);
  or (_10252_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_10253_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_10254_, _10253_, _10252_);
  and (_10255_, _10254_, _01954_);
  or (_10256_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_10257_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_10258_, _10257_, _10256_);
  and (_10259_, _10258_, _02150_);
  or (_10260_, _10259_, _10255_);
  and (_10261_, _10260_, _02144_);
  or (_10262_, _10261_, _10251_);
  and (_10263_, _10262_, _02077_);
  or (_10264_, _10263_, _10241_);
  and (_10265_, _10264_, _02065_);
  or (_10266_, _10265_, _10219_);
  and (_10267_, _10266_, _02005_);
  and (_10268_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_10269_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_10270_, _10269_, _10268_);
  and (_10271_, _10270_, _01954_);
  and (_10272_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_10273_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_10274_, _10273_, _10272_);
  and (_10275_, _10274_, _02150_);
  or (_10276_, _10275_, _10271_);
  or (_10277_, _10276_, _02144_);
  and (_10278_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_10279_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_10280_, _10279_, _10278_);
  and (_10281_, _10280_, _01954_);
  and (_10282_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_10283_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_10284_, _10283_, _10282_);
  and (_10285_, _10284_, _02150_);
  or (_10286_, _10285_, _10281_);
  or (_10287_, _10286_, _02131_);
  and (_10288_, _10287_, _02157_);
  and (_10289_, _10288_, _10277_);
  or (_10290_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_10291_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_10292_, _10291_, _10290_);
  and (_10293_, _10292_, _01954_);
  or (_10294_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_10295_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_10296_, _10295_, _10294_);
  and (_10297_, _10296_, _02150_);
  or (_10298_, _10297_, _10293_);
  or (_10299_, _10298_, _02144_);
  or (_10300_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_10301_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_10302_, _10301_, _10300_);
  and (_10303_, _10302_, _01954_);
  or (_10304_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_10305_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_10306_, _10305_, _10304_);
  and (_10307_, _10306_, _02150_);
  or (_10308_, _10307_, _10303_);
  or (_10309_, _10308_, _02131_);
  and (_10310_, _10309_, _02077_);
  and (_10311_, _10310_, _10299_);
  or (_10312_, _10311_, _10289_);
  and (_10313_, _10312_, _02065_);
  and (_10314_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_10315_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_10316_, _10315_, _10314_);
  and (_10317_, _10316_, _01954_);
  and (_10318_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_10319_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_10320_, _10319_, _10318_);
  and (_10321_, _10320_, _02150_);
  or (_10322_, _10321_, _10317_);
  or (_10323_, _10322_, _02144_);
  and (_10324_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_10325_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_10326_, _10325_, _10324_);
  and (_10327_, _10326_, _01954_);
  and (_10328_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_10329_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_10330_, _10329_, _10328_);
  and (_10331_, _10330_, _02150_);
  or (_10332_, _10331_, _10327_);
  or (_10333_, _10332_, _02131_);
  and (_10334_, _10333_, _02157_);
  and (_10335_, _10334_, _10323_);
  or (_10336_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_10337_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_10338_, _10337_, _02150_);
  and (_10339_, _10338_, _10336_);
  or (_10340_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_10341_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_10342_, _10341_, _01954_);
  and (_10343_, _10342_, _10340_);
  or (_10344_, _10343_, _10339_);
  or (_10345_, _10344_, _02144_);
  or (_10346_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_10347_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_10348_, _10347_, _02150_);
  and (_10349_, _10348_, _10346_);
  or (_10350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_10351_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_10352_, _10351_, _01954_);
  and (_10353_, _10352_, _10350_);
  or (_10354_, _10353_, _10349_);
  or (_10355_, _10354_, _02131_);
  and (_10356_, _10355_, _02077_);
  and (_10357_, _10356_, _10345_);
  or (_10358_, _10357_, _10335_);
  and (_10359_, _10358_, _02194_);
  or (_10360_, _10359_, _10313_);
  and (_10361_, _10360_, _02143_);
  or (_10362_, _10361_, _10267_);
  or (_10363_, _10362_, _02054_);
  and (_10364_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_10365_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_10366_, _10365_, _10364_);
  and (_10367_, _10366_, _02150_);
  and (_10368_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_10369_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_10370_, _10369_, _10368_);
  and (_10371_, _10370_, _01954_);
  or (_10372_, _10371_, _10367_);
  or (_10373_, _10372_, _02144_);
  and (_10374_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_10375_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_10376_, _10375_, _10374_);
  and (_10377_, _10376_, _02150_);
  and (_10378_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_10379_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_10380_, _10379_, _10378_);
  and (_10381_, _10380_, _01954_);
  or (_10382_, _10381_, _10377_);
  or (_10383_, _10382_, _02131_);
  and (_10384_, _10383_, _02157_);
  and (_10385_, _10384_, _10373_);
  or (_10386_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_10387_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_10388_, _10387_, _01954_);
  and (_10389_, _10388_, _10386_);
  or (_10390_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_10391_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_10392_, _10391_, _02150_);
  and (_10393_, _10392_, _10390_);
  or (_10394_, _10393_, _10389_);
  or (_10395_, _10394_, _02144_);
  or (_10396_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_10397_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_10398_, _10397_, _01954_);
  and (_10399_, _10398_, _10396_);
  or (_10400_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_10401_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_10402_, _10401_, _02150_);
  and (_10403_, _10402_, _10400_);
  or (_10404_, _10403_, _10399_);
  or (_10405_, _10404_, _02131_);
  and (_10406_, _10405_, _02077_);
  and (_10407_, _10406_, _10395_);
  or (_10408_, _10407_, _10385_);
  and (_10409_, _10408_, _02194_);
  and (_10410_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_10411_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_10412_, _10411_, _01954_);
  or (_10413_, _10412_, _10410_);
  and (_10414_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_10415_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_10416_, _10415_, _02150_);
  or (_10417_, _10416_, _10414_);
  and (_10418_, _10417_, _10413_);
  or (_10419_, _10418_, _02144_);
  and (_10420_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_10421_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_10422_, _10421_, _01954_);
  or (_10423_, _10422_, _10420_);
  and (_10424_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_10425_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_10426_, _10425_, _02150_);
  or (_10427_, _10426_, _10424_);
  and (_10428_, _10427_, _10423_);
  or (_10429_, _10428_, _02131_);
  and (_10430_, _10429_, _02157_);
  and (_10431_, _10430_, _10419_);
  or (_10432_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_10433_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_10434_, _10433_, _10432_);
  or (_10435_, _10434_, _02150_);
  or (_10436_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_10437_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_10438_, _10437_, _10436_);
  or (_10439_, _10438_, _01954_);
  and (_10440_, _10439_, _10435_);
  or (_10441_, _10440_, _02144_);
  or (_10442_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_10443_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_10444_, _10443_, _10442_);
  or (_10445_, _10444_, _02150_);
  or (_10446_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_10447_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_10448_, _10447_, _10446_);
  or (_10449_, _10448_, _01954_);
  and (_10450_, _10449_, _10445_);
  or (_10451_, _10450_, _02131_);
  and (_10452_, _10451_, _02077_);
  and (_10453_, _10452_, _10441_);
  or (_10454_, _10453_, _10431_);
  and (_10455_, _10454_, _02065_);
  or (_10456_, _10455_, _10409_);
  and (_10457_, _10456_, _02143_);
  and (_10458_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_10459_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_10460_, _10459_, _10458_);
  and (_10461_, _10460_, _01954_);
  and (_10462_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_10463_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_10464_, _10463_, _10462_);
  and (_10465_, _10464_, _02150_);
  or (_10466_, _10465_, _10461_);
  and (_10467_, _10466_, _02131_);
  and (_10468_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_10469_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_10470_, _10469_, _10468_);
  and (_10471_, _10470_, _01954_);
  and (_10472_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_10473_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_10474_, _10473_, _10472_);
  and (_10475_, _10474_, _02150_);
  or (_10476_, _10475_, _10471_);
  and (_10477_, _10476_, _02144_);
  or (_10478_, _10477_, _10467_);
  and (_10479_, _10478_, _02157_);
  or (_10480_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_10481_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_10482_, _10481_, _10480_);
  and (_10483_, _10482_, _01954_);
  or (_10484_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_10485_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_10486_, _10485_, _10484_);
  and (_10487_, _10486_, _02150_);
  or (_10488_, _10487_, _10483_);
  and (_10489_, _10488_, _02131_);
  or (_10490_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_10491_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_10492_, _10491_, _10490_);
  and (_10493_, _10492_, _01954_);
  or (_10494_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_10495_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_10496_, _10495_, _10494_);
  and (_10497_, _10496_, _02150_);
  or (_10498_, _10497_, _10493_);
  and (_10499_, _10498_, _02144_);
  or (_10500_, _10499_, _10489_);
  and (_10501_, _10500_, _02077_);
  or (_10502_, _10501_, _10479_);
  and (_10503_, _10502_, _02065_);
  and (_10504_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and (_10505_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or (_10506_, _10505_, _10504_);
  and (_10507_, _10506_, _01954_);
  and (_10508_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and (_10509_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_10510_, _10509_, _10508_);
  and (_10511_, _10510_, _02150_);
  or (_10512_, _10511_, _10507_);
  and (_10513_, _10512_, _02131_);
  and (_10514_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and (_10515_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or (_10516_, _10515_, _10514_);
  and (_10517_, _10516_, _01954_);
  and (_10518_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and (_10519_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_10520_, _10519_, _10518_);
  and (_10521_, _10520_, _02150_);
  or (_10522_, _10521_, _10517_);
  and (_10523_, _10522_, _02144_);
  or (_10524_, _10523_, _10513_);
  and (_10525_, _10524_, _02157_);
  or (_10526_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_10527_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and (_10528_, _10527_, _10526_);
  and (_10529_, _10528_, _01954_);
  or (_10530_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or (_10531_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and (_10532_, _10531_, _10530_);
  and (_10533_, _10532_, _02150_);
  or (_10534_, _10533_, _10529_);
  and (_10535_, _10534_, _02131_);
  or (_10536_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_10537_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and (_10538_, _10537_, _10536_);
  and (_10539_, _10538_, _01954_);
  or (_10540_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_10541_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and (_10542_, _10541_, _10540_);
  and (_10543_, _10542_, _02150_);
  or (_10544_, _10543_, _10539_);
  and (_10545_, _10544_, _02144_);
  or (_10546_, _10545_, _10535_);
  and (_10547_, _10546_, _02077_);
  or (_10548_, _10547_, _10525_);
  and (_10549_, _10548_, _02194_);
  or (_10550_, _10549_, _10503_);
  and (_10551_, _10550_, _02005_);
  or (_10552_, _10551_, _10457_);
  or (_10553_, _10552_, _02374_);
  and (_10554_, _10553_, _10363_);
  or (_10555_, _10554_, _01748_);
  and (_10556_, _10555_, _10173_);
  or (_10557_, _10556_, _02141_);
  or (_10558_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_10559_, _10558_, _27355_);
  and (_15236_, _10559_, _10557_);
  and (_10560_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_10561_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_10562_, _10561_, _10560_);
  and (_10563_, _10562_, _01954_);
  and (_10564_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_10565_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_10566_, _10565_, _10564_);
  and (_10567_, _10566_, _02150_);
  or (_10568_, _10567_, _10563_);
  or (_10569_, _10568_, _02144_);
  and (_10570_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_10571_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_10572_, _10571_, _10570_);
  and (_10573_, _10572_, _01954_);
  and (_10574_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and (_10575_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_10576_, _10575_, _10574_);
  and (_10577_, _10576_, _02150_);
  or (_10578_, _10577_, _10573_);
  or (_10579_, _10578_, _02131_);
  and (_10580_, _10579_, _02157_);
  and (_10581_, _10580_, _10569_);
  or (_10582_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_10583_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_10584_, _10583_, _10582_);
  and (_10585_, _10584_, _01954_);
  or (_10586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_10587_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_10588_, _10587_, _10586_);
  and (_10589_, _10588_, _02150_);
  or (_10590_, _10589_, _10585_);
  or (_10591_, _10590_, _02144_);
  or (_10592_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_10593_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and (_10594_, _10593_, _10592_);
  and (_10595_, _10594_, _01954_);
  or (_10596_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_10597_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_10598_, _10597_, _10596_);
  and (_10599_, _10598_, _02150_);
  or (_10600_, _10599_, _10595_);
  or (_10601_, _10600_, _02131_);
  and (_10602_, _10601_, _02077_);
  and (_10603_, _10602_, _10591_);
  or (_10604_, _10603_, _10581_);
  or (_10605_, _10604_, _02194_);
  and (_10606_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_10607_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_10608_, _10607_, _10606_);
  and (_10609_, _10608_, _01954_);
  and (_10610_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_10611_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_10612_, _10611_, _10610_);
  and (_10613_, _10612_, _02150_);
  or (_10614_, _10613_, _10609_);
  or (_10615_, _10614_, _02144_);
  and (_10616_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and (_10617_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_10618_, _10617_, _10616_);
  and (_10619_, _10618_, _01954_);
  and (_10620_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_10621_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_10622_, _10621_, _10620_);
  and (_10623_, _10622_, _02150_);
  or (_10624_, _10623_, _10619_);
  or (_10625_, _10624_, _02131_);
  and (_10626_, _10625_, _02157_);
  and (_10627_, _10626_, _10615_);
  or (_10628_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_10629_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and (_10630_, _10629_, _02150_);
  and (_10631_, _10630_, _10628_);
  or (_10632_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_10633_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_10634_, _10633_, _01954_);
  and (_10635_, _10634_, _10632_);
  or (_10636_, _10635_, _10631_);
  or (_10637_, _10636_, _02144_);
  or (_10638_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_10639_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and (_10640_, _10639_, _02150_);
  and (_10641_, _10640_, _10638_);
  or (_10642_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_10643_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_10644_, _10643_, _01954_);
  and (_10645_, _10644_, _10642_);
  or (_10646_, _10645_, _10641_);
  or (_10647_, _10646_, _02131_);
  and (_10648_, _10647_, _02077_);
  and (_10649_, _10648_, _10637_);
  or (_10650_, _10649_, _10627_);
  or (_10651_, _10650_, _02065_);
  and (_10652_, _10651_, _02143_);
  and (_10653_, _10652_, _10605_);
  and (_10654_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_10655_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_10656_, _10655_, _10654_);
  and (_10657_, _10656_, _01954_);
  and (_10658_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_10659_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_10660_, _10659_, _10658_);
  and (_10661_, _10660_, _02150_);
  or (_10662_, _10661_, _10657_);
  and (_10663_, _10662_, _02131_);
  and (_10664_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_10665_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_10666_, _10665_, _10664_);
  and (_10667_, _10666_, _01954_);
  and (_10668_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_10669_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_10670_, _10669_, _10668_);
  and (_10671_, _10670_, _02150_);
  or (_10672_, _10671_, _10667_);
  and (_10673_, _10672_, _02144_);
  or (_10674_, _10673_, _02077_);
  or (_10675_, _10674_, _10663_);
  or (_10676_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_10677_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_10678_, _10677_, _02150_);
  and (_10679_, _10678_, _10676_);
  or (_10680_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_10681_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_10682_, _10681_, _01954_);
  and (_10683_, _10682_, _10680_);
  or (_10684_, _10683_, _10679_);
  and (_10685_, _10684_, _02131_);
  or (_10686_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_10687_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_10688_, _10687_, _02150_);
  and (_10689_, _10688_, _10686_);
  or (_10690_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_10691_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_10692_, _10691_, _01954_);
  and (_10693_, _10692_, _10690_);
  or (_10694_, _10693_, _10689_);
  and (_10695_, _10694_, _02144_);
  or (_10696_, _10695_, _02157_);
  or (_10697_, _10696_, _10685_);
  and (_10698_, _10697_, _10675_);
  or (_10699_, _10698_, _02065_);
  and (_10700_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and (_10701_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_10702_, _10701_, _10700_);
  and (_10703_, _10702_, _01954_);
  and (_10704_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_10705_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_10706_, _10705_, _10704_);
  and (_10707_, _10706_, _02150_);
  or (_10708_, _10707_, _10703_);
  and (_10709_, _10708_, _02131_);
  and (_10710_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_10711_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_10712_, _10711_, _10710_);
  and (_10713_, _10712_, _01954_);
  and (_10714_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_10715_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_10716_, _10715_, _10714_);
  and (_10717_, _10716_, _02150_);
  or (_10719_, _10717_, _10713_);
  and (_10720_, _10719_, _02144_);
  or (_10721_, _10720_, _02077_);
  or (_10722_, _10721_, _10709_);
  or (_10723_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_10724_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and (_10725_, _10724_, _10723_);
  and (_10726_, _10725_, _01954_);
  or (_10727_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_10728_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_10730_, _10728_, _10727_);
  and (_10731_, _10730_, _02150_);
  or (_10732_, _10731_, _10726_);
  and (_10733_, _10732_, _02131_);
  or (_10734_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_10735_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_10736_, _10735_, _10734_);
  and (_10737_, _10736_, _01954_);
  or (_10738_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_10739_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_10741_, _10739_, _10738_);
  and (_10742_, _10741_, _02150_);
  or (_10743_, _10742_, _10737_);
  and (_10744_, _10743_, _02144_);
  or (_10745_, _10744_, _02157_);
  or (_10746_, _10745_, _10733_);
  and (_10747_, _10746_, _10722_);
  or (_10748_, _10747_, _02194_);
  and (_10749_, _10748_, _02005_);
  and (_10750_, _10749_, _10699_);
  or (_10752_, _10750_, _10653_);
  or (_10753_, _10752_, _02054_);
  and (_10754_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and (_10755_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_10756_, _10755_, _10754_);
  and (_10757_, _10756_, _01954_);
  and (_10758_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and (_10759_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_10760_, _10759_, _10758_);
  and (_10761_, _10760_, _02150_);
  or (_10763_, _10761_, _10757_);
  and (_10764_, _10763_, _02131_);
  and (_10765_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  and (_10766_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_10767_, _10766_, _10765_);
  and (_10768_, _10767_, _01954_);
  and (_10769_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and (_10770_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_10771_, _10770_, _10769_);
  and (_10772_, _10771_, _02150_);
  or (_10774_, _10772_, _10768_);
  and (_10775_, _10774_, _02144_);
  or (_10776_, _10775_, _02077_);
  or (_10777_, _10776_, _10764_);
  or (_10778_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_10779_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and (_10780_, _10779_, _10778_);
  and (_10781_, _10780_, _01954_);
  or (_10782_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_10783_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  and (_10785_, _10783_, _10782_);
  and (_10786_, _10785_, _02150_);
  or (_10787_, _10786_, _10781_);
  and (_10788_, _10787_, _02131_);
  or (_10789_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_10790_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  and (_10791_, _10790_, _10789_);
  and (_10792_, _10791_, _01954_);
  or (_10793_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_10794_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and (_10795_, _10794_, _10793_);
  and (_10796_, _10795_, _02150_);
  or (_10797_, _10796_, _10792_);
  and (_10798_, _10797_, _02144_);
  or (_10799_, _10798_, _02157_);
  or (_10800_, _10799_, _10788_);
  and (_10801_, _10800_, _10777_);
  or (_10802_, _10801_, _02065_);
  and (_10803_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_10804_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_10805_, _10804_, _10803_);
  and (_10806_, _10805_, _01954_);
  and (_10807_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and (_10808_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_10809_, _10808_, _10807_);
  and (_10810_, _10809_, _02150_);
  or (_10811_, _10810_, _10806_);
  and (_10812_, _10811_, _02131_);
  and (_10813_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_10814_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_10815_, _10814_, _10813_);
  and (_10816_, _10815_, _01954_);
  and (_10817_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and (_10818_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_10819_, _10818_, _10817_);
  and (_10820_, _10819_, _02150_);
  or (_10821_, _10820_, _10816_);
  and (_10822_, _10821_, _02144_);
  or (_10823_, _10822_, _02077_);
  or (_10824_, _10823_, _10812_);
  or (_10825_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_10826_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_10827_, _10826_, _10825_);
  and (_10828_, _10827_, _01954_);
  or (_10829_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_10830_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and (_10831_, _10830_, _10829_);
  and (_10832_, _10831_, _02150_);
  or (_10833_, _10832_, _10828_);
  and (_10834_, _10833_, _02131_);
  or (_10835_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_10836_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_10837_, _10836_, _10835_);
  and (_10838_, _10837_, _01954_);
  or (_10839_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_10840_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and (_10841_, _10840_, _10839_);
  and (_10842_, _10841_, _02150_);
  or (_10843_, _10842_, _10838_);
  and (_10844_, _10843_, _02144_);
  or (_10845_, _10844_, _02157_);
  or (_10846_, _10845_, _10834_);
  and (_10847_, _10846_, _10824_);
  or (_10848_, _10847_, _02194_);
  and (_10849_, _10848_, _02005_);
  and (_10850_, _10849_, _10802_);
  and (_10851_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_10852_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_10853_, _10852_, _10851_);
  and (_10854_, _10853_, _02150_);
  and (_10855_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and (_10856_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_10857_, _10856_, _10855_);
  and (_10858_, _10857_, _01954_);
  or (_10859_, _10858_, _10854_);
  or (_10860_, _10859_, _02144_);
  and (_10861_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_10862_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_10863_, _10862_, _10861_);
  and (_10864_, _10863_, _02150_);
  and (_10865_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and (_10866_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_10867_, _10866_, _10865_);
  and (_10868_, _10867_, _01954_);
  or (_10869_, _10868_, _10864_);
  or (_10870_, _10869_, _02131_);
  and (_10871_, _10870_, _02157_);
  and (_10872_, _10871_, _10860_);
  or (_10873_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_10874_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_10875_, _10874_, _01954_);
  and (_10876_, _10875_, _10873_);
  or (_10877_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_10878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_10879_, _10878_, _02150_);
  and (_10880_, _10879_, _10877_);
  or (_10881_, _10880_, _10876_);
  or (_10882_, _10881_, _02144_);
  or (_10883_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_10884_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and (_10885_, _10884_, _01954_);
  and (_10886_, _10885_, _10883_);
  or (_10887_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_10888_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_10889_, _10888_, _02150_);
  and (_10890_, _10889_, _10887_);
  or (_10891_, _10890_, _10886_);
  or (_10892_, _10891_, _02131_);
  and (_10893_, _10892_, _02077_);
  and (_10894_, _10893_, _10882_);
  or (_10895_, _10894_, _10872_);
  and (_10896_, _10895_, _02194_);
  and (_10897_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_10898_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_10899_, _10898_, _01954_);
  or (_10900_, _10899_, _10897_);
  and (_10901_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_10902_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_10903_, _10902_, _02150_);
  or (_10904_, _10903_, _10901_);
  and (_10905_, _10904_, _10900_);
  or (_10906_, _10905_, _02144_);
  and (_10907_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_10908_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_10909_, _10908_, _01954_);
  or (_10910_, _10909_, _10907_);
  and (_10911_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_10912_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_10913_, _10912_, _02150_);
  or (_10914_, _10913_, _10911_);
  and (_10915_, _10914_, _10910_);
  or (_10916_, _10915_, _02131_);
  and (_10917_, _10916_, _02157_);
  and (_10918_, _10917_, _10906_);
  or (_10919_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_10920_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_10921_, _10920_, _10919_);
  or (_10922_, _10921_, _02150_);
  or (_10923_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_10924_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_10925_, _10924_, _10923_);
  or (_10926_, _10925_, _01954_);
  and (_10927_, _10926_, _10922_);
  or (_10928_, _10927_, _02144_);
  or (_10929_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_10930_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_10931_, _10930_, _10929_);
  or (_10932_, _10931_, _02150_);
  or (_10933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_10934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_10935_, _10934_, _10933_);
  or (_10936_, _10935_, _01954_);
  and (_10937_, _10936_, _10932_);
  or (_10938_, _10937_, _02131_);
  and (_10939_, _10938_, _02077_);
  and (_10940_, _10939_, _10928_);
  or (_10941_, _10940_, _10918_);
  and (_10942_, _10941_, _02065_);
  or (_10943_, _10942_, _10896_);
  and (_10944_, _10943_, _02143_);
  or (_10945_, _10944_, _10850_);
  or (_10946_, _10945_, _02374_);
  and (_10947_, _10946_, _10753_);
  or (_10948_, _10947_, _02142_);
  and (_10949_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_10950_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_10951_, _10950_, _10949_);
  and (_10952_, _10951_, _01954_);
  and (_10953_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_10954_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_10955_, _10954_, _10953_);
  and (_10956_, _10955_, _02150_);
  or (_10957_, _10956_, _10952_);
  or (_10958_, _10957_, _02144_);
  and (_10959_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_10960_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_10961_, _10960_, _10959_);
  and (_10962_, _10961_, _01954_);
  and (_10963_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_10964_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_10965_, _10964_, _10963_);
  and (_10966_, _10965_, _02150_);
  or (_10967_, _10966_, _10962_);
  or (_10968_, _10967_, _02131_);
  and (_10969_, _10968_, _02157_);
  and (_10970_, _10969_, _10958_);
  or (_10971_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_10972_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_10973_, _10972_, _10971_);
  and (_10974_, _10973_, _01954_);
  or (_10975_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_10976_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_10977_, _10976_, _10975_);
  and (_10978_, _10977_, _02150_);
  or (_10979_, _10978_, _10974_);
  or (_10980_, _10979_, _02144_);
  or (_10981_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_10982_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_10983_, _10982_, _10981_);
  and (_10984_, _10983_, _01954_);
  or (_10985_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_10986_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_10987_, _10986_, _10985_);
  and (_10988_, _10987_, _02150_);
  or (_10989_, _10988_, _10984_);
  or (_10990_, _10989_, _02131_);
  and (_10991_, _10990_, _02077_);
  and (_10992_, _10991_, _10980_);
  or (_10993_, _10992_, _10970_);
  and (_10994_, _10993_, _02065_);
  and (_10995_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_10996_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_10997_, _10996_, _10995_);
  and (_10998_, _10997_, _01954_);
  and (_10999_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_11000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_11001_, _11000_, _10999_);
  and (_11002_, _11001_, _02150_);
  or (_11003_, _11002_, _10998_);
  or (_11004_, _11003_, _02144_);
  and (_11005_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_11006_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_11007_, _11006_, _11005_);
  and (_11008_, _11007_, _01954_);
  and (_11009_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_11010_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_11011_, _11010_, _11009_);
  and (_11012_, _11011_, _02150_);
  or (_11013_, _11012_, _11008_);
  or (_11014_, _11013_, _02131_);
  and (_11015_, _11014_, _02157_);
  and (_11016_, _11015_, _11004_);
  or (_11017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_11018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_11019_, _11018_, _02150_);
  and (_11020_, _11019_, _11017_);
  or (_11021_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_11022_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_11023_, _11022_, _01954_);
  and (_11024_, _11023_, _11021_);
  or (_11025_, _11024_, _11020_);
  or (_11026_, _11025_, _02144_);
  or (_11027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_11028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_11029_, _11028_, _02150_);
  and (_11030_, _11029_, _11027_);
  or (_11031_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_11032_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_11033_, _11032_, _01954_);
  and (_11034_, _11033_, _11031_);
  or (_11035_, _11034_, _11030_);
  or (_11036_, _11035_, _02131_);
  and (_11037_, _11036_, _02077_);
  and (_11038_, _11037_, _11026_);
  or (_11039_, _11038_, _11016_);
  and (_11040_, _11039_, _02194_);
  or (_11041_, _11040_, _10994_);
  and (_11042_, _11041_, _02143_);
  and (_11043_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and (_11044_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_11045_, _11044_, _11043_);
  and (_11046_, _11045_, _01954_);
  and (_11047_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_11048_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_11049_, _11048_, _11047_);
  and (_11050_, _11049_, _02150_);
  or (_11051_, _11050_, _11046_);
  and (_11052_, _11051_, _02131_);
  and (_11053_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_11054_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_11055_, _11054_, _11053_);
  and (_11056_, _11055_, _01954_);
  and (_11057_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_11058_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_11059_, _11058_, _11057_);
  and (_11060_, _11059_, _02150_);
  or (_11061_, _11060_, _11056_);
  and (_11062_, _11061_, _02144_);
  or (_11063_, _11062_, _11052_);
  and (_11064_, _11063_, _02157_);
  or (_11065_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_11066_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_11067_, _11066_, _02150_);
  and (_11068_, _11067_, _11065_);
  or (_11069_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_11070_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_11071_, _11070_, _01954_);
  and (_11072_, _11071_, _11069_);
  or (_11073_, _11072_, _11068_);
  and (_11074_, _11073_, _02131_);
  or (_11075_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_11076_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and (_11077_, _11076_, _02150_);
  and (_11078_, _11077_, _11075_);
  or (_11079_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_11080_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_11081_, _11080_, _01954_);
  and (_11082_, _11081_, _11079_);
  or (_11083_, _11082_, _11078_);
  and (_11084_, _11083_, _02144_);
  or (_11085_, _11084_, _11074_);
  and (_11086_, _11085_, _02077_);
  or (_11087_, _11086_, _11064_);
  and (_11088_, _11087_, _02194_);
  and (_11089_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_11090_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_11091_, _11090_, _11089_);
  and (_11092_, _11091_, _01954_);
  and (_11093_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_11094_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_11095_, _11094_, _11093_);
  and (_11096_, _11095_, _02150_);
  or (_11097_, _11096_, _11092_);
  and (_11098_, _11097_, _02131_);
  and (_11099_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_11100_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_11101_, _11100_, _11099_);
  and (_11102_, _11101_, _01954_);
  and (_11103_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_11104_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_11105_, _11104_, _11103_);
  and (_11106_, _11105_, _02150_);
  or (_11107_, _11106_, _11102_);
  and (_11108_, _11107_, _02144_);
  or (_11109_, _11108_, _11098_);
  and (_11110_, _11109_, _02157_);
  or (_11111_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_11112_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_11113_, _11112_, _11111_);
  and (_11114_, _11113_, _01954_);
  or (_11115_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_11116_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_11117_, _11116_, _11115_);
  and (_11118_, _11117_, _02150_);
  or (_11119_, _11118_, _11114_);
  and (_11120_, _11119_, _02131_);
  or (_11121_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_11122_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_11123_, _11122_, _11121_);
  and (_11124_, _11123_, _01954_);
  or (_11125_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_11126_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_11127_, _11126_, _11125_);
  and (_11128_, _11127_, _02150_);
  or (_11129_, _11128_, _11124_);
  and (_11130_, _11129_, _02144_);
  or (_11131_, _11130_, _11120_);
  and (_11132_, _11131_, _02077_);
  or (_11133_, _11132_, _11110_);
  and (_11134_, _11133_, _02065_);
  or (_11135_, _11134_, _11088_);
  and (_11136_, _11135_, _02005_);
  or (_11137_, _11136_, _11042_);
  or (_11138_, _11137_, _02054_);
  and (_11139_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_11140_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_11141_, _11140_, _11139_);
  and (_11142_, _11141_, _01954_);
  and (_11143_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_11144_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_11145_, _11144_, _11143_);
  and (_11146_, _11145_, _02150_);
  or (_11147_, _11146_, _11142_);
  or (_11148_, _11147_, _02144_);
  and (_11149_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_11150_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_11151_, _11150_, _11149_);
  and (_11152_, _11151_, _01954_);
  and (_11153_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_11154_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_11155_, _11154_, _11153_);
  and (_11156_, _11155_, _02150_);
  or (_11157_, _11156_, _11152_);
  or (_11158_, _11157_, _02131_);
  and (_11159_, _11158_, _02157_);
  and (_11160_, _11159_, _11148_);
  or (_11161_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_11162_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_11163_, _11162_, _02150_);
  and (_11164_, _11163_, _11161_);
  or (_11165_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_11166_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_11167_, _11166_, _01954_);
  and (_11168_, _11167_, _11165_);
  or (_11169_, _11168_, _11164_);
  or (_11170_, _11169_, _02144_);
  or (_11171_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_11172_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_11173_, _11172_, _02150_);
  and (_11174_, _11173_, _11171_);
  or (_11175_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_11176_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_11177_, _11176_, _01954_);
  and (_11178_, _11177_, _11175_);
  or (_11179_, _11178_, _11174_);
  or (_11180_, _11179_, _02131_);
  and (_11181_, _11180_, _02077_);
  and (_11182_, _11181_, _11170_);
  or (_11183_, _11182_, _11160_);
  and (_11184_, _11183_, _02194_);
  and (_11185_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_11186_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_11187_, _11186_, _11185_);
  and (_11188_, _11187_, _01954_);
  and (_11189_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_11190_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_11191_, _11190_, _11189_);
  and (_11192_, _11191_, _02150_);
  or (_11193_, _11192_, _11188_);
  or (_11194_, _11193_, _02144_);
  and (_11195_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_11196_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_11197_, _11196_, _11195_);
  and (_11198_, _11197_, _01954_);
  and (_11199_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_11200_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_11201_, _11200_, _11199_);
  and (_11202_, _11201_, _02150_);
  or (_11203_, _11202_, _11198_);
  or (_11204_, _11203_, _02131_);
  and (_11205_, _11204_, _02157_);
  and (_11206_, _11205_, _11194_);
  or (_11207_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_11208_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_11209_, _11208_, _11207_);
  and (_11210_, _11209_, _01954_);
  or (_11211_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_11212_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_11213_, _11212_, _11211_);
  and (_11214_, _11213_, _02150_);
  or (_11215_, _11214_, _11210_);
  or (_11216_, _11215_, _02144_);
  or (_11217_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_11218_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_11219_, _11218_, _11217_);
  and (_11220_, _11219_, _01954_);
  or (_11221_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_11222_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_11223_, _11222_, _11221_);
  and (_11224_, _11223_, _02150_);
  or (_11225_, _11224_, _11220_);
  or (_11226_, _11225_, _02131_);
  and (_11227_, _11226_, _02077_);
  and (_11228_, _11227_, _11216_);
  or (_11229_, _11228_, _11206_);
  and (_11230_, _11229_, _02065_);
  or (_11231_, _11230_, _11184_);
  and (_11232_, _11231_, _02143_);
  or (_11233_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_11234_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_11235_, _11234_, _11233_);
  and (_11236_, _11235_, _01954_);
  or (_11237_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_11238_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_11239_, _11238_, _11237_);
  and (_11240_, _11239_, _02150_);
  or (_11241_, _11240_, _11236_);
  and (_11242_, _11241_, _02144_);
  or (_11243_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_11244_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_11245_, _11244_, _11243_);
  and (_11246_, _11245_, _01954_);
  or (_11247_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_11248_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_11249_, _11248_, _11247_);
  and (_11250_, _11249_, _02150_);
  or (_11251_, _11250_, _11246_);
  and (_11252_, _11251_, _02131_);
  or (_11253_, _11252_, _11242_);
  and (_11254_, _11253_, _02077_);
  and (_11255_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_11256_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_11257_, _11256_, _11255_);
  and (_11258_, _11257_, _01954_);
  and (_11259_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_11260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_11261_, _11260_, _11259_);
  and (_11262_, _11261_, _02150_);
  or (_11263_, _11262_, _11258_);
  and (_11264_, _11263_, _02144_);
  and (_11265_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_11266_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_11267_, _11266_, _11265_);
  and (_11268_, _11267_, _01954_);
  and (_11269_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_11270_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_11271_, _11270_, _11269_);
  and (_11272_, _11271_, _02150_);
  or (_11273_, _11272_, _11268_);
  and (_11274_, _11273_, _02131_);
  or (_11275_, _11274_, _11264_);
  and (_11276_, _11275_, _02157_);
  or (_11277_, _11276_, _11254_);
  and (_11278_, _11277_, _02065_);
  or (_11279_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_11280_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_11281_, _11280_, _02150_);
  and (_11282_, _11281_, _11279_);
  or (_11283_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_11284_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_11285_, _11284_, _01954_);
  and (_11286_, _11285_, _11283_);
  or (_11287_, _11286_, _11282_);
  and (_11288_, _11287_, _02144_);
  or (_11289_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_11290_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_11291_, _11290_, _02150_);
  and (_11292_, _11291_, _11289_);
  or (_11293_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_11294_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_11295_, _11294_, _01954_);
  and (_11296_, _11295_, _11293_);
  or (_11297_, _11296_, _11292_);
  and (_11298_, _11297_, _02131_);
  or (_11299_, _11298_, _11288_);
  and (_11300_, _11299_, _02077_);
  and (_11301_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_11302_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_11303_, _11302_, _11301_);
  and (_11304_, _11303_, _01954_);
  and (_11305_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_11306_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_11307_, _11306_, _11305_);
  and (_11308_, _11307_, _02150_);
  or (_11309_, _11308_, _11304_);
  and (_11310_, _11309_, _02144_);
  and (_11311_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_11312_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_11313_, _11312_, _11311_);
  and (_11314_, _11313_, _01954_);
  and (_11315_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_11316_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_11317_, _11316_, _11315_);
  and (_11318_, _11317_, _02150_);
  or (_11319_, _11318_, _11314_);
  and (_11320_, _11319_, _02131_);
  or (_11321_, _11320_, _11310_);
  and (_11322_, _11321_, _02157_);
  or (_11323_, _11322_, _11300_);
  and (_11324_, _11323_, _02194_);
  or (_11325_, _11324_, _11278_);
  and (_11326_, _11325_, _02005_);
  or (_11327_, _11326_, _11232_);
  or (_11328_, _11327_, _02374_);
  and (_11329_, _11328_, _11138_);
  or (_11330_, _11329_, _01748_);
  and (_11331_, _11330_, _10948_);
  or (_11332_, _11331_, _02141_);
  or (_11333_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_11334_, _11333_, _27355_);
  and (_15238_, _11334_, _11332_);
  and (_11335_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_11336_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_11337_, _11336_, _11335_);
  and (_11338_, _11337_, _01954_);
  and (_11339_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_11340_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_11341_, _11340_, _11339_);
  and (_11342_, _11341_, _02150_);
  or (_11343_, _11342_, _11338_);
  or (_11344_, _11343_, _02144_);
  and (_11345_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_11346_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_11347_, _11346_, _11345_);
  and (_11348_, _11347_, _01954_);
  and (_11349_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_11350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_11351_, _11350_, _11349_);
  and (_11352_, _11351_, _02150_);
  or (_11353_, _11352_, _11348_);
  or (_11354_, _11353_, _02131_);
  and (_11355_, _11354_, _02157_);
  and (_11356_, _11355_, _11344_);
  or (_11357_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_11358_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_11359_, _11358_, _11357_);
  and (_11360_, _11359_, _01954_);
  or (_11361_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_11362_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_11363_, _11362_, _11361_);
  and (_11364_, _11363_, _02150_);
  or (_11365_, _11364_, _11360_);
  or (_11366_, _11365_, _02144_);
  or (_11367_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_11368_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_11369_, _11368_, _11367_);
  and (_11370_, _11369_, _01954_);
  or (_11371_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_11372_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_11373_, _11372_, _11371_);
  and (_11374_, _11373_, _02150_);
  or (_11375_, _11374_, _11370_);
  or (_11376_, _11375_, _02131_);
  and (_11377_, _11376_, _02077_);
  and (_11378_, _11377_, _11366_);
  or (_11379_, _11378_, _11356_);
  and (_11380_, _11379_, _02065_);
  and (_11381_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_11382_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_11383_, _11382_, _11381_);
  and (_11384_, _11383_, _01954_);
  and (_11385_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_11386_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_11387_, _11386_, _11385_);
  and (_11388_, _11387_, _02150_);
  or (_11389_, _11388_, _11384_);
  or (_11390_, _11389_, _02144_);
  and (_11391_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_11392_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_11393_, _11392_, _11391_);
  and (_11394_, _11393_, _01954_);
  and (_11395_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_11396_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_11397_, _11396_, _11395_);
  and (_11398_, _11397_, _02150_);
  or (_11399_, _11398_, _11394_);
  or (_11400_, _11399_, _02131_);
  and (_11401_, _11400_, _02157_);
  and (_11402_, _11401_, _11390_);
  or (_11403_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_11404_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and (_11405_, _11404_, _02150_);
  and (_11406_, _11405_, _11403_);
  or (_11407_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_11408_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and (_11409_, _11408_, _01954_);
  and (_11410_, _11409_, _11407_);
  or (_11411_, _11410_, _11406_);
  or (_11412_, _11411_, _02144_);
  or (_11413_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_11414_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_11415_, _11414_, _02150_);
  and (_11416_, _11415_, _11413_);
  or (_11417_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_11418_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_11419_, _11418_, _01954_);
  and (_11420_, _11419_, _11417_);
  or (_11421_, _11420_, _11416_);
  or (_11422_, _11421_, _02131_);
  and (_11423_, _11422_, _02077_);
  and (_11424_, _11423_, _11412_);
  or (_11425_, _11424_, _11402_);
  and (_11426_, _11425_, _02194_);
  or (_11427_, _11426_, _11380_);
  and (_11428_, _11427_, _02143_);
  and (_11429_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_11430_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_11431_, _11430_, _11429_);
  and (_11432_, _11431_, _01954_);
  and (_11433_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_11434_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_11435_, _11434_, _11433_);
  and (_11436_, _11435_, _02150_);
  or (_11437_, _11436_, _11432_);
  and (_11438_, _11437_, _02131_);
  and (_11439_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_11440_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_11441_, _11440_, _11439_);
  and (_11442_, _11441_, _01954_);
  and (_11443_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_11444_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_11445_, _11444_, _11443_);
  and (_11446_, _11445_, _02150_);
  or (_11447_, _11446_, _11442_);
  and (_11448_, _11447_, _02144_);
  or (_11449_, _11448_, _11438_);
  and (_11450_, _11449_, _02157_);
  or (_11451_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_11452_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_11453_, _11452_, _02150_);
  and (_11454_, _11453_, _11451_);
  or (_11455_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_11456_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_11457_, _11456_, _01954_);
  and (_11458_, _11457_, _11455_);
  or (_11459_, _11458_, _11454_);
  and (_11460_, _11459_, _02131_);
  or (_11461_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_11462_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_11463_, _11462_, _02150_);
  and (_11464_, _11463_, _11461_);
  or (_11465_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_11466_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_11467_, _11466_, _01954_);
  and (_11468_, _11467_, _11465_);
  or (_11469_, _11468_, _11464_);
  and (_11470_, _11469_, _02144_);
  or (_11471_, _11470_, _11460_);
  and (_11472_, _11471_, _02077_);
  or (_11473_, _11472_, _11450_);
  and (_11474_, _11473_, _02194_);
  and (_11475_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_11476_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_11477_, _11476_, _11475_);
  and (_11478_, _11477_, _01954_);
  and (_11479_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and (_11480_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_11481_, _11480_, _11479_);
  and (_11482_, _11481_, _02150_);
  or (_11483_, _11482_, _11478_);
  and (_11484_, _11483_, _02131_);
  and (_11485_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_11486_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_11487_, _11486_, _11485_);
  and (_11488_, _11487_, _01954_);
  and (_11489_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_11490_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_11491_, _11490_, _11489_);
  and (_11492_, _11491_, _02150_);
  or (_11493_, _11492_, _11488_);
  and (_11494_, _11493_, _02144_);
  or (_11495_, _11494_, _11484_);
  and (_11496_, _11495_, _02157_);
  or (_11497_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_11498_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_11499_, _11498_, _11497_);
  and (_11500_, _11499_, _01954_);
  or (_11501_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_11502_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_11503_, _11502_, _11501_);
  and (_11504_, _11503_, _02150_);
  or (_11505_, _11504_, _11500_);
  and (_11506_, _11505_, _02131_);
  or (_11507_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_11508_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_11509_, _11508_, _11507_);
  and (_11510_, _11509_, _01954_);
  or (_11511_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_11512_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_11513_, _11512_, _11511_);
  and (_11514_, _11513_, _02150_);
  or (_11515_, _11514_, _11510_);
  and (_11516_, _11515_, _02144_);
  or (_11517_, _11516_, _11506_);
  and (_11518_, _11517_, _02077_);
  or (_11519_, _11518_, _11496_);
  and (_11520_, _11519_, _02065_);
  or (_11521_, _11520_, _11474_);
  and (_11522_, _11521_, _02005_);
  or (_11523_, _11522_, _11428_);
  or (_11524_, _11523_, _02054_);
  and (_11525_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_11526_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_11527_, _11526_, _11525_);
  and (_11528_, _11527_, _01954_);
  and (_11529_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_11530_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_11531_, _11530_, _11529_);
  and (_11532_, _11531_, _02150_);
  or (_11533_, _11532_, _11528_);
  or (_11534_, _11533_, _02144_);
  and (_11535_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_11536_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_11537_, _11536_, _11535_);
  and (_11538_, _11537_, _01954_);
  and (_11539_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_11540_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_11541_, _11540_, _11539_);
  and (_11542_, _11541_, _02150_);
  or (_11543_, _11542_, _11538_);
  or (_11544_, _11543_, _02131_);
  and (_11545_, _11544_, _02157_);
  and (_11546_, _11545_, _11534_);
  or (_11547_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_11548_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_11549_, _11548_, _02150_);
  and (_11550_, _11549_, _11547_);
  or (_11551_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_11552_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_11553_, _11552_, _01954_);
  and (_11554_, _11553_, _11551_);
  or (_11555_, _11554_, _11550_);
  or (_11556_, _11555_, _02144_);
  or (_11557_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_11558_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_11559_, _11558_, _02150_);
  and (_11560_, _11559_, _11557_);
  or (_11561_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_11562_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and (_11563_, _11562_, _01954_);
  and (_11564_, _11563_, _11561_);
  or (_11565_, _11564_, _11560_);
  or (_11566_, _11565_, _02131_);
  and (_11567_, _11566_, _02077_);
  and (_11568_, _11567_, _11556_);
  or (_11569_, _11568_, _11546_);
  and (_11570_, _11569_, _02194_);
  and (_11571_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_11572_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_11573_, _11572_, _11571_);
  and (_11574_, _11573_, _01954_);
  and (_11575_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_11576_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_11577_, _11576_, _11575_);
  and (_11578_, _11577_, _02150_);
  or (_11579_, _11578_, _11574_);
  or (_11580_, _11579_, _02144_);
  and (_11581_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_11582_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_11583_, _11582_, _11581_);
  and (_11584_, _11583_, _01954_);
  and (_11585_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_11586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_11587_, _11586_, _11585_);
  and (_11588_, _11587_, _02150_);
  or (_11589_, _11588_, _11584_);
  or (_11590_, _11589_, _02131_);
  and (_11591_, _11590_, _02157_);
  and (_11592_, _11591_, _11580_);
  or (_11593_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_11594_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_11595_, _11594_, _11593_);
  and (_11596_, _11595_, _01954_);
  or (_11597_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_11598_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_11599_, _11598_, _11597_);
  and (_11600_, _11599_, _02150_);
  or (_11601_, _11600_, _11596_);
  or (_11602_, _11601_, _02144_);
  or (_11603_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_11604_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_11605_, _11604_, _11603_);
  and (_11606_, _11605_, _01954_);
  or (_11607_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_11608_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_11609_, _11608_, _11607_);
  and (_11610_, _11609_, _02150_);
  or (_11611_, _11610_, _11606_);
  or (_11612_, _11611_, _02131_);
  and (_11613_, _11612_, _02077_);
  and (_11614_, _11613_, _11602_);
  or (_11615_, _11614_, _11592_);
  and (_11616_, _11615_, _02065_);
  or (_11617_, _11616_, _11570_);
  and (_11618_, _11617_, _02143_);
  or (_11619_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_11620_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_11621_, _11620_, _11619_);
  and (_11622_, _11621_, _01954_);
  or (_11623_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_11624_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and (_11625_, _11624_, _11623_);
  and (_11626_, _11625_, _02150_);
  or (_11627_, _11626_, _11622_);
  and (_11628_, _11627_, _02144_);
  or (_11629_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_11630_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_11631_, _11630_, _11629_);
  and (_11632_, _11631_, _01954_);
  or (_11633_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_11634_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_11635_, _11634_, _11633_);
  and (_11636_, _11635_, _02150_);
  or (_11637_, _11636_, _11632_);
  and (_11638_, _11637_, _02131_);
  or (_11639_, _11638_, _11628_);
  and (_11640_, _11639_, _02077_);
  and (_11641_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_11642_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_11643_, _11642_, _11641_);
  and (_11644_, _11643_, _01954_);
  and (_11645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_11646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_11647_, _11646_, _11645_);
  and (_11648_, _11647_, _02150_);
  or (_11649_, _11648_, _11644_);
  and (_11650_, _11649_, _02144_);
  and (_11651_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_11652_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_11653_, _11652_, _11651_);
  and (_11654_, _11653_, _01954_);
  and (_11655_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_11656_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_11657_, _11656_, _11655_);
  and (_11658_, _11657_, _02150_);
  or (_11659_, _11658_, _11654_);
  and (_11660_, _11659_, _02131_);
  or (_11661_, _11660_, _11650_);
  and (_11662_, _11661_, _02157_);
  or (_11663_, _11662_, _11640_);
  and (_11664_, _11663_, _02065_);
  or (_11665_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_11666_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and (_11667_, _11666_, _02150_);
  and (_11668_, _11667_, _11665_);
  or (_11669_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_11670_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_11671_, _11670_, _01954_);
  and (_11672_, _11671_, _11669_);
  or (_11673_, _11672_, _11668_);
  and (_11674_, _11673_, _02144_);
  or (_11675_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_11676_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and (_11677_, _11676_, _02150_);
  and (_11678_, _11677_, _11675_);
  or (_11679_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_11680_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_11681_, _11680_, _01954_);
  and (_11682_, _11681_, _11679_);
  or (_11683_, _11682_, _11678_);
  and (_11684_, _11683_, _02131_);
  or (_11685_, _11684_, _11674_);
  and (_11686_, _11685_, _02077_);
  and (_11687_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_11688_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_11689_, _11688_, _11687_);
  and (_11690_, _11689_, _01954_);
  and (_11691_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and (_11692_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_11693_, _11692_, _11691_);
  and (_11694_, _11693_, _02150_);
  or (_11695_, _11694_, _11690_);
  and (_11696_, _11695_, _02144_);
  and (_11697_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and (_11698_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_11699_, _11698_, _11697_);
  and (_11700_, _11699_, _01954_);
  and (_11701_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_11702_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_11703_, _11702_, _11701_);
  and (_11704_, _11703_, _02150_);
  or (_11705_, _11704_, _11700_);
  and (_11706_, _11705_, _02131_);
  or (_11707_, _11706_, _11696_);
  and (_11708_, _11707_, _02157_);
  or (_11709_, _11708_, _11686_);
  and (_11710_, _11709_, _02194_);
  or (_11711_, _11710_, _11664_);
  and (_11712_, _11711_, _02005_);
  or (_11713_, _11712_, _11618_);
  or (_11714_, _11713_, _02374_);
  and (_11715_, _11714_, _11524_);
  or (_11716_, _11715_, _02142_);
  and (_11717_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_11718_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_11719_, _11718_, _11717_);
  and (_11720_, _11719_, _01954_);
  and (_11721_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_11722_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_11723_, _11722_, _11721_);
  and (_11724_, _11723_, _02150_);
  or (_11725_, _11724_, _11720_);
  or (_11726_, _11725_, _02144_);
  and (_11727_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_11728_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_11729_, _11728_, _11727_);
  and (_11730_, _11729_, _01954_);
  and (_11731_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_11732_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_11733_, _11732_, _11731_);
  and (_11734_, _11733_, _02150_);
  or (_11735_, _11734_, _11730_);
  or (_11736_, _11735_, _02131_);
  and (_11737_, _11736_, _02157_);
  and (_11738_, _11737_, _11726_);
  or (_11739_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_11740_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_11741_, _11740_, _11739_);
  and (_11742_, _11741_, _01954_);
  or (_11743_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_11744_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_11745_, _11744_, _11743_);
  and (_11746_, _11745_, _02150_);
  or (_11747_, _11746_, _11742_);
  or (_11748_, _11747_, _02144_);
  or (_11749_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_11750_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_11751_, _11750_, _11749_);
  and (_11752_, _11751_, _01954_);
  or (_11753_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_11754_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_11755_, _11754_, _11753_);
  and (_11756_, _11755_, _02150_);
  or (_11757_, _11756_, _11752_);
  or (_11758_, _11757_, _02131_);
  and (_11759_, _11758_, _02077_);
  and (_11760_, _11759_, _11748_);
  or (_11761_, _11760_, _11738_);
  and (_11762_, _11761_, _02065_);
  and (_11763_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_11764_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_11765_, _11764_, _11763_);
  and (_11766_, _11765_, _01954_);
  and (_11767_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_11768_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_11769_, _11768_, _11767_);
  and (_11770_, _11769_, _02150_);
  or (_11771_, _11770_, _11766_);
  or (_11772_, _11771_, _02144_);
  and (_11773_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_11774_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_11775_, _11774_, _11773_);
  and (_11776_, _11775_, _01954_);
  and (_11777_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_11778_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_11779_, _11778_, _11777_);
  and (_11780_, _11779_, _02150_);
  or (_11781_, _11780_, _11776_);
  or (_11782_, _11781_, _02131_);
  and (_11783_, _11782_, _02157_);
  and (_11784_, _11783_, _11772_);
  or (_11785_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_11786_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_11787_, _11786_, _02150_);
  and (_11788_, _11787_, _11785_);
  or (_11789_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_11790_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_11791_, _11790_, _01954_);
  and (_11792_, _11791_, _11789_);
  or (_11793_, _11792_, _11788_);
  or (_11794_, _11793_, _02144_);
  or (_11795_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_11796_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_11797_, _11796_, _02150_);
  and (_11798_, _11797_, _11795_);
  or (_11799_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_11800_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_11801_, _11800_, _01954_);
  and (_11802_, _11801_, _11799_);
  or (_11803_, _11802_, _11798_);
  or (_11804_, _11803_, _02131_);
  and (_11805_, _11804_, _02077_);
  and (_11806_, _11805_, _11794_);
  or (_11807_, _11806_, _11784_);
  and (_11808_, _11807_, _02194_);
  or (_11809_, _11808_, _11762_);
  and (_11810_, _11809_, _02143_);
  and (_11811_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_11812_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_11813_, _11812_, _11811_);
  and (_11814_, _11813_, _01954_);
  and (_11815_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_11816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_11817_, _11816_, _11815_);
  and (_11818_, _11817_, _02150_);
  or (_11819_, _11818_, _11814_);
  and (_11820_, _11819_, _02131_);
  and (_11821_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and (_11822_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_11823_, _11822_, _11821_);
  and (_11824_, _11823_, _01954_);
  and (_11825_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_11826_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_11827_, _11826_, _11825_);
  and (_11828_, _11827_, _02150_);
  or (_11829_, _11828_, _11824_);
  and (_11830_, _11829_, _02144_);
  or (_11831_, _11830_, _11820_);
  and (_11832_, _11831_, _02157_);
  or (_11833_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_11834_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and (_11835_, _11834_, _02150_);
  and (_11836_, _11835_, _11833_);
  or (_11837_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_11838_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and (_11839_, _11838_, _01954_);
  and (_11840_, _11839_, _11837_);
  or (_11841_, _11840_, _11836_);
  and (_11842_, _11841_, _02131_);
  or (_11843_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_11844_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and (_11845_, _11844_, _02150_);
  and (_11846_, _11845_, _11843_);
  or (_11847_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_11848_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_11849_, _11848_, _01954_);
  and (_11850_, _11849_, _11847_);
  or (_11851_, _11850_, _11846_);
  and (_11852_, _11851_, _02144_);
  or (_11853_, _11852_, _11842_);
  and (_11854_, _11853_, _02077_);
  or (_11855_, _11854_, _11832_);
  and (_11856_, _11855_, _02194_);
  and (_11857_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_11858_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_11859_, _11858_, _11857_);
  and (_11860_, _11859_, _01954_);
  and (_11861_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_11862_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_11863_, _11862_, _11861_);
  and (_11864_, _11863_, _02150_);
  or (_11865_, _11864_, _11860_);
  and (_11866_, _11865_, _02131_);
  and (_11867_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_11868_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_11869_, _11868_, _11867_);
  and (_11870_, _11869_, _01954_);
  and (_11871_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_11872_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_11873_, _11872_, _11871_);
  and (_11874_, _11873_, _02150_);
  or (_11875_, _11874_, _11870_);
  and (_11876_, _11875_, _02144_);
  or (_11877_, _11876_, _11866_);
  and (_11878_, _11877_, _02157_);
  or (_11879_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_11880_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_11881_, _11880_, _11879_);
  and (_11882_, _11881_, _01954_);
  or (_11883_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_11884_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_11885_, _11884_, _11883_);
  and (_11886_, _11885_, _02150_);
  or (_11887_, _11886_, _11882_);
  and (_11888_, _11887_, _02131_);
  or (_11889_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_11890_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_11891_, _11890_, _11889_);
  and (_11892_, _11891_, _01954_);
  or (_11893_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_11894_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_11895_, _11894_, _11893_);
  and (_11896_, _11895_, _02150_);
  or (_11897_, _11896_, _11892_);
  and (_11898_, _11897_, _02144_);
  or (_11899_, _11898_, _11888_);
  and (_11900_, _11899_, _02077_);
  or (_11901_, _11900_, _11878_);
  and (_11902_, _11901_, _02065_);
  or (_11903_, _11902_, _11856_);
  and (_11904_, _11903_, _02005_);
  or (_11905_, _11904_, _11810_);
  or (_11906_, _11905_, _02054_);
  and (_11907_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_11908_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_11909_, _11908_, _11907_);
  and (_11910_, _11909_, _01954_);
  and (_11911_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_11912_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_11913_, _11912_, _11911_);
  and (_11914_, _11913_, _02150_);
  or (_11915_, _11914_, _11910_);
  or (_11916_, _11915_, _02144_);
  and (_11917_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_11918_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_11919_, _11918_, _11917_);
  and (_11920_, _11919_, _01954_);
  and (_11921_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_11922_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_11923_, _11922_, _11921_);
  and (_11924_, _11923_, _02150_);
  or (_11925_, _11924_, _11920_);
  or (_11926_, _11925_, _02131_);
  and (_11927_, _11926_, _02157_);
  and (_11928_, _11927_, _11916_);
  or (_11929_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_11930_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_11931_, _11930_, _02150_);
  and (_11932_, _11931_, _11929_);
  or (_11933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_11934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_11935_, _11934_, _01954_);
  and (_11936_, _11935_, _11933_);
  or (_11937_, _11936_, _11932_);
  or (_11938_, _11937_, _02144_);
  or (_11939_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_11940_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_11941_, _11940_, _02150_);
  and (_11942_, _11941_, _11939_);
  or (_11943_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_11944_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_11945_, _11944_, _01954_);
  and (_11946_, _11945_, _11943_);
  or (_11947_, _11946_, _11942_);
  or (_11948_, _11947_, _02131_);
  and (_11949_, _11948_, _02077_);
  and (_11950_, _11949_, _11938_);
  or (_11951_, _11950_, _11928_);
  and (_11952_, _11951_, _02194_);
  and (_11953_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_11954_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_11955_, _11954_, _11953_);
  and (_11956_, _11955_, _01954_);
  and (_11957_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_11958_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_11959_, _11958_, _11957_);
  and (_11960_, _11959_, _02150_);
  or (_11961_, _11960_, _11956_);
  or (_11962_, _11961_, _02144_);
  and (_11963_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_11964_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_11965_, _11964_, _11963_);
  and (_11966_, _11965_, _01954_);
  and (_11967_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_11968_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_11969_, _11968_, _11967_);
  and (_11970_, _11969_, _02150_);
  or (_11971_, _11970_, _11966_);
  or (_11972_, _11971_, _02131_);
  and (_11973_, _11972_, _02157_);
  and (_11974_, _11973_, _11962_);
  or (_11975_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_11976_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_11977_, _11976_, _11975_);
  and (_11978_, _11977_, _01954_);
  or (_11979_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_11980_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_11981_, _11980_, _11979_);
  and (_11982_, _11981_, _02150_);
  or (_11983_, _11982_, _11978_);
  or (_11984_, _11983_, _02144_);
  or (_11985_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_11986_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_11987_, _11986_, _11985_);
  and (_11988_, _11987_, _01954_);
  or (_11989_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_11990_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_11991_, _11990_, _11989_);
  and (_11992_, _11991_, _02150_);
  or (_11993_, _11992_, _11988_);
  or (_11994_, _11993_, _02131_);
  and (_11995_, _11994_, _02077_);
  and (_11996_, _11995_, _11984_);
  or (_11997_, _11996_, _11974_);
  and (_11998_, _11997_, _02065_);
  or (_11999_, _11998_, _11952_);
  and (_12000_, _11999_, _02143_);
  or (_12001_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_12002_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_12003_, _12002_, _12001_);
  and (_12004_, _12003_, _01954_);
  or (_12005_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_12006_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_12007_, _12006_, _12005_);
  and (_12008_, _12007_, _02150_);
  or (_12009_, _12008_, _12004_);
  and (_12010_, _12009_, _02144_);
  or (_12011_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_12012_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_12013_, _12012_, _12011_);
  and (_12014_, _12013_, _01954_);
  or (_12015_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_12016_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_12017_, _12016_, _12015_);
  and (_12018_, _12017_, _02150_);
  or (_12019_, _12018_, _12014_);
  and (_12020_, _12019_, _02131_);
  or (_12021_, _12020_, _12010_);
  and (_12022_, _12021_, _02077_);
  and (_12023_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_12024_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_12025_, _12024_, _12023_);
  and (_12026_, _12025_, _01954_);
  and (_12027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_12028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_12029_, _12028_, _12027_);
  and (_12030_, _12029_, _02150_);
  or (_12031_, _12030_, _12026_);
  and (_12032_, _12031_, _02144_);
  and (_12033_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_12034_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_12035_, _12034_, _12033_);
  and (_12036_, _12035_, _01954_);
  and (_12037_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_12038_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_12039_, _12038_, _12037_);
  and (_12040_, _12039_, _02150_);
  or (_12041_, _12040_, _12036_);
  and (_12042_, _12041_, _02131_);
  or (_12043_, _12042_, _12032_);
  and (_12044_, _12043_, _02157_);
  or (_12045_, _12044_, _12022_);
  and (_12046_, _12045_, _02065_);
  or (_12047_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_12048_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_12049_, _12048_, _02150_);
  and (_12050_, _12049_, _12047_);
  or (_12051_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_12052_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_12053_, _12052_, _01954_);
  and (_12054_, _12053_, _12051_);
  or (_12055_, _12054_, _12050_);
  and (_12056_, _12055_, _02144_);
  or (_12057_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_12058_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_12059_, _12058_, _02150_);
  and (_12060_, _12059_, _12057_);
  or (_12061_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_12062_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_12063_, _12062_, _01954_);
  and (_12064_, _12063_, _12061_);
  or (_12065_, _12064_, _12060_);
  and (_12066_, _12065_, _02131_);
  or (_12067_, _12066_, _12056_);
  and (_12068_, _12067_, _02077_);
  and (_12069_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_12070_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_12071_, _12070_, _12069_);
  and (_12072_, _12071_, _01954_);
  and (_12073_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_12074_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_12075_, _12074_, _12073_);
  and (_12076_, _12075_, _02150_);
  or (_12077_, _12076_, _12072_);
  and (_12078_, _12077_, _02144_);
  and (_12079_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_12080_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_12081_, _12080_, _12079_);
  and (_12082_, _12081_, _01954_);
  and (_12083_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_12084_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_12085_, _12084_, _12083_);
  and (_12086_, _12085_, _02150_);
  or (_12087_, _12086_, _12082_);
  and (_12088_, _12087_, _02131_);
  or (_12089_, _12088_, _12078_);
  and (_12090_, _12089_, _02157_);
  or (_12091_, _12090_, _12068_);
  and (_12092_, _12091_, _02194_);
  or (_12093_, _12092_, _12046_);
  and (_12094_, _12093_, _02005_);
  or (_12095_, _12094_, _12000_);
  or (_12096_, _12095_, _02374_);
  and (_12097_, _12096_, _11906_);
  or (_12098_, _12097_, _01748_);
  and (_12099_, _12098_, _11716_);
  or (_12100_, _12099_, _02141_);
  or (_12101_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_12102_, _12101_, _27355_);
  and (_15240_, _12102_, _12100_);
  and (_12103_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_12104_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_12105_, _12104_, _12103_);
  and (_12106_, _12105_, _01954_);
  and (_12107_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_12108_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_12109_, _12108_, _12107_);
  and (_12110_, _12109_, _02150_);
  or (_12111_, _12110_, _12106_);
  or (_12112_, _12111_, _02144_);
  and (_12113_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_12114_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_12115_, _12114_, _12113_);
  and (_12116_, _12115_, _01954_);
  and (_12117_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and (_12118_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_12119_, _12118_, _12117_);
  and (_12120_, _12119_, _02150_);
  or (_12121_, _12120_, _12116_);
  or (_12122_, _12121_, _02131_);
  and (_12123_, _12122_, _02157_);
  and (_12124_, _12123_, _12112_);
  or (_12125_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_12126_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and (_12127_, _12126_, _12125_);
  and (_12128_, _12127_, _01954_);
  or (_12129_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_12130_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_12131_, _12130_, _12129_);
  and (_12132_, _12131_, _02150_);
  or (_12133_, _12132_, _12128_);
  or (_12134_, _12133_, _02144_);
  or (_12135_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_12136_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_12137_, _12136_, _12135_);
  and (_12138_, _12137_, _01954_);
  or (_12139_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_12140_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_12141_, _12140_, _12139_);
  and (_12142_, _12141_, _02150_);
  or (_12143_, _12142_, _12138_);
  or (_12144_, _12143_, _02131_);
  and (_12145_, _12144_, _02077_);
  and (_12146_, _12145_, _12134_);
  or (_12147_, _12146_, _12124_);
  and (_12148_, _12147_, _02065_);
  and (_12149_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_12150_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_12151_, _12150_, _12149_);
  and (_12152_, _12151_, _01954_);
  and (_12153_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_12154_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_12155_, _12154_, _12153_);
  and (_12156_, _12155_, _02150_);
  or (_12157_, _12156_, _12152_);
  or (_12158_, _12157_, _02144_);
  and (_12159_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and (_12160_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_12161_, _12160_, _12159_);
  and (_12162_, _12161_, _01954_);
  and (_12163_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_12164_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_12165_, _12164_, _12163_);
  and (_12166_, _12165_, _02150_);
  or (_12167_, _12166_, _12162_);
  or (_12168_, _12167_, _02131_);
  and (_12169_, _12168_, _02157_);
  and (_12170_, _12169_, _12158_);
  or (_12171_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_12172_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_12173_, _12172_, _02150_);
  and (_12174_, _12173_, _12171_);
  or (_12175_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_12176_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_12177_, _12176_, _01954_);
  and (_12178_, _12177_, _12175_);
  or (_12179_, _12178_, _12174_);
  or (_12180_, _12179_, _02144_);
  or (_12181_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_12182_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and (_12183_, _12182_, _02150_);
  and (_12184_, _12183_, _12181_);
  or (_12185_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_12186_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_12187_, _12186_, _01954_);
  and (_12188_, _12187_, _12185_);
  or (_12189_, _12188_, _12184_);
  or (_12190_, _12189_, _02131_);
  and (_12191_, _12190_, _02077_);
  and (_12192_, _12191_, _12180_);
  or (_12193_, _12192_, _12170_);
  and (_12194_, _12193_, _02194_);
  or (_12195_, _12194_, _12148_);
  and (_12196_, _12195_, _02143_);
  and (_12197_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_12198_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_12199_, _12198_, _12197_);
  and (_12200_, _12199_, _01954_);
  and (_12201_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_12202_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_12203_, _12202_, _12201_);
  and (_12204_, _12203_, _02150_);
  or (_12205_, _12204_, _12200_);
  and (_12206_, _12205_, _02131_);
  and (_12207_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_12208_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_12209_, _12208_, _12207_);
  and (_12210_, _12209_, _01954_);
  and (_12211_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_12212_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_12213_, _12212_, _12211_);
  and (_12214_, _12213_, _02150_);
  or (_12215_, _12214_, _12210_);
  and (_12216_, _12215_, _02144_);
  or (_12217_, _12216_, _12206_);
  and (_12218_, _12217_, _02157_);
  or (_12219_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_12220_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_12221_, _12220_, _02150_);
  and (_12222_, _12221_, _12219_);
  or (_12223_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_12224_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_12225_, _12224_, _01954_);
  and (_12226_, _12225_, _12223_);
  or (_12227_, _12226_, _12222_);
  and (_12228_, _12227_, _02131_);
  or (_12229_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_12230_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_12231_, _12230_, _02150_);
  and (_12232_, _12231_, _12229_);
  or (_12233_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_12234_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_12235_, _12234_, _01954_);
  and (_12236_, _12235_, _12233_);
  or (_12237_, _12236_, _12232_);
  and (_12238_, _12237_, _02144_);
  or (_12239_, _12238_, _12228_);
  and (_12240_, _12239_, _02077_);
  or (_12241_, _12240_, _12218_);
  and (_12242_, _12241_, _02194_);
  and (_12243_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_12244_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_12245_, _12244_, _12243_);
  and (_12246_, _12245_, _01954_);
  and (_12247_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_12248_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_12249_, _12248_, _12247_);
  and (_12250_, _12249_, _02150_);
  or (_12251_, _12250_, _12246_);
  and (_12252_, _12251_, _02131_);
  and (_12253_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_12254_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_12255_, _12254_, _12253_);
  and (_12256_, _12255_, _01954_);
  and (_12257_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and (_12258_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_12259_, _12258_, _12257_);
  and (_12260_, _12259_, _02150_);
  or (_12261_, _12260_, _12256_);
  and (_12262_, _12261_, _02144_);
  or (_12263_, _12262_, _12252_);
  and (_12264_, _12263_, _02157_);
  or (_12265_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_12266_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and (_12267_, _12266_, _12265_);
  and (_12268_, _12267_, _01954_);
  or (_12269_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_12270_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_12271_, _12270_, _12269_);
  and (_12272_, _12271_, _02150_);
  or (_12273_, _12272_, _12268_);
  and (_12274_, _12273_, _02131_);
  or (_12275_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_12276_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_12277_, _12276_, _12275_);
  and (_12278_, _12277_, _01954_);
  or (_12279_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_12280_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_12281_, _12280_, _12279_);
  and (_12282_, _12281_, _02150_);
  or (_12283_, _12282_, _12278_);
  and (_12284_, _12283_, _02144_);
  or (_12285_, _12284_, _12274_);
  and (_12286_, _12285_, _02077_);
  or (_12287_, _12286_, _12264_);
  and (_12288_, _12287_, _02065_);
  or (_12289_, _12288_, _12242_);
  and (_12290_, _12289_, _02005_);
  or (_12291_, _12290_, _12196_);
  or (_12292_, _12291_, _02054_);
  and (_12293_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_12294_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_12295_, _12294_, _12293_);
  and (_12296_, _12295_, _01954_);
  and (_12297_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and (_12298_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_12299_, _12298_, _12297_);
  and (_12300_, _12299_, _02150_);
  or (_12301_, _12300_, _12296_);
  or (_12302_, _12301_, _02144_);
  and (_12303_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_12304_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_12305_, _12304_, _12303_);
  and (_12306_, _12305_, _01954_);
  and (_12307_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_12308_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_12309_, _12308_, _12307_);
  and (_12310_, _12309_, _02150_);
  or (_12311_, _12310_, _12306_);
  or (_12312_, _12311_, _02131_);
  and (_12313_, _12312_, _02157_);
  and (_12314_, _12313_, _12302_);
  or (_12315_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_12316_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and (_12317_, _12316_, _02150_);
  and (_12318_, _12317_, _12315_);
  or (_12319_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_12320_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_12321_, _12320_, _01954_);
  and (_12322_, _12321_, _12319_);
  or (_12323_, _12322_, _12318_);
  or (_12324_, _12323_, _02144_);
  or (_12325_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_12326_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and (_12327_, _12326_, _02150_);
  and (_12328_, _12327_, _12325_);
  or (_12329_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_12330_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_12331_, _12330_, _01954_);
  and (_12332_, _12331_, _12329_);
  or (_12333_, _12332_, _12328_);
  or (_12334_, _12333_, _02131_);
  and (_12335_, _12334_, _02077_);
  and (_12336_, _12335_, _12324_);
  or (_12337_, _12336_, _12314_);
  and (_12338_, _12337_, _02194_);
  and (_12339_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_12340_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_12341_, _12340_, _12339_);
  and (_12342_, _12341_, _01954_);
  and (_12343_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_12344_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_12345_, _12344_, _12343_);
  and (_12346_, _12345_, _02150_);
  or (_12347_, _12346_, _12342_);
  or (_12348_, _12347_, _02144_);
  and (_12349_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_12350_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_12351_, _12350_, _12349_);
  and (_12352_, _12351_, _01954_);
  and (_12353_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_12354_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_12355_, _12354_, _12353_);
  and (_12356_, _12355_, _02150_);
  or (_12357_, _12356_, _12352_);
  or (_12358_, _12357_, _02131_);
  and (_12359_, _12358_, _02157_);
  and (_12360_, _12359_, _12348_);
  or (_12361_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_12362_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_12363_, _12362_, _12361_);
  and (_12364_, _12363_, _01954_);
  or (_12365_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_12366_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_12367_, _12366_, _12365_);
  and (_12368_, _12367_, _02150_);
  or (_12369_, _12368_, _12364_);
  or (_12370_, _12369_, _02144_);
  or (_12371_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_12372_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_12373_, _12372_, _12371_);
  and (_12374_, _12373_, _01954_);
  or (_12375_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_12376_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_12377_, _12376_, _12375_);
  and (_12378_, _12377_, _02150_);
  or (_12379_, _12378_, _12374_);
  or (_12380_, _12379_, _02131_);
  and (_12381_, _12380_, _02077_);
  and (_12382_, _12381_, _12370_);
  or (_12383_, _12382_, _12360_);
  and (_12384_, _12383_, _02065_);
  or (_12385_, _12384_, _12338_);
  and (_12386_, _12385_, _02143_);
  or (_12387_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_12388_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_12389_, _12388_, _12387_);
  and (_12390_, _12389_, _01954_);
  or (_12391_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_12392_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and (_12393_, _12392_, _12391_);
  and (_12394_, _12393_, _02150_);
  or (_12395_, _12394_, _12390_);
  and (_12396_, _12395_, _02144_);
  or (_12397_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_12398_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_12399_, _12398_, _12397_);
  and (_12400_, _12399_, _01954_);
  or (_12401_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_12402_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_12403_, _12402_, _12401_);
  and (_12404_, _12403_, _02150_);
  or (_12405_, _12404_, _12400_);
  and (_12406_, _12405_, _02131_);
  or (_12407_, _12406_, _12396_);
  and (_12408_, _12407_, _02077_);
  and (_12409_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and (_12410_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_12411_, _12410_, _12409_);
  and (_12412_, _12411_, _01954_);
  and (_12413_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_12414_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_12415_, _12414_, _12413_);
  and (_12416_, _12415_, _02150_);
  or (_12417_, _12416_, _12412_);
  and (_12418_, _12417_, _02144_);
  and (_12419_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_12420_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_12421_, _12420_, _12419_);
  and (_12422_, _12421_, _01954_);
  and (_12423_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_12424_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_12425_, _12424_, _12423_);
  and (_12426_, _12425_, _02150_);
  or (_12427_, _12426_, _12422_);
  and (_12428_, _12427_, _02131_);
  or (_12429_, _12428_, _12418_);
  and (_12430_, _12429_, _02157_);
  or (_12431_, _12430_, _12408_);
  and (_12432_, _12431_, _02065_);
  or (_12433_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_12434_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and (_12435_, _12434_, _02150_);
  and (_12436_, _12435_, _12433_);
  or (_12437_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_12438_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and (_12439_, _12438_, _01954_);
  and (_12440_, _12439_, _12437_);
  or (_12441_, _12440_, _12436_);
  and (_12442_, _12441_, _02144_);
  or (_12443_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_12444_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_12445_, _12444_, _02150_);
  and (_12446_, _12445_, _12443_);
  or (_12447_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_12448_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and (_12449_, _12448_, _01954_);
  and (_12450_, _12449_, _12447_);
  or (_12451_, _12450_, _12446_);
  and (_12452_, _12451_, _02131_);
  or (_12453_, _12452_, _12442_);
  and (_12454_, _12453_, _02077_);
  and (_12455_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and (_12456_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_12457_, _12456_, _12455_);
  and (_12458_, _12457_, _01954_);
  and (_12459_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_12460_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_12461_, _12460_, _12459_);
  and (_12462_, _12461_, _02150_);
  or (_12463_, _12462_, _12458_);
  and (_12464_, _12463_, _02144_);
  and (_12465_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and (_12466_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_12467_, _12466_, _12465_);
  and (_12468_, _12467_, _01954_);
  and (_12469_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_12470_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_12471_, _12470_, _12469_);
  and (_12472_, _12471_, _02150_);
  or (_12473_, _12472_, _12468_);
  and (_12474_, _12473_, _02131_);
  or (_12475_, _12474_, _12464_);
  and (_12476_, _12475_, _02157_);
  or (_12477_, _12476_, _12454_);
  and (_12478_, _12477_, _02194_);
  or (_12479_, _12478_, _12432_);
  and (_12480_, _12479_, _02005_);
  or (_12481_, _12480_, _12386_);
  or (_12482_, _12481_, _02374_);
  and (_12483_, _12482_, _12292_);
  or (_12484_, _12483_, _02142_);
  and (_12485_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_12486_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_12487_, _12486_, _12485_);
  and (_12488_, _12487_, _01954_);
  and (_12489_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_12490_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_12491_, _12490_, _12489_);
  and (_12492_, _12491_, _02150_);
  or (_12493_, _12492_, _12488_);
  or (_12494_, _12493_, _02144_);
  and (_12495_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_12496_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_12497_, _12496_, _12495_);
  and (_12498_, _12497_, _01954_);
  and (_12499_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_12500_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_12501_, _12500_, _12499_);
  and (_12502_, _12501_, _02150_);
  or (_12503_, _12502_, _12498_);
  or (_12504_, _12503_, _02131_);
  and (_12505_, _12504_, _02157_);
  and (_12506_, _12505_, _12494_);
  or (_12507_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_12508_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_12509_, _12508_, _12507_);
  and (_12510_, _12509_, _01954_);
  or (_12511_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_12512_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_12513_, _12512_, _12511_);
  and (_12514_, _12513_, _02150_);
  or (_12515_, _12514_, _12510_);
  or (_12516_, _12515_, _02144_);
  or (_12517_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_12518_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_12519_, _12518_, _12517_);
  and (_12520_, _12519_, _01954_);
  or (_12521_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_12522_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_12523_, _12522_, _12521_);
  and (_12524_, _12523_, _02150_);
  or (_12525_, _12524_, _12520_);
  or (_12526_, _12525_, _02131_);
  and (_12527_, _12526_, _02077_);
  and (_12528_, _12527_, _12516_);
  or (_12529_, _12528_, _12506_);
  and (_12530_, _12529_, _02065_);
  and (_12531_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_12532_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_12533_, _12532_, _12531_);
  and (_12534_, _12533_, _01954_);
  and (_12535_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_12536_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_12537_, _12536_, _12535_);
  and (_12538_, _12537_, _02150_);
  or (_12539_, _12538_, _12534_);
  or (_12540_, _12539_, _02144_);
  and (_12541_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_12542_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_12543_, _12542_, _12541_);
  and (_12544_, _12543_, _01954_);
  and (_12545_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_12546_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_12547_, _12546_, _12545_);
  and (_12548_, _12547_, _02150_);
  or (_12549_, _12548_, _12544_);
  or (_12550_, _12549_, _02131_);
  and (_12551_, _12550_, _02157_);
  and (_12552_, _12551_, _12540_);
  or (_12553_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_12554_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_12555_, _12554_, _02150_);
  and (_12556_, _12555_, _12553_);
  or (_12557_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_12558_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_12559_, _12558_, _01954_);
  and (_12560_, _12559_, _12557_);
  or (_12561_, _12560_, _12556_);
  or (_12562_, _12561_, _02144_);
  or (_12563_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_12564_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_12565_, _12564_, _02150_);
  and (_12566_, _12565_, _12563_);
  or (_12567_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_12568_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_12569_, _12568_, _01954_);
  and (_12570_, _12569_, _12567_);
  or (_12571_, _12570_, _12566_);
  or (_12572_, _12571_, _02131_);
  and (_12573_, _12572_, _02077_);
  and (_12574_, _12573_, _12562_);
  or (_12575_, _12574_, _12552_);
  and (_12576_, _12575_, _02194_);
  or (_12577_, _12576_, _12530_);
  and (_12578_, _12577_, _02143_);
  and (_12579_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_12580_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_12581_, _12580_, _12579_);
  and (_12582_, _12581_, _01954_);
  and (_12583_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_12584_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_12585_, _12584_, _12583_);
  and (_12586_, _12585_, _02150_);
  or (_12587_, _12586_, _12582_);
  and (_12588_, _12587_, _02131_);
  and (_12589_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_12590_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_12591_, _12590_, _12589_);
  and (_12592_, _12591_, _01954_);
  and (_12593_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_12594_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_12595_, _12594_, _12593_);
  and (_12596_, _12595_, _02150_);
  or (_12597_, _12596_, _12592_);
  and (_12598_, _12597_, _02144_);
  or (_12599_, _12598_, _12588_);
  and (_12600_, _12599_, _02157_);
  or (_12601_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_12602_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_12603_, _12602_, _02150_);
  and (_12604_, _12603_, _12601_);
  or (_12605_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_12606_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_12607_, _12606_, _01954_);
  and (_12608_, _12607_, _12605_);
  or (_12609_, _12608_, _12604_);
  and (_12610_, _12609_, _02131_);
  or (_12611_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_12612_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_12613_, _12612_, _02150_);
  and (_12614_, _12613_, _12611_);
  or (_12615_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_12616_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_12617_, _12616_, _01954_);
  and (_12618_, _12617_, _12615_);
  or (_12619_, _12618_, _12614_);
  and (_12620_, _12619_, _02144_);
  or (_12621_, _12620_, _12610_);
  and (_12622_, _12621_, _02077_);
  or (_12623_, _12622_, _12600_);
  and (_12624_, _12623_, _02194_);
  and (_12625_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_12626_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_12627_, _12626_, _12625_);
  and (_12628_, _12627_, _01954_);
  and (_12629_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_12630_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_12631_, _12630_, _12629_);
  and (_12632_, _12631_, _02150_);
  or (_12633_, _12632_, _12628_);
  and (_12634_, _12633_, _02131_);
  and (_12635_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_12636_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_12637_, _12636_, _12635_);
  and (_12638_, _12637_, _01954_);
  and (_12639_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_12640_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_12641_, _12640_, _12639_);
  and (_12642_, _12641_, _02150_);
  or (_12643_, _12642_, _12638_);
  and (_12644_, _12643_, _02144_);
  or (_12645_, _12644_, _12634_);
  and (_12646_, _12645_, _02157_);
  or (_12647_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_12648_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_12649_, _12648_, _12647_);
  and (_12650_, _12649_, _01954_);
  or (_12651_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_12652_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_12653_, _12652_, _12651_);
  and (_12654_, _12653_, _02150_);
  or (_12655_, _12654_, _12650_);
  and (_12656_, _12655_, _02131_);
  or (_12657_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_12658_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_12659_, _12658_, _12657_);
  and (_12660_, _12659_, _01954_);
  or (_12661_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_12662_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_12663_, _12662_, _12661_);
  and (_12664_, _12663_, _02150_);
  or (_12665_, _12664_, _12660_);
  and (_12666_, _12665_, _02144_);
  or (_12667_, _12666_, _12656_);
  and (_12668_, _12667_, _02077_);
  or (_12669_, _12668_, _12646_);
  and (_12670_, _12669_, _02065_);
  or (_12671_, _12670_, _12624_);
  and (_12672_, _12671_, _02005_);
  or (_12673_, _12672_, _12578_);
  or (_12674_, _12673_, _02054_);
  and (_12675_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_12676_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_12677_, _12676_, _12675_);
  and (_12678_, _12677_, _01954_);
  and (_12679_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_12680_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_12681_, _12680_, _12679_);
  and (_12682_, _12681_, _02150_);
  or (_12683_, _12682_, _12678_);
  or (_12684_, _12683_, _02144_);
  and (_12685_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_12686_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_12687_, _12686_, _12685_);
  and (_12688_, _12687_, _01954_);
  and (_12689_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_12690_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_12691_, _12690_, _12689_);
  and (_12692_, _12691_, _02150_);
  or (_12693_, _12692_, _12688_);
  or (_12694_, _12693_, _02131_);
  and (_12695_, _12694_, _02157_);
  and (_12696_, _12695_, _12684_);
  or (_12697_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_12698_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_12699_, _12698_, _02150_);
  and (_12700_, _12699_, _12697_);
  or (_12701_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_12702_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_12703_, _12702_, _01954_);
  and (_12704_, _12703_, _12701_);
  or (_12705_, _12704_, _12700_);
  or (_12706_, _12705_, _02144_);
  or (_12707_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_12708_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_12709_, _12708_, _02150_);
  and (_12710_, _12709_, _12707_);
  or (_12711_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_12712_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_12713_, _12712_, _01954_);
  and (_12714_, _12713_, _12711_);
  or (_12715_, _12714_, _12710_);
  or (_12716_, _12715_, _02131_);
  and (_12717_, _12716_, _02077_);
  and (_12718_, _12717_, _12706_);
  or (_12719_, _12718_, _12696_);
  and (_12720_, _12719_, _02194_);
  and (_12721_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_12722_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_12723_, _12722_, _12721_);
  and (_12724_, _12723_, _01954_);
  and (_12725_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_12726_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_12727_, _12726_, _12725_);
  and (_12728_, _12727_, _02150_);
  or (_12729_, _12728_, _12724_);
  or (_12730_, _12729_, _02144_);
  and (_12731_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_12732_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_12733_, _12732_, _12731_);
  and (_12734_, _12733_, _01954_);
  and (_12735_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_12736_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_12737_, _12736_, _12735_);
  and (_12738_, _12737_, _02150_);
  or (_12739_, _12738_, _12734_);
  or (_12740_, _12739_, _02131_);
  and (_12741_, _12740_, _02157_);
  and (_12742_, _12741_, _12730_);
  or (_12744_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_12745_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_12746_, _12745_, _12744_);
  and (_12747_, _12746_, _01954_);
  or (_12748_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_12749_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_12750_, _12749_, _12748_);
  and (_12751_, _12750_, _02150_);
  or (_12752_, _12751_, _12747_);
  or (_12753_, _12752_, _02144_);
  or (_12754_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_12755_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_12756_, _12755_, _12754_);
  and (_12757_, _12756_, _01954_);
  or (_12758_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_12759_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_12760_, _12759_, _12758_);
  and (_12761_, _12760_, _02150_);
  or (_12762_, _12761_, _12757_);
  or (_12763_, _12762_, _02131_);
  and (_12765_, _12763_, _02077_);
  and (_12766_, _12765_, _12753_);
  or (_12767_, _12766_, _12742_);
  and (_12768_, _12767_, _02065_);
  or (_12769_, _12768_, _12720_);
  and (_12770_, _12769_, _02143_);
  or (_12771_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_12772_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_12773_, _12772_, _12771_);
  and (_12774_, _12773_, _01954_);
  or (_12775_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_12776_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_12777_, _12776_, _12775_);
  and (_12778_, _12777_, _02150_);
  or (_12779_, _12778_, _12774_);
  and (_12780_, _12779_, _02144_);
  or (_12781_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_12782_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_12783_, _12782_, _12781_);
  and (_12784_, _12783_, _01954_);
  or (_12785_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_12786_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_12787_, _12786_, _12785_);
  and (_12788_, _12787_, _02150_);
  or (_12789_, _12788_, _12784_);
  and (_12790_, _12789_, _02131_);
  or (_12791_, _12790_, _12780_);
  and (_12792_, _12791_, _02077_);
  and (_12793_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_12794_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_12795_, _12794_, _12793_);
  and (_12796_, _12795_, _01954_);
  and (_12797_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_12798_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_12799_, _12798_, _12797_);
  and (_12800_, _12799_, _02150_);
  or (_12801_, _12800_, _12796_);
  and (_12802_, _12801_, _02144_);
  and (_12803_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_12804_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_12805_, _12804_, _12803_);
  and (_12806_, _12805_, _01954_);
  and (_12807_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_12808_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_12809_, _12808_, _12807_);
  and (_12810_, _12809_, _02150_);
  or (_12811_, _12810_, _12806_);
  and (_12812_, _12811_, _02131_);
  or (_12813_, _12812_, _12802_);
  and (_12814_, _12813_, _02157_);
  or (_12815_, _12814_, _12792_);
  and (_12816_, _12815_, _02065_);
  or (_12817_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_12818_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_12819_, _12818_, _02150_);
  and (_12820_, _12819_, _12817_);
  or (_12821_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_12822_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_12823_, _12822_, _01954_);
  and (_12824_, _12823_, _12821_);
  or (_12825_, _12824_, _12820_);
  and (_12826_, _12825_, _02144_);
  or (_12827_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_12828_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_12829_, _12828_, _02150_);
  and (_12830_, _12829_, _12827_);
  or (_12831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_12832_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_12833_, _12832_, _01954_);
  and (_12834_, _12833_, _12831_);
  or (_12835_, _12834_, _12830_);
  and (_12836_, _12835_, _02131_);
  or (_12837_, _12836_, _12826_);
  and (_12838_, _12837_, _02077_);
  and (_12839_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_12840_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_12841_, _12840_, _12839_);
  and (_12842_, _12841_, _01954_);
  and (_12843_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_12844_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_12845_, _12844_, _12843_);
  and (_12846_, _12845_, _02150_);
  or (_12847_, _12846_, _12842_);
  and (_12848_, _12847_, _02144_);
  and (_12849_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_12850_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_12851_, _12850_, _12849_);
  and (_12852_, _12851_, _01954_);
  and (_12853_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_12854_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_12855_, _12854_, _12853_);
  and (_12856_, _12855_, _02150_);
  or (_12857_, _12856_, _12852_);
  and (_12858_, _12857_, _02131_);
  or (_12859_, _12858_, _12848_);
  and (_12860_, _12859_, _02157_);
  or (_12861_, _12860_, _12838_);
  and (_12862_, _12861_, _02194_);
  or (_12863_, _12862_, _12816_);
  and (_12864_, _12863_, _02005_);
  or (_12865_, _12864_, _12770_);
  or (_12866_, _12865_, _02374_);
  and (_12867_, _12866_, _12674_);
  or (_12868_, _12867_, _01748_);
  and (_12869_, _12868_, _12484_);
  or (_12870_, _12869_, _02141_);
  or (_12871_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_12872_, _12871_, _27355_);
  and (_15242_, _12872_, _12870_);
  and (_12873_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_12874_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_12875_, _12874_, _12873_);
  and (_12876_, _12875_, _01954_);
  and (_12877_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_12878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_12879_, _12878_, _12877_);
  and (_12880_, _12879_, _02150_);
  or (_12881_, _12880_, _12876_);
  or (_12882_, _12881_, _02144_);
  and (_12883_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_12884_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_12885_, _12884_, _12883_);
  and (_12886_, _12885_, _01954_);
  and (_12887_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and (_12888_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_12889_, _12888_, _12887_);
  and (_12890_, _12889_, _02150_);
  or (_12891_, _12890_, _12886_);
  or (_12892_, _12891_, _02131_);
  and (_12893_, _12892_, _02157_);
  and (_12894_, _12893_, _12882_);
  or (_12895_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_12896_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_12897_, _12896_, _12895_);
  and (_12898_, _12897_, _01954_);
  or (_12899_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_12900_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and (_12901_, _12900_, _12899_);
  and (_12902_, _12901_, _02150_);
  or (_12903_, _12902_, _12898_);
  or (_12904_, _12903_, _02144_);
  or (_12905_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_12906_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_12907_, _12906_, _12905_);
  and (_12908_, _12907_, _01954_);
  or (_12909_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_12910_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_12911_, _12910_, _12909_);
  and (_12912_, _12911_, _02150_);
  or (_12913_, _12912_, _12908_);
  or (_12914_, _12913_, _02131_);
  and (_12915_, _12914_, _02077_);
  and (_12916_, _12915_, _12904_);
  or (_12917_, _12916_, _12894_);
  and (_12918_, _12917_, _02065_);
  and (_12919_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_12920_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_12921_, _12920_, _12919_);
  and (_12922_, _12921_, _01954_);
  and (_12923_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and (_12924_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_12925_, _12924_, _12923_);
  and (_12926_, _12925_, _02150_);
  or (_12927_, _12926_, _12922_);
  or (_12928_, _12927_, _02144_);
  and (_12929_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_12930_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_12931_, _12930_, _12929_);
  and (_12932_, _12931_, _01954_);
  and (_12933_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_12934_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_12935_, _12934_, _12933_);
  and (_12936_, _12935_, _02150_);
  or (_12937_, _12936_, _12932_);
  or (_12938_, _12937_, _02131_);
  and (_12939_, _12938_, _02157_);
  and (_12940_, _12939_, _12928_);
  or (_12941_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_12942_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_12943_, _12942_, _02150_);
  and (_12944_, _12943_, _12941_);
  or (_12945_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_12946_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_12947_, _12946_, _01954_);
  and (_12948_, _12947_, _12945_);
  or (_12949_, _12948_, _12944_);
  or (_12950_, _12949_, _02144_);
  or (_12951_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_12952_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_12953_, _12952_, _02150_);
  and (_12954_, _12953_, _12951_);
  or (_12955_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_12956_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and (_12957_, _12956_, _01954_);
  and (_12958_, _12957_, _12955_);
  or (_12959_, _12958_, _12954_);
  or (_12960_, _12959_, _02131_);
  and (_12961_, _12960_, _02077_);
  and (_12962_, _12961_, _12950_);
  or (_12963_, _12962_, _12940_);
  and (_12964_, _12963_, _02194_);
  or (_12965_, _12964_, _12918_);
  and (_12966_, _12965_, _02143_);
  and (_12967_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_12968_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_12969_, _12968_, _12967_);
  and (_12970_, _12969_, _01954_);
  and (_12971_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_12972_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_12973_, _12972_, _12971_);
  and (_12974_, _12973_, _02150_);
  or (_12975_, _12974_, _12970_);
  and (_12976_, _12975_, _02131_);
  and (_12977_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_12978_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_12979_, _12978_, _12977_);
  and (_12980_, _12979_, _01954_);
  and (_12981_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_12982_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_12983_, _12982_, _12981_);
  and (_12984_, _12983_, _02150_);
  or (_12985_, _12984_, _12980_);
  and (_12986_, _12985_, _02144_);
  or (_12987_, _12986_, _12976_);
  and (_12988_, _12987_, _02157_);
  or (_12989_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_12990_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_12991_, _12990_, _02150_);
  and (_12992_, _12991_, _12989_);
  or (_12993_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_12994_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_12995_, _12994_, _01954_);
  and (_12996_, _12995_, _12993_);
  or (_12997_, _12996_, _12992_);
  and (_12998_, _12997_, _02131_);
  or (_12999_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_13000_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_13001_, _13000_, _02150_);
  and (_13002_, _13001_, _12999_);
  or (_13003_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_13004_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_13005_, _13004_, _01954_);
  and (_13006_, _13005_, _13003_);
  or (_13007_, _13006_, _13002_);
  and (_13008_, _13007_, _02144_);
  or (_13009_, _13008_, _12998_);
  and (_13010_, _13009_, _02077_);
  or (_13011_, _13010_, _12988_);
  and (_13012_, _13011_, _02194_);
  and (_13013_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_13014_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_13015_, _13014_, _13013_);
  and (_13016_, _13015_, _01954_);
  and (_13017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_13018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_13019_, _13018_, _13017_);
  and (_13020_, _13019_, _02150_);
  or (_13021_, _13020_, _13016_);
  and (_13022_, _13021_, _02131_);
  and (_13023_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_13024_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_13025_, _13024_, _13023_);
  and (_13026_, _13025_, _01954_);
  and (_13027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_13028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_13029_, _13028_, _13027_);
  and (_13030_, _13029_, _02150_);
  or (_13031_, _13030_, _13026_);
  and (_13032_, _13031_, _02144_);
  or (_13033_, _13032_, _13022_);
  and (_13034_, _13033_, _02157_);
  or (_13035_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_13036_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_13037_, _13036_, _13035_);
  and (_13038_, _13037_, _01954_);
  or (_13039_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_13040_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_13041_, _13040_, _13039_);
  and (_13042_, _13041_, _02150_);
  or (_13043_, _13042_, _13038_);
  and (_13044_, _13043_, _02131_);
  or (_13045_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_13046_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_13047_, _13046_, _13045_);
  and (_13048_, _13047_, _01954_);
  or (_13049_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_13050_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_13051_, _13050_, _13049_);
  and (_13052_, _13051_, _02150_);
  or (_13053_, _13052_, _13048_);
  and (_13054_, _13053_, _02144_);
  or (_13055_, _13054_, _13044_);
  and (_13056_, _13055_, _02077_);
  or (_13057_, _13056_, _13034_);
  and (_13058_, _13057_, _02065_);
  or (_13059_, _13058_, _13012_);
  and (_13060_, _13059_, _02005_);
  or (_13061_, _13060_, _12966_);
  or (_13062_, _13061_, _02054_);
  and (_13063_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and (_13064_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_13065_, _13064_, _13063_);
  and (_13066_, _13065_, _01954_);
  and (_13067_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_13068_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_13069_, _13068_, _13067_);
  and (_13070_, _13069_, _02150_);
  or (_13071_, _13070_, _13066_);
  or (_13072_, _13071_, _02144_);
  and (_13073_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_13074_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_13075_, _13074_, _13073_);
  and (_13076_, _13075_, _01954_);
  and (_13077_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_13078_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_13079_, _13078_, _13077_);
  and (_13080_, _13079_, _02150_);
  or (_13081_, _13080_, _13076_);
  or (_13082_, _13081_, _02131_);
  and (_13083_, _13082_, _02157_);
  and (_13084_, _13083_, _13072_);
  or (_13085_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_13086_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_13087_, _13086_, _02150_);
  and (_13088_, _13087_, _13085_);
  or (_13089_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_13090_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_13091_, _13090_, _01954_);
  and (_13092_, _13091_, _13089_);
  or (_13093_, _13092_, _13088_);
  or (_13094_, _13093_, _02144_);
  or (_13095_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_13096_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_13097_, _13096_, _02150_);
  and (_13098_, _13097_, _13095_);
  or (_13099_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_13100_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and (_13101_, _13100_, _01954_);
  and (_13102_, _13101_, _13099_);
  or (_13103_, _13102_, _13098_);
  or (_13104_, _13103_, _02131_);
  and (_13105_, _13104_, _02077_);
  and (_13106_, _13105_, _13094_);
  or (_13107_, _13106_, _13084_);
  and (_13108_, _13107_, _02194_);
  and (_13109_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_13110_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_13111_, _13110_, _13109_);
  and (_13112_, _13111_, _01954_);
  and (_13113_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_13114_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_13115_, _13114_, _13113_);
  and (_13116_, _13115_, _02150_);
  or (_13117_, _13116_, _13112_);
  or (_13118_, _13117_, _02144_);
  and (_13119_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_13120_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_13121_, _13120_, _13119_);
  and (_13122_, _13121_, _01954_);
  and (_13123_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_13124_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_13125_, _13124_, _13123_);
  and (_13126_, _13125_, _02150_);
  or (_13127_, _13126_, _13122_);
  or (_13128_, _13127_, _02131_);
  and (_13129_, _13128_, _02157_);
  and (_13130_, _13129_, _13118_);
  or (_13131_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_13132_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_13133_, _13132_, _13131_);
  and (_13134_, _13133_, _01954_);
  or (_13135_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_13136_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_13137_, _13136_, _13135_);
  and (_13138_, _13137_, _02150_);
  or (_13139_, _13138_, _13134_);
  or (_13140_, _13139_, _02144_);
  or (_13141_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_13142_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_13143_, _13142_, _13141_);
  and (_13144_, _13143_, _01954_);
  or (_13145_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_13146_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_13147_, _13146_, _13145_);
  and (_13148_, _13147_, _02150_);
  or (_13149_, _13148_, _13144_);
  or (_13150_, _13149_, _02131_);
  and (_13151_, _13150_, _02077_);
  and (_13152_, _13151_, _13140_);
  or (_13153_, _13152_, _13130_);
  and (_13154_, _13153_, _02065_);
  or (_13155_, _13154_, _13108_);
  and (_13156_, _13155_, _02143_);
  or (_13157_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_13158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and (_13159_, _13158_, _13157_);
  and (_13160_, _13159_, _01954_);
  or (_13161_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_13162_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_13163_, _13162_, _13161_);
  and (_13164_, _13163_, _02150_);
  or (_13165_, _13164_, _13160_);
  and (_13166_, _13165_, _02144_);
  or (_13167_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_13168_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_13169_, _13168_, _13167_);
  and (_13170_, _13169_, _01954_);
  or (_13171_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_13172_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and (_13173_, _13172_, _13171_);
  and (_13174_, _13173_, _02150_);
  or (_13175_, _13174_, _13170_);
  and (_13176_, _13175_, _02131_);
  or (_13177_, _13176_, _13166_);
  and (_13178_, _13177_, _02077_);
  and (_13179_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_13180_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_13181_, _13180_, _13179_);
  and (_13182_, _13181_, _01954_);
  and (_13183_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_13184_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_13185_, _13184_, _13183_);
  and (_13186_, _13185_, _02150_);
  or (_13187_, _13186_, _13182_);
  and (_13188_, _13187_, _02144_);
  and (_13189_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_13190_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_13191_, _13190_, _13189_);
  and (_13192_, _13191_, _01954_);
  and (_13193_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_13194_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_13195_, _13194_, _13193_);
  and (_13196_, _13195_, _02150_);
  or (_13197_, _13196_, _13192_);
  and (_13198_, _13197_, _02131_);
  or (_13199_, _13198_, _13188_);
  and (_13200_, _13199_, _02157_);
  or (_13201_, _13200_, _13178_);
  and (_13202_, _13201_, _02065_);
  or (_13203_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_13204_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and (_13205_, _13204_, _02150_);
  and (_13206_, _13205_, _13203_);
  or (_13207_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_13208_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and (_13209_, _13208_, _01954_);
  and (_13210_, _13209_, _13207_);
  or (_13211_, _13210_, _13206_);
  and (_13212_, _13211_, _02144_);
  or (_13213_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_13214_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and (_13215_, _13214_, _02150_);
  and (_13216_, _13215_, _13213_);
  or (_13217_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_13218_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and (_13219_, _13218_, _01954_);
  and (_13220_, _13219_, _13217_);
  or (_13221_, _13220_, _13216_);
  and (_13222_, _13221_, _02131_);
  or (_13223_, _13222_, _13212_);
  and (_13224_, _13223_, _02077_);
  and (_13225_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and (_13226_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_13227_, _13226_, _13225_);
  and (_13228_, _13227_, _01954_);
  and (_13229_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and (_13230_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_13231_, _13230_, _13229_);
  and (_13232_, _13231_, _02150_);
  or (_13233_, _13232_, _13228_);
  and (_13234_, _13233_, _02144_);
  and (_13235_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and (_13236_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_13237_, _13236_, _13235_);
  and (_13238_, _13237_, _01954_);
  and (_13239_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and (_13240_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_13241_, _13240_, _13239_);
  and (_13242_, _13241_, _02150_);
  or (_13243_, _13242_, _13238_);
  and (_13244_, _13243_, _02131_);
  or (_13245_, _13244_, _13234_);
  and (_13246_, _13245_, _02157_);
  or (_13247_, _13246_, _13224_);
  and (_13248_, _13247_, _02194_);
  or (_13249_, _13248_, _13202_);
  and (_13250_, _13249_, _02005_);
  or (_13251_, _13250_, _13156_);
  or (_13252_, _13251_, _02374_);
  and (_13253_, _13252_, _13062_);
  or (_13254_, _13253_, _02142_);
  and (_13255_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_13256_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_13257_, _13256_, _13255_);
  and (_13258_, _13257_, _01954_);
  and (_13259_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_13260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_13261_, _13260_, _13259_);
  and (_13262_, _13261_, _02150_);
  or (_13263_, _13262_, _13258_);
  or (_13264_, _13263_, _02144_);
  and (_13265_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_13266_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_13267_, _13266_, _13265_);
  and (_13268_, _13267_, _01954_);
  and (_13269_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_13270_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_13271_, _13270_, _13269_);
  and (_13272_, _13271_, _02150_);
  or (_13273_, _13272_, _13268_);
  or (_13274_, _13273_, _02131_);
  and (_13275_, _13274_, _02157_);
  and (_13276_, _13275_, _13264_);
  or (_13277_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_13278_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_13279_, _13278_, _13277_);
  and (_13280_, _13279_, _01954_);
  or (_13281_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_13282_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_13283_, _13282_, _13281_);
  and (_13284_, _13283_, _02150_);
  or (_13285_, _13284_, _13280_);
  or (_13286_, _13285_, _02144_);
  or (_13287_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_13288_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_13289_, _13288_, _13287_);
  and (_13290_, _13289_, _01954_);
  or (_13291_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_13292_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_13293_, _13292_, _13291_);
  and (_13294_, _13293_, _02150_);
  or (_13295_, _13294_, _13290_);
  or (_13296_, _13295_, _02131_);
  and (_13297_, _13296_, _02077_);
  and (_13298_, _13297_, _13286_);
  or (_13299_, _13298_, _13276_);
  and (_13300_, _13299_, _02065_);
  and (_13301_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_13302_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_13303_, _13302_, _13301_);
  and (_13304_, _13303_, _01954_);
  and (_13305_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_13306_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_13307_, _13306_, _13305_);
  and (_13308_, _13307_, _02150_);
  or (_13309_, _13308_, _13304_);
  or (_13310_, _13309_, _02144_);
  and (_13311_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_13312_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_13313_, _13312_, _13311_);
  and (_13314_, _13313_, _01954_);
  and (_13315_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_13316_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_13317_, _13316_, _13315_);
  and (_13318_, _13317_, _02150_);
  or (_13319_, _13318_, _13314_);
  or (_13320_, _13319_, _02131_);
  and (_13321_, _13320_, _02157_);
  and (_13322_, _13321_, _13310_);
  or (_13323_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_13324_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_13325_, _13324_, _02150_);
  and (_13326_, _13325_, _13323_);
  or (_13327_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_13328_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_13329_, _13328_, _01954_);
  and (_13330_, _13329_, _13327_);
  or (_13331_, _13330_, _13326_);
  or (_13332_, _13331_, _02144_);
  or (_13333_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_13334_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_13335_, _13334_, _02150_);
  and (_13336_, _13335_, _13333_);
  or (_13337_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_13338_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_13339_, _13338_, _01954_);
  and (_13340_, _13339_, _13337_);
  or (_13341_, _13340_, _13336_);
  or (_13342_, _13341_, _02131_);
  and (_13343_, _13342_, _02077_);
  and (_13344_, _13343_, _13332_);
  or (_13345_, _13344_, _13322_);
  and (_13346_, _13345_, _02194_);
  or (_13347_, _13346_, _13300_);
  and (_13348_, _13347_, _02143_);
  and (_13349_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_13350_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_13351_, _13350_, _13349_);
  and (_13352_, _13351_, _01954_);
  and (_13353_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_13354_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_13355_, _13354_, _13353_);
  and (_13356_, _13355_, _02150_);
  or (_13357_, _13356_, _13352_);
  and (_13358_, _13357_, _02131_);
  and (_13359_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_13360_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_13361_, _13360_, _13359_);
  and (_13362_, _13361_, _01954_);
  and (_13363_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_13364_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_13365_, _13364_, _13363_);
  and (_13366_, _13365_, _02150_);
  or (_13367_, _13366_, _13362_);
  and (_13368_, _13367_, _02144_);
  or (_13369_, _13368_, _13358_);
  and (_13370_, _13369_, _02157_);
  or (_13371_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_13372_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_13373_, _13372_, _02150_);
  and (_13374_, _13373_, _13371_);
  or (_13375_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_13376_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_13377_, _13376_, _01954_);
  and (_13378_, _13377_, _13375_);
  or (_13379_, _13378_, _13374_);
  and (_13380_, _13379_, _02131_);
  or (_13381_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_13382_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_13383_, _13382_, _02150_);
  and (_13384_, _13383_, _13381_);
  or (_13385_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_13386_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_13387_, _13386_, _01954_);
  and (_13388_, _13387_, _13385_);
  or (_13389_, _13388_, _13384_);
  and (_13390_, _13389_, _02144_);
  or (_13391_, _13390_, _13380_);
  and (_13392_, _13391_, _02077_);
  or (_13393_, _13392_, _13370_);
  and (_13394_, _13393_, _02194_);
  and (_13395_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_13396_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_13397_, _13396_, _13395_);
  and (_13398_, _13397_, _01954_);
  and (_13399_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_13400_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_13401_, _13400_, _13399_);
  and (_13402_, _13401_, _02150_);
  or (_13403_, _13402_, _13398_);
  and (_13404_, _13403_, _02131_);
  and (_13405_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_13406_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_13407_, _13406_, _13405_);
  and (_13408_, _13407_, _01954_);
  and (_13409_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_13410_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_13411_, _13410_, _13409_);
  and (_13412_, _13411_, _02150_);
  or (_13413_, _13412_, _13408_);
  and (_13414_, _13413_, _02144_);
  or (_13415_, _13414_, _13404_);
  and (_13416_, _13415_, _02157_);
  or (_13417_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_13418_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_13419_, _13418_, _13417_);
  and (_13420_, _13419_, _01954_);
  or (_13421_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_13422_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_13423_, _13422_, _13421_);
  and (_13424_, _13423_, _02150_);
  or (_13425_, _13424_, _13420_);
  and (_13426_, _13425_, _02131_);
  or (_13427_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_13428_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_13429_, _13428_, _13427_);
  and (_13430_, _13429_, _01954_);
  or (_13431_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_13432_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_13433_, _13432_, _13431_);
  and (_13434_, _13433_, _02150_);
  or (_13435_, _13434_, _13430_);
  and (_13436_, _13435_, _02144_);
  or (_13437_, _13436_, _13426_);
  and (_13438_, _13437_, _02077_);
  or (_13439_, _13438_, _13416_);
  and (_13440_, _13439_, _02065_);
  or (_13441_, _13440_, _13394_);
  and (_13442_, _13441_, _02005_);
  or (_13443_, _13442_, _13348_);
  or (_13444_, _13443_, _02054_);
  and (_13445_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_13446_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_13447_, _13446_, _13445_);
  and (_13448_, _13447_, _01954_);
  and (_13449_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_13450_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_13451_, _13450_, _13449_);
  and (_13452_, _13451_, _02150_);
  or (_13453_, _13452_, _13448_);
  or (_13454_, _13453_, _02144_);
  and (_13455_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_13456_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_13457_, _13456_, _13455_);
  and (_13458_, _13457_, _01954_);
  and (_13459_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_13460_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_13461_, _13460_, _13459_);
  and (_13462_, _13461_, _02150_);
  or (_13463_, _13462_, _13458_);
  or (_13464_, _13463_, _02131_);
  and (_13465_, _13464_, _02157_);
  and (_13466_, _13465_, _13454_);
  or (_13467_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_13468_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_13469_, _13468_, _02150_);
  and (_13470_, _13469_, _13467_);
  or (_13471_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_13472_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_13473_, _13472_, _01954_);
  and (_13474_, _13473_, _13471_);
  or (_13475_, _13474_, _13470_);
  or (_13476_, _13475_, _02144_);
  or (_13477_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_13478_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_13479_, _13478_, _02150_);
  and (_13480_, _13479_, _13477_);
  or (_13481_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_13482_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_13483_, _13482_, _01954_);
  and (_13484_, _13483_, _13481_);
  or (_13485_, _13484_, _13480_);
  or (_13486_, _13485_, _02131_);
  and (_13487_, _13486_, _02077_);
  and (_13488_, _13487_, _13476_);
  or (_13489_, _13488_, _13466_);
  and (_13490_, _13489_, _02194_);
  and (_13491_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_13492_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_13493_, _13492_, _13491_);
  and (_13494_, _13493_, _01954_);
  and (_13495_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_13496_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_13497_, _13496_, _13495_);
  and (_13498_, _13497_, _02150_);
  or (_13499_, _13498_, _13494_);
  or (_13500_, _13499_, _02144_);
  and (_13501_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_13502_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_13503_, _13502_, _13501_);
  and (_13504_, _13503_, _01954_);
  and (_13505_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_13506_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_13507_, _13506_, _13505_);
  and (_13508_, _13507_, _02150_);
  or (_13509_, _13508_, _13504_);
  or (_13510_, _13509_, _02131_);
  and (_13511_, _13510_, _02157_);
  and (_13512_, _13511_, _13500_);
  or (_13513_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_13514_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_13515_, _13514_, _13513_);
  and (_13516_, _13515_, _01954_);
  or (_13517_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_13518_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_13519_, _13518_, _13517_);
  and (_13520_, _13519_, _02150_);
  or (_13521_, _13520_, _13516_);
  or (_13522_, _13521_, _02144_);
  or (_13523_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_13524_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_13525_, _13524_, _13523_);
  and (_13526_, _13525_, _01954_);
  or (_13527_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_13528_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_13529_, _13528_, _13527_);
  and (_13530_, _13529_, _02150_);
  or (_13531_, _13530_, _13526_);
  or (_13532_, _13531_, _02131_);
  and (_13533_, _13532_, _02077_);
  and (_13534_, _13533_, _13522_);
  or (_13535_, _13534_, _13512_);
  and (_13536_, _13535_, _02065_);
  or (_13537_, _13536_, _13490_);
  and (_13538_, _13537_, _02143_);
  or (_13539_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_13540_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_13541_, _13540_, _13539_);
  and (_13542_, _13541_, _01954_);
  or (_13543_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_13544_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_13545_, _13544_, _13543_);
  and (_13546_, _13545_, _02150_);
  or (_13547_, _13546_, _13542_);
  and (_13548_, _13547_, _02144_);
  or (_13549_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_13550_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_13551_, _13550_, _13549_);
  and (_13552_, _13551_, _01954_);
  or (_13553_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_13554_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_13555_, _13554_, _13553_);
  and (_13556_, _13555_, _02150_);
  or (_13557_, _13556_, _13552_);
  and (_13558_, _13557_, _02131_);
  or (_13559_, _13558_, _13548_);
  and (_13560_, _13559_, _02077_);
  and (_13561_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_13562_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_13563_, _13562_, _13561_);
  and (_13564_, _13563_, _01954_);
  and (_13565_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_13566_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_13567_, _13566_, _13565_);
  and (_13568_, _13567_, _02150_);
  or (_13569_, _13568_, _13564_);
  and (_13570_, _13569_, _02144_);
  and (_13571_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_13572_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_13573_, _13572_, _13571_);
  and (_13574_, _13573_, _01954_);
  and (_13575_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_13576_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_13577_, _13576_, _13575_);
  and (_13578_, _13577_, _02150_);
  or (_13579_, _13578_, _13574_);
  and (_13580_, _13579_, _02131_);
  or (_13581_, _13580_, _13570_);
  and (_13582_, _13581_, _02157_);
  or (_13583_, _13582_, _13560_);
  and (_13584_, _13583_, _02065_);
  or (_13585_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_13586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_13587_, _13586_, _02150_);
  and (_13588_, _13587_, _13585_);
  or (_13589_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_13590_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_13591_, _13590_, _01954_);
  and (_13592_, _13591_, _13589_);
  or (_13593_, _13592_, _13588_);
  and (_13594_, _13593_, _02144_);
  or (_13595_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_13596_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_13597_, _13596_, _02150_);
  and (_13598_, _13597_, _13595_);
  or (_13599_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_13600_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_13601_, _13600_, _01954_);
  and (_13602_, _13601_, _13599_);
  or (_13603_, _13602_, _13598_);
  and (_13604_, _13603_, _02131_);
  or (_13605_, _13604_, _13594_);
  and (_13606_, _13605_, _02077_);
  and (_13607_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_13608_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_13609_, _13608_, _13607_);
  and (_13610_, _13609_, _01954_);
  and (_13611_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_13612_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_13613_, _13612_, _13611_);
  and (_13614_, _13613_, _02150_);
  or (_13615_, _13614_, _13610_);
  and (_13616_, _13615_, _02144_);
  and (_13617_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_13618_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_13619_, _13618_, _13617_);
  and (_13620_, _13619_, _01954_);
  and (_13621_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_13622_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_13623_, _13622_, _13621_);
  and (_13624_, _13623_, _02150_);
  or (_13625_, _13624_, _13620_);
  and (_13626_, _13625_, _02131_);
  or (_13627_, _13626_, _13616_);
  and (_13628_, _13627_, _02157_);
  or (_13629_, _13628_, _13606_);
  and (_13630_, _13629_, _02194_);
  or (_13631_, _13630_, _13584_);
  and (_13632_, _13631_, _02005_);
  or (_13633_, _13632_, _13538_);
  or (_13634_, _13633_, _02374_);
  and (_13635_, _13634_, _13444_);
  or (_13636_, _13635_, _01748_);
  and (_13637_, _13636_, _13254_);
  or (_13638_, _13637_, _02141_);
  or (_13639_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_13640_, _13639_, _27355_);
  and (_15244_, _13640_, _13638_);
  and (_13641_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_13642_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_13643_, _13642_, _13641_);
  and (_13644_, _13643_, _01954_);
  and (_13645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_13646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_13647_, _13646_, _13645_);
  and (_13648_, _13647_, _02150_);
  or (_13649_, _13648_, _13644_);
  or (_13650_, _13649_, _02144_);
  and (_13651_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_13652_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_13653_, _13652_, _13651_);
  and (_13654_, _13653_, _01954_);
  and (_13655_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and (_13656_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_13657_, _13656_, _13655_);
  and (_13658_, _13657_, _02150_);
  or (_13659_, _13658_, _13654_);
  or (_13660_, _13659_, _02131_);
  and (_13661_, _13660_, _02157_);
  and (_13662_, _13661_, _13650_);
  or (_13663_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_13664_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_13665_, _13664_, _13663_);
  and (_13666_, _13665_, _01954_);
  or (_13667_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_13668_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_13669_, _13668_, _13667_);
  and (_13670_, _13669_, _02150_);
  or (_13671_, _13670_, _13666_);
  or (_13672_, _13671_, _02144_);
  or (_13673_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_13674_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_13675_, _13674_, _13673_);
  and (_13676_, _13675_, _01954_);
  or (_13677_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_13678_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_13679_, _13678_, _13677_);
  and (_13680_, _13679_, _02150_);
  or (_13681_, _13680_, _13676_);
  or (_13682_, _13681_, _02131_);
  and (_13684_, _13682_, _02077_);
  and (_13685_, _13684_, _13672_);
  or (_13686_, _13685_, _13662_);
  and (_13687_, _13686_, _02065_);
  and (_13688_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_13689_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_13690_, _13689_, _13688_);
  and (_13691_, _13690_, _01954_);
  and (_13692_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_13693_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_13695_, _13693_, _13692_);
  and (_13696_, _13695_, _02150_);
  or (_13697_, _13696_, _13691_);
  or (_13698_, _13697_, _02144_);
  and (_13699_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_13700_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_13701_, _13700_, _13699_);
  and (_13702_, _13701_, _01954_);
  and (_13703_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_13704_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_13706_, _13704_, _13703_);
  and (_13707_, _13706_, _02150_);
  or (_13708_, _13707_, _13702_);
  or (_13709_, _13708_, _02131_);
  and (_13710_, _13709_, _02157_);
  and (_13711_, _13710_, _13698_);
  or (_13712_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_13713_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and (_13714_, _13713_, _02150_);
  and (_13715_, _13714_, _13712_);
  or (_13717_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_13718_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_13719_, _13718_, _01954_);
  and (_13720_, _13719_, _13717_);
  or (_13721_, _13720_, _13715_);
  or (_13722_, _13721_, _02144_);
  or (_13723_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_13724_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and (_13725_, _13724_, _02150_);
  and (_13726_, _13725_, _13723_);
  or (_13728_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_13729_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_13730_, _13729_, _01954_);
  and (_13731_, _13730_, _13728_);
  or (_13732_, _13731_, _13726_);
  or (_13733_, _13732_, _02131_);
  and (_13734_, _13733_, _02077_);
  and (_13735_, _13734_, _13722_);
  or (_13736_, _13735_, _13711_);
  and (_13737_, _13736_, _02194_);
  or (_13739_, _13737_, _13687_);
  and (_13740_, _13739_, _02143_);
  and (_13741_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_13742_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_13743_, _13742_, _13741_);
  and (_13744_, _13743_, _01954_);
  and (_13745_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_13746_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_13747_, _13746_, _13745_);
  and (_13748_, _13747_, _02150_);
  or (_13750_, _13748_, _13744_);
  and (_13751_, _13750_, _02131_);
  and (_13752_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_13753_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_13754_, _13753_, _13752_);
  and (_13755_, _13754_, _01954_);
  and (_13756_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_13757_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_13758_, _13757_, _13756_);
  and (_13759_, _13758_, _02150_);
  or (_13761_, _13759_, _13755_);
  and (_13762_, _13761_, _02144_);
  or (_13763_, _13762_, _13751_);
  and (_13764_, _13763_, _02157_);
  or (_13765_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_13766_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_13767_, _13766_, _02150_);
  and (_13768_, _13767_, _13765_);
  or (_13769_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_13770_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_13772_, _13770_, _01954_);
  and (_13773_, _13772_, _13769_);
  or (_13774_, _13773_, _13768_);
  and (_13775_, _13774_, _02131_);
  or (_13776_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_13777_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_13778_, _13777_, _02150_);
  and (_13779_, _13778_, _13776_);
  or (_13780_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_13781_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_13783_, _13781_, _01954_);
  and (_13784_, _13783_, _13780_);
  or (_13785_, _13784_, _13779_);
  and (_13786_, _13785_, _02144_);
  or (_13787_, _13786_, _13775_);
  and (_13788_, _13787_, _02077_);
  or (_13789_, _13788_, _13764_);
  and (_13790_, _13789_, _02194_);
  and (_13791_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_13792_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_13794_, _13792_, _13791_);
  and (_13795_, _13794_, _01954_);
  and (_13796_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_13797_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_13798_, _13797_, _13796_);
  and (_13799_, _13798_, _02150_);
  or (_13800_, _13799_, _13795_);
  and (_13801_, _13800_, _02131_);
  and (_13802_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_13803_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_13805_, _13803_, _13802_);
  and (_13806_, _13805_, _01954_);
  and (_13807_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and (_13808_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_13809_, _13808_, _13807_);
  and (_13810_, _13809_, _02150_);
  or (_13811_, _13810_, _13806_);
  and (_13812_, _13811_, _02144_);
  or (_13813_, _13812_, _13801_);
  and (_13814_, _13813_, _02157_);
  or (_13816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_13817_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and (_13818_, _13817_, _13816_);
  and (_13819_, _13818_, _01954_);
  or (_13820_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_13821_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_13822_, _13821_, _13820_);
  and (_13823_, _13822_, _02150_);
  or (_13824_, _13823_, _13819_);
  and (_13825_, _13824_, _02131_);
  or (_13827_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_13828_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and (_13829_, _13828_, _13827_);
  and (_13830_, _13829_, _01954_);
  or (_13831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_13832_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_13833_, _13832_, _13831_);
  and (_13834_, _13833_, _02150_);
  or (_13835_, _13834_, _13830_);
  and (_13836_, _13835_, _02144_);
  or (_13837_, _13836_, _13825_);
  and (_13838_, _13837_, _02077_);
  or (_13839_, _13838_, _13814_);
  and (_13840_, _13839_, _02065_);
  or (_13841_, _13840_, _13790_);
  and (_13842_, _13841_, _02005_);
  or (_13843_, _13842_, _13740_);
  or (_13844_, _13843_, _02054_);
  and (_13845_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_13846_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_13847_, _13846_, _13845_);
  and (_13848_, _13847_, _01954_);
  and (_13849_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_13850_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_13851_, _13850_, _13849_);
  and (_13852_, _13851_, _02150_);
  or (_13853_, _13852_, _13848_);
  or (_13854_, _13853_, _02144_);
  and (_13855_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_13856_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_13857_, _13856_, _13855_);
  and (_13858_, _13857_, _01954_);
  and (_13859_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_13860_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_13861_, _13860_, _13859_);
  and (_13862_, _13861_, _02150_);
  or (_13863_, _13862_, _13858_);
  or (_13864_, _13863_, _02131_);
  and (_13865_, _13864_, _02157_);
  and (_13866_, _13865_, _13854_);
  or (_13867_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_13868_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_13869_, _13868_, _02150_);
  and (_13870_, _13869_, _13867_);
  or (_13871_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_13872_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_13873_, _13872_, _01954_);
  and (_13874_, _13873_, _13871_);
  or (_13875_, _13874_, _13870_);
  or (_13876_, _13875_, _02144_);
  or (_13877_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_13878_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and (_13879_, _13878_, _02150_);
  and (_13880_, _13879_, _13877_);
  or (_13881_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_13882_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and (_13883_, _13882_, _01954_);
  and (_13884_, _13883_, _13881_);
  or (_13885_, _13884_, _13880_);
  or (_13886_, _13885_, _02131_);
  and (_13887_, _13886_, _02077_);
  and (_13888_, _13887_, _13876_);
  or (_13889_, _13888_, _13866_);
  and (_13890_, _13889_, _02194_);
  and (_13891_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_13892_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_13893_, _13892_, _13891_);
  and (_13894_, _13893_, _01954_);
  and (_13895_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_13896_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_13897_, _13896_, _13895_);
  and (_13898_, _13897_, _02150_);
  or (_13899_, _13898_, _13894_);
  or (_13900_, _13899_, _02144_);
  and (_13901_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_13902_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_13903_, _13902_, _13901_);
  and (_13904_, _13903_, _01954_);
  and (_13905_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_13906_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_13907_, _13906_, _13905_);
  and (_13908_, _13907_, _02150_);
  or (_13909_, _13908_, _13904_);
  or (_13910_, _13909_, _02131_);
  and (_13911_, _13910_, _02157_);
  and (_13912_, _13911_, _13900_);
  or (_13913_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_13914_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_13915_, _13914_, _13913_);
  and (_13916_, _13915_, _01954_);
  or (_13917_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_13918_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_13919_, _13918_, _13917_);
  and (_13920_, _13919_, _02150_);
  or (_13921_, _13920_, _13916_);
  or (_13922_, _13921_, _02144_);
  or (_13923_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_13924_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_13925_, _13924_, _13923_);
  and (_13926_, _13925_, _01954_);
  or (_13927_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_13928_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_13929_, _13928_, _13927_);
  and (_13930_, _13929_, _02150_);
  or (_13931_, _13930_, _13926_);
  or (_13932_, _13931_, _02131_);
  and (_13933_, _13932_, _02077_);
  and (_13934_, _13933_, _13922_);
  or (_13935_, _13934_, _13912_);
  and (_13936_, _13935_, _02065_);
  or (_13937_, _13936_, _13890_);
  and (_13938_, _13937_, _02143_);
  or (_13939_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_13940_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and (_13941_, _13940_, _13939_);
  and (_13942_, _13941_, _01954_);
  or (_13943_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_13944_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_13945_, _13944_, _13943_);
  and (_13946_, _13945_, _02150_);
  or (_13947_, _13946_, _13942_);
  and (_13948_, _13947_, _02144_);
  or (_13949_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_13950_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_13951_, _13950_, _13949_);
  and (_13952_, _13951_, _01954_);
  or (_13953_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_13954_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_13955_, _13954_, _13953_);
  and (_13956_, _13955_, _02150_);
  or (_13957_, _13956_, _13952_);
  and (_13958_, _13957_, _02131_);
  or (_13959_, _13958_, _13948_);
  and (_13960_, _13959_, _02077_);
  and (_13961_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and (_13962_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_13963_, _13962_, _13961_);
  and (_13964_, _13963_, _01954_);
  and (_13965_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and (_13966_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_13967_, _13966_, _13965_);
  and (_13968_, _13967_, _02150_);
  or (_13969_, _13968_, _13964_);
  and (_13970_, _13969_, _02144_);
  and (_13971_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and (_13972_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_13973_, _13972_, _13971_);
  and (_13974_, _13973_, _01954_);
  and (_13975_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_13976_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_13977_, _13976_, _13975_);
  and (_13978_, _13977_, _02150_);
  or (_13979_, _13978_, _13974_);
  and (_13980_, _13979_, _02131_);
  or (_13981_, _13980_, _13970_);
  and (_13982_, _13981_, _02157_);
  or (_13983_, _13982_, _13960_);
  and (_13984_, _13983_, _02065_);
  or (_13985_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_13986_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_13987_, _13986_, _02150_);
  and (_13988_, _13987_, _13985_);
  or (_13989_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_13990_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_13991_, _13990_, _01954_);
  and (_13992_, _13991_, _13989_);
  or (_13993_, _13992_, _13988_);
  and (_13994_, _13993_, _02144_);
  or (_13995_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_13996_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_13997_, _13996_, _02150_);
  and (_13998_, _13997_, _13995_);
  or (_13999_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_14000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and (_14001_, _14000_, _01954_);
  and (_14002_, _14001_, _13999_);
  or (_14003_, _14002_, _13998_);
  and (_14004_, _14003_, _02131_);
  or (_14005_, _14004_, _13994_);
  and (_14006_, _14005_, _02077_);
  and (_14007_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and (_14008_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_14009_, _14008_, _14007_);
  and (_14010_, _14009_, _01954_);
  and (_14011_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_14012_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_14013_, _14012_, _14011_);
  and (_14014_, _14013_, _02150_);
  or (_14015_, _14014_, _14010_);
  and (_14016_, _14015_, _02144_);
  and (_14017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_14018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_14019_, _14018_, _14017_);
  and (_14020_, _14019_, _01954_);
  and (_14021_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_14022_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_14023_, _14022_, _14021_);
  and (_14024_, _14023_, _02150_);
  or (_14025_, _14024_, _14020_);
  and (_14026_, _14025_, _02131_);
  or (_14027_, _14026_, _14016_);
  and (_14028_, _14027_, _02157_);
  or (_14029_, _14028_, _14006_);
  and (_14030_, _14029_, _02194_);
  or (_14031_, _14030_, _13984_);
  and (_14032_, _14031_, _02005_);
  or (_14033_, _14032_, _13938_);
  or (_14034_, _14033_, _02374_);
  and (_14035_, _14034_, _13844_);
  or (_14036_, _14035_, _02142_);
  and (_14037_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_14038_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_14039_, _14038_, _14037_);
  and (_14040_, _14039_, _01954_);
  and (_14041_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_14042_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_14043_, _14042_, _14041_);
  and (_14044_, _14043_, _02150_);
  or (_14045_, _14044_, _14040_);
  or (_14046_, _14045_, _02144_);
  and (_14047_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_14048_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_14049_, _14048_, _14047_);
  and (_14050_, _14049_, _01954_);
  and (_14051_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_14052_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_14053_, _14052_, _14051_);
  and (_14054_, _14053_, _02150_);
  or (_14055_, _14054_, _14050_);
  or (_14056_, _14055_, _02131_);
  and (_14057_, _14056_, _02157_);
  and (_14058_, _14057_, _14046_);
  or (_14059_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_14060_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_14061_, _14060_, _14059_);
  and (_14062_, _14061_, _01954_);
  or (_14063_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_14064_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_14065_, _14064_, _14063_);
  and (_14066_, _14065_, _02150_);
  or (_14067_, _14066_, _14062_);
  or (_14068_, _14067_, _02144_);
  or (_14069_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_14070_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_14071_, _14070_, _14069_);
  and (_14072_, _14071_, _01954_);
  or (_14073_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_14074_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_14075_, _14074_, _14073_);
  and (_14076_, _14075_, _02150_);
  or (_14077_, _14076_, _14072_);
  or (_14078_, _14077_, _02131_);
  and (_14079_, _14078_, _02077_);
  and (_14080_, _14079_, _14068_);
  or (_14081_, _14080_, _14058_);
  and (_14082_, _14081_, _02065_);
  and (_14083_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_14084_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_14085_, _14084_, _14083_);
  and (_14086_, _14085_, _01954_);
  and (_14087_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_14088_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_14089_, _14088_, _14087_);
  and (_14090_, _14089_, _02150_);
  or (_14091_, _14090_, _14086_);
  or (_14092_, _14091_, _02144_);
  and (_14093_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_14094_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_14095_, _14094_, _14093_);
  and (_14096_, _14095_, _01954_);
  and (_14097_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_14098_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_14099_, _14098_, _14097_);
  and (_14100_, _14099_, _02150_);
  or (_14101_, _14100_, _14096_);
  or (_14102_, _14101_, _02131_);
  and (_14103_, _14102_, _02157_);
  and (_14104_, _14103_, _14092_);
  or (_14105_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_14106_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_14107_, _14106_, _02150_);
  and (_14108_, _14107_, _14105_);
  or (_14109_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_14110_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_14111_, _14110_, _01954_);
  and (_14112_, _14111_, _14109_);
  or (_14113_, _14112_, _14108_);
  or (_14114_, _14113_, _02144_);
  or (_14115_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_14116_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_14117_, _14116_, _02150_);
  and (_14118_, _14117_, _14115_);
  or (_14119_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_14120_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_14121_, _14120_, _01954_);
  and (_14122_, _14121_, _14119_);
  or (_14123_, _14122_, _14118_);
  or (_14124_, _14123_, _02131_);
  and (_14125_, _14124_, _02077_);
  and (_14126_, _14125_, _14114_);
  or (_14127_, _14126_, _14104_);
  and (_14128_, _14127_, _02194_);
  or (_14129_, _14128_, _14082_);
  and (_14130_, _14129_, _02143_);
  and (_14131_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_14132_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_14133_, _14132_, _14131_);
  and (_14134_, _14133_, _01954_);
  and (_14135_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_14136_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_14137_, _14136_, _14135_);
  and (_14138_, _14137_, _02150_);
  or (_14139_, _14138_, _14134_);
  and (_14140_, _14139_, _02131_);
  and (_14141_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_14142_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_14143_, _14142_, _14141_);
  and (_14144_, _14143_, _01954_);
  and (_14145_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_14146_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_14147_, _14146_, _14145_);
  and (_14148_, _14147_, _02150_);
  or (_14149_, _14148_, _14144_);
  and (_14150_, _14149_, _02144_);
  or (_14151_, _14150_, _14140_);
  and (_14152_, _14151_, _02157_);
  or (_14153_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_14154_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_14155_, _14154_, _02150_);
  and (_14156_, _14155_, _14153_);
  or (_14157_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_14158_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_14159_, _14158_, _01954_);
  and (_14160_, _14159_, _14157_);
  or (_14161_, _14160_, _14156_);
  and (_14162_, _14161_, _02131_);
  or (_14163_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_14164_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_14165_, _14164_, _02150_);
  and (_14166_, _14165_, _14163_);
  or (_14167_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_14168_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_14169_, _14168_, _01954_);
  and (_14170_, _14169_, _14167_);
  or (_14171_, _14170_, _14166_);
  and (_14172_, _14171_, _02144_);
  or (_14173_, _14172_, _14162_);
  and (_14174_, _14173_, _02077_);
  or (_14175_, _14174_, _14152_);
  and (_14176_, _14175_, _02194_);
  and (_14177_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_14178_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_14179_, _14178_, _14177_);
  and (_14180_, _14179_, _01954_);
  and (_14181_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_14182_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_14183_, _14182_, _14181_);
  and (_14184_, _14183_, _02150_);
  or (_14185_, _14184_, _14180_);
  and (_14186_, _14185_, _02131_);
  and (_14187_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_14188_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_14189_, _14188_, _14187_);
  and (_14190_, _14189_, _01954_);
  and (_14191_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_14192_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_14193_, _14192_, _14191_);
  and (_14194_, _14193_, _02150_);
  or (_14195_, _14194_, _14190_);
  and (_14196_, _14195_, _02144_);
  or (_14197_, _14196_, _14186_);
  and (_14198_, _14197_, _02157_);
  or (_14199_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_14200_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_14201_, _14200_, _14199_);
  and (_14202_, _14201_, _01954_);
  or (_14203_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_14204_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_14205_, _14204_, _14203_);
  and (_14206_, _14205_, _02150_);
  or (_14207_, _14206_, _14202_);
  and (_14208_, _14207_, _02131_);
  or (_14209_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_14210_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_14211_, _14210_, _14209_);
  and (_14212_, _14211_, _01954_);
  or (_14213_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_14214_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_14215_, _14214_, _14213_);
  and (_14216_, _14215_, _02150_);
  or (_14217_, _14216_, _14212_);
  and (_14218_, _14217_, _02144_);
  or (_14219_, _14218_, _14208_);
  and (_14220_, _14219_, _02077_);
  or (_14221_, _14220_, _14198_);
  and (_14222_, _14221_, _02065_);
  or (_14223_, _14222_, _14176_);
  and (_14224_, _14223_, _02005_);
  or (_14225_, _14224_, _14130_);
  or (_14226_, _14225_, _02054_);
  and (_14227_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_14228_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_14229_, _14228_, _14227_);
  and (_14230_, _14229_, _01954_);
  and (_14231_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_14232_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_14233_, _14232_, _14231_);
  and (_14234_, _14233_, _02150_);
  or (_14235_, _14234_, _14230_);
  or (_14236_, _14235_, _02144_);
  and (_14237_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_14238_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_14239_, _14238_, _14237_);
  and (_14240_, _14239_, _01954_);
  and (_14241_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_14242_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_14243_, _14242_, _14241_);
  and (_14244_, _14243_, _02150_);
  or (_14245_, _14244_, _14240_);
  or (_14246_, _14245_, _02131_);
  and (_14247_, _14246_, _02157_);
  and (_14248_, _14247_, _14236_);
  or (_14249_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_14250_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_14251_, _14250_, _02150_);
  and (_14252_, _14251_, _14249_);
  or (_14253_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_14254_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_14255_, _14254_, _01954_);
  and (_14256_, _14255_, _14253_);
  or (_14257_, _14256_, _14252_);
  or (_14258_, _14257_, _02144_);
  or (_14259_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_14260_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_14261_, _14260_, _02150_);
  and (_14262_, _14261_, _14259_);
  or (_14263_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_14264_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_14265_, _14264_, _01954_);
  and (_14266_, _14265_, _14263_);
  or (_14267_, _14266_, _14262_);
  or (_14268_, _14267_, _02131_);
  and (_14269_, _14268_, _02077_);
  and (_14270_, _14269_, _14258_);
  or (_14271_, _14270_, _14248_);
  and (_14272_, _14271_, _02194_);
  and (_14273_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_14274_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_14275_, _14274_, _14273_);
  and (_14276_, _14275_, _01954_);
  and (_14277_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_14278_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_14279_, _14278_, _14277_);
  and (_14280_, _14279_, _02150_);
  or (_14281_, _14280_, _14276_);
  or (_14282_, _14281_, _02144_);
  and (_14283_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_14284_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_14285_, _14284_, _14283_);
  and (_14286_, _14285_, _01954_);
  and (_14287_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_14288_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_14289_, _14288_, _14287_);
  and (_14290_, _14289_, _02150_);
  or (_14291_, _14290_, _14286_);
  or (_14292_, _14291_, _02131_);
  and (_14293_, _14292_, _02157_);
  and (_14294_, _14293_, _14282_);
  or (_14295_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_14296_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_14297_, _14296_, _14295_);
  and (_14298_, _14297_, _01954_);
  or (_14299_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_14300_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_14301_, _14300_, _14299_);
  and (_14302_, _14301_, _02150_);
  or (_14303_, _14302_, _14298_);
  or (_14304_, _14303_, _02144_);
  or (_14305_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_14306_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_14307_, _14306_, _14305_);
  and (_14308_, _14307_, _01954_);
  or (_14309_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_14310_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_14311_, _14310_, _14309_);
  and (_14312_, _14311_, _02150_);
  or (_14313_, _14312_, _14308_);
  or (_14314_, _14313_, _02131_);
  and (_14315_, _14314_, _02077_);
  and (_14316_, _14315_, _14304_);
  or (_14317_, _14316_, _14294_);
  and (_14318_, _14317_, _02065_);
  or (_14319_, _14318_, _14272_);
  and (_14320_, _14319_, _02143_);
  or (_14321_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_14322_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_14323_, _14322_, _14321_);
  and (_14324_, _14323_, _01954_);
  or (_14325_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_14326_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_14327_, _14326_, _14325_);
  and (_14328_, _14327_, _02150_);
  or (_14329_, _14328_, _14324_);
  and (_14330_, _14329_, _02144_);
  or (_14331_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_14332_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_14333_, _14332_, _14331_);
  and (_14334_, _14333_, _01954_);
  or (_14335_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_14336_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_14337_, _14336_, _14335_);
  and (_14338_, _14337_, _02150_);
  or (_14339_, _14338_, _14334_);
  and (_14340_, _14339_, _02131_);
  or (_14341_, _14340_, _14330_);
  and (_14342_, _14341_, _02077_);
  and (_14343_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_14344_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_14345_, _14344_, _14343_);
  and (_14346_, _14345_, _01954_);
  and (_14347_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_14348_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_14349_, _14348_, _14347_);
  and (_14350_, _14349_, _02150_);
  or (_14351_, _14350_, _14346_);
  and (_14352_, _14351_, _02144_);
  and (_14353_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_14354_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_14355_, _14354_, _14353_);
  and (_14356_, _14355_, _01954_);
  and (_14357_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_14358_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_14359_, _14358_, _14357_);
  and (_14360_, _14359_, _02150_);
  or (_14361_, _14360_, _14356_);
  and (_14362_, _14361_, _02131_);
  or (_14363_, _14362_, _14352_);
  and (_14364_, _14363_, _02157_);
  or (_14365_, _14364_, _14342_);
  and (_14366_, _14365_, _02065_);
  or (_14367_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_14368_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and (_14369_, _14368_, _02150_);
  and (_14370_, _14369_, _14367_);
  or (_14371_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_14372_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and (_14373_, _14372_, _01954_);
  and (_14374_, _14373_, _14371_);
  or (_14375_, _14374_, _14370_);
  and (_14376_, _14375_, _02144_);
  or (_14377_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_14378_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and (_14379_, _14378_, _02150_);
  and (_14380_, _14379_, _14377_);
  or (_14381_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_14382_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and (_14383_, _14382_, _01954_);
  and (_14384_, _14383_, _14381_);
  or (_14385_, _14384_, _14380_);
  and (_14386_, _14385_, _02131_);
  or (_14387_, _14386_, _14376_);
  and (_14388_, _14387_, _02077_);
  and (_14389_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and (_14390_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_14391_, _14390_, _14389_);
  and (_14392_, _14391_, _01954_);
  and (_14393_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and (_14394_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_14395_, _14394_, _14393_);
  and (_14396_, _14395_, _02150_);
  or (_14397_, _14396_, _14392_);
  and (_14398_, _14397_, _02144_);
  and (_14399_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and (_14400_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_14401_, _14400_, _14399_);
  and (_14402_, _14401_, _01954_);
  and (_14403_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and (_14404_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_14405_, _14404_, _14403_);
  and (_14406_, _14405_, _02150_);
  or (_14407_, _14406_, _14402_);
  and (_14408_, _14407_, _02131_);
  or (_14409_, _14408_, _14398_);
  and (_14410_, _14409_, _02157_);
  or (_14411_, _14410_, _14388_);
  and (_14412_, _14411_, _02194_);
  or (_14413_, _14412_, _14366_);
  and (_14414_, _14413_, _02005_);
  or (_14415_, _14414_, _14320_);
  or (_14416_, _14415_, _02374_);
  and (_14417_, _14416_, _14226_);
  or (_14418_, _14417_, _01748_);
  and (_14419_, _14418_, _14036_);
  or (_14420_, _14419_, _02141_);
  or (_14421_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_14422_, _14421_, _27355_);
  and (_15246_, _14422_, _14420_);
  and (_14423_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_14424_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_14425_, _14424_, _14423_);
  and (_14426_, _14425_, _01954_);
  and (_14427_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_14428_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_14429_, _14428_, _14427_);
  and (_14430_, _14429_, _02150_);
  or (_14431_, _14430_, _14426_);
  or (_14432_, _14431_, _02144_);
  and (_14433_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_14434_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_14435_, _14434_, _14433_);
  and (_14436_, _14435_, _01954_);
  and (_14437_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_14438_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_14439_, _14438_, _14437_);
  and (_14440_, _14439_, _02150_);
  or (_14441_, _14440_, _14436_);
  or (_14442_, _14441_, _02131_);
  and (_14443_, _14442_, _02157_);
  and (_14444_, _14443_, _14432_);
  or (_14445_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_14446_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_14447_, _14446_, _14445_);
  and (_14448_, _14447_, _01954_);
  or (_14449_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_14450_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_14451_, _14450_, _14449_);
  and (_14452_, _14451_, _02150_);
  or (_14453_, _14452_, _14448_);
  or (_14454_, _14453_, _02144_);
  or (_14455_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_14456_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and (_14457_, _14456_, _14455_);
  and (_14458_, _14457_, _01954_);
  or (_14459_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_14460_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_14461_, _14460_, _14459_);
  and (_14462_, _14461_, _02150_);
  or (_14463_, _14462_, _14458_);
  or (_14464_, _14463_, _02131_);
  and (_14465_, _14464_, _02077_);
  and (_14466_, _14465_, _14454_);
  or (_14467_, _14466_, _14444_);
  and (_14468_, _14467_, _02065_);
  and (_14469_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_14470_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_14471_, _14470_, _14469_);
  and (_14472_, _14471_, _01954_);
  and (_14473_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_14474_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_14475_, _14474_, _14473_);
  and (_14476_, _14475_, _02150_);
  or (_14477_, _14476_, _14472_);
  or (_14478_, _14477_, _02144_);
  and (_14479_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_14480_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_14481_, _14480_, _14479_);
  and (_14482_, _14481_, _01954_);
  and (_14483_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_14484_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_14485_, _14484_, _14483_);
  and (_14486_, _14485_, _02150_);
  or (_14487_, _14486_, _14482_);
  or (_14488_, _14487_, _02131_);
  and (_14489_, _14488_, _02157_);
  and (_14490_, _14489_, _14478_);
  or (_14491_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_14492_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_14493_, _14492_, _02150_);
  and (_14494_, _14493_, _14491_);
  or (_14495_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_14496_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_14497_, _14496_, _01954_);
  and (_14498_, _14497_, _14495_);
  or (_14499_, _14498_, _14494_);
  or (_14500_, _14499_, _02144_);
  or (_14501_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_14502_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_14503_, _14502_, _02150_);
  and (_14504_, _14503_, _14501_);
  or (_14505_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_14506_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_14507_, _14506_, _01954_);
  and (_14508_, _14507_, _14505_);
  or (_14509_, _14508_, _14504_);
  or (_14510_, _14509_, _02131_);
  and (_14511_, _14510_, _02077_);
  and (_14512_, _14511_, _14500_);
  or (_14513_, _14512_, _14490_);
  and (_14514_, _14513_, _02194_);
  or (_14515_, _14514_, _14468_);
  and (_14516_, _14515_, _02143_);
  and (_14517_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_14518_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_14519_, _14518_, _14517_);
  and (_14520_, _14519_, _01954_);
  and (_14521_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_14522_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_14523_, _14522_, _14521_);
  and (_14524_, _14523_, _02150_);
  or (_14525_, _14524_, _14520_);
  and (_14526_, _14525_, _02131_);
  and (_14527_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_14528_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_14529_, _14528_, _14527_);
  and (_14530_, _14529_, _01954_);
  and (_14531_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_14532_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_14533_, _14532_, _14531_);
  and (_14534_, _14533_, _02150_);
  or (_14535_, _14534_, _14530_);
  and (_14536_, _14535_, _02144_);
  or (_14537_, _14536_, _14526_);
  and (_14538_, _14537_, _02157_);
  or (_14539_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_14540_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_14541_, _14540_, _02150_);
  and (_14542_, _14541_, _14539_);
  or (_14543_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_14544_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_14545_, _14544_, _01954_);
  and (_14546_, _14545_, _14543_);
  or (_14547_, _14546_, _14542_);
  and (_14548_, _14547_, _02131_);
  or (_14549_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_14550_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_14551_, _14550_, _02150_);
  and (_14552_, _14551_, _14549_);
  or (_14553_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_14554_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_14555_, _14554_, _01954_);
  and (_14556_, _14555_, _14553_);
  or (_14557_, _14556_, _14552_);
  and (_14558_, _14557_, _02144_);
  or (_14559_, _14558_, _14548_);
  and (_14560_, _14559_, _02077_);
  or (_14561_, _14560_, _14538_);
  and (_14562_, _14561_, _02194_);
  and (_14563_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and (_14564_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_14565_, _14564_, _14563_);
  and (_14566_, _14565_, _01954_);
  and (_14567_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_14568_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_14569_, _14568_, _14567_);
  and (_14570_, _14569_, _02150_);
  or (_14571_, _14570_, _14566_);
  and (_14572_, _14571_, _02131_);
  and (_14573_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and (_14574_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_14575_, _14574_, _14573_);
  and (_14576_, _14575_, _01954_);
  and (_14577_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and (_14578_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_14579_, _14578_, _14577_);
  and (_14580_, _14579_, _02150_);
  or (_14581_, _14580_, _14576_);
  and (_14582_, _14581_, _02144_);
  or (_14583_, _14582_, _14572_);
  and (_14584_, _14583_, _02157_);
  or (_14585_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_14586_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and (_14587_, _14586_, _14585_);
  and (_14588_, _14587_, _01954_);
  or (_14589_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_14590_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_14591_, _14590_, _14589_);
  and (_14592_, _14591_, _02150_);
  or (_14593_, _14592_, _14588_);
  and (_14594_, _14593_, _02131_);
  or (_14595_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_14596_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and (_14597_, _14596_, _14595_);
  and (_14598_, _14597_, _01954_);
  or (_14599_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_14600_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_14601_, _14600_, _14599_);
  and (_14602_, _14601_, _02150_);
  or (_14603_, _14602_, _14598_);
  and (_14604_, _14603_, _02144_);
  or (_14605_, _14604_, _14594_);
  and (_14606_, _14605_, _02077_);
  or (_14607_, _14606_, _14584_);
  and (_14608_, _14607_, _02065_);
  or (_14609_, _14608_, _14562_);
  and (_14610_, _14609_, _02005_);
  or (_14611_, _14610_, _14516_);
  or (_14612_, _14611_, _02054_);
  and (_14613_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and (_14614_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_14615_, _14614_, _14613_);
  and (_14616_, _14615_, _01954_);
  and (_14617_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_14618_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_14619_, _14618_, _14617_);
  and (_14620_, _14619_, _02150_);
  or (_14621_, _14620_, _14616_);
  or (_14622_, _14621_, _02144_);
  and (_14623_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_14624_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_14625_, _14624_, _14623_);
  and (_14626_, _14625_, _01954_);
  and (_14627_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and (_14628_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_14629_, _14628_, _14627_);
  and (_14630_, _14629_, _02150_);
  or (_14631_, _14630_, _14626_);
  or (_14632_, _14631_, _02131_);
  and (_14633_, _14632_, _02157_);
  and (_14634_, _14633_, _14622_);
  or (_14635_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_14636_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_14637_, _14636_, _02150_);
  and (_14638_, _14637_, _14635_);
  or (_14639_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_14640_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_14641_, _14640_, _01954_);
  and (_14642_, _14641_, _14639_);
  or (_14643_, _14642_, _14638_);
  or (_14644_, _14643_, _02144_);
  or (_14645_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_14646_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_14647_, _14646_, _02150_);
  and (_14648_, _14647_, _14645_);
  or (_14649_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_14650_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_14651_, _14650_, _01954_);
  and (_14652_, _14651_, _14649_);
  or (_14653_, _14652_, _14648_);
  or (_14654_, _14653_, _02131_);
  and (_14655_, _14654_, _02077_);
  and (_14656_, _14655_, _14644_);
  or (_14657_, _14656_, _14634_);
  and (_14658_, _14657_, _02194_);
  and (_14659_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_14660_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_14661_, _14660_, _14659_);
  and (_14662_, _14661_, _01954_);
  and (_14663_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_14664_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_14665_, _14664_, _14663_);
  and (_14666_, _14665_, _02150_);
  or (_14667_, _14666_, _14662_);
  or (_14668_, _14667_, _02144_);
  and (_14669_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_14670_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_14671_, _14670_, _14669_);
  and (_14672_, _14671_, _01954_);
  and (_14673_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_14674_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_14675_, _14674_, _14673_);
  and (_14676_, _14675_, _02150_);
  or (_14677_, _14676_, _14672_);
  or (_14678_, _14677_, _02131_);
  and (_14679_, _14678_, _02157_);
  and (_14680_, _14679_, _14668_);
  or (_14681_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_14682_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_14683_, _14682_, _14681_);
  and (_14684_, _14683_, _01954_);
  or (_14685_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_14686_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_14687_, _14686_, _14685_);
  and (_14688_, _14687_, _02150_);
  or (_14689_, _14688_, _14684_);
  or (_14690_, _14689_, _02144_);
  or (_14691_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_14692_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_14693_, _14692_, _14691_);
  and (_14694_, _14693_, _01954_);
  or (_14695_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_14696_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_14697_, _14696_, _14695_);
  and (_14698_, _14697_, _02150_);
  or (_14699_, _14698_, _14694_);
  or (_14700_, _14699_, _02131_);
  and (_14701_, _14700_, _02077_);
  and (_14702_, _14701_, _14690_);
  or (_14703_, _14702_, _14680_);
  and (_14704_, _14703_, _02065_);
  or (_14705_, _14704_, _14658_);
  and (_14706_, _14705_, _02143_);
  or (_14707_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_14708_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_14709_, _14708_, _14707_);
  and (_14710_, _14709_, _01954_);
  or (_14711_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_14712_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and (_14713_, _14712_, _14711_);
  and (_14714_, _14713_, _02150_);
  or (_14715_, _14714_, _14710_);
  and (_14716_, _14715_, _02144_);
  or (_14717_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_14718_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_14719_, _14718_, _14717_);
  and (_14720_, _14719_, _01954_);
  or (_14721_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_14722_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_14723_, _14722_, _14721_);
  and (_14724_, _14723_, _02150_);
  or (_14725_, _14724_, _14720_);
  and (_14726_, _14725_, _02131_);
  or (_14727_, _14726_, _14716_);
  and (_14728_, _14727_, _02077_);
  and (_14729_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_14730_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_14731_, _14730_, _14729_);
  and (_14732_, _14731_, _01954_);
  and (_14733_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_14734_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_14735_, _14734_, _14733_);
  and (_14736_, _14735_, _02150_);
  or (_14737_, _14736_, _14732_);
  and (_14738_, _14737_, _02144_);
  and (_14739_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_14740_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_14741_, _14740_, _14739_);
  and (_14742_, _14741_, _01954_);
  and (_14743_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and (_14744_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_14745_, _14744_, _14743_);
  and (_14746_, _14745_, _02150_);
  or (_14747_, _14746_, _14742_);
  and (_14748_, _14747_, _02131_);
  or (_14749_, _14748_, _14738_);
  and (_14750_, _14749_, _02157_);
  or (_14751_, _14750_, _14728_);
  and (_14752_, _14751_, _02065_);
  or (_14753_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_14754_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and (_14755_, _14754_, _02150_);
  and (_14756_, _14755_, _14753_);
  or (_14757_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_14758_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_14759_, _14758_, _01954_);
  and (_14760_, _14759_, _14757_);
  or (_14761_, _14760_, _14756_);
  and (_14762_, _14761_, _02144_);
  or (_14763_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_14764_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and (_14765_, _14764_, _02150_);
  and (_14766_, _14765_, _14763_);
  or (_14767_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_14768_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and (_14769_, _14768_, _01954_);
  and (_14770_, _14769_, _14767_);
  or (_14771_, _14770_, _14766_);
  and (_14772_, _14771_, _02131_);
  or (_14773_, _14772_, _14762_);
  and (_14774_, _14773_, _02077_);
  and (_14775_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_14776_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_14777_, _14776_, _14775_);
  and (_14778_, _14777_, _01954_);
  and (_14779_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_14780_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_14781_, _14780_, _14779_);
  and (_14782_, _14781_, _02150_);
  or (_14783_, _14782_, _14778_);
  and (_14784_, _14783_, _02144_);
  and (_14785_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_14786_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_14787_, _14786_, _14785_);
  and (_14788_, _14787_, _01954_);
  and (_14789_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_14790_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_14791_, _14790_, _14789_);
  and (_14792_, _14791_, _02150_);
  or (_14793_, _14792_, _14788_);
  and (_14794_, _14793_, _02131_);
  or (_14795_, _14794_, _14784_);
  and (_14796_, _14795_, _02157_);
  or (_14797_, _14796_, _14774_);
  and (_14798_, _14797_, _02194_);
  or (_14799_, _14798_, _14752_);
  and (_14800_, _14799_, _02005_);
  or (_14801_, _14800_, _14706_);
  or (_14802_, _14801_, _02374_);
  and (_14803_, _14802_, _14612_);
  or (_14804_, _14803_, _02142_);
  and (_14805_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_14806_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_14807_, _14806_, _14805_);
  and (_14808_, _14807_, _01954_);
  and (_14809_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_14810_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_14811_, _14810_, _14809_);
  and (_14812_, _14811_, _02150_);
  or (_14813_, _14812_, _14808_);
  or (_14814_, _14813_, _02144_);
  and (_14815_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_14816_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_14817_, _14816_, _14815_);
  and (_14818_, _14817_, _01954_);
  and (_14819_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_14820_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_14821_, _14820_, _14819_);
  and (_14822_, _14821_, _02150_);
  or (_14823_, _14822_, _14818_);
  or (_14824_, _14823_, _02131_);
  and (_14825_, _14824_, _02157_);
  and (_14826_, _14825_, _14814_);
  or (_14827_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_14828_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_14829_, _14828_, _14827_);
  and (_14830_, _14829_, _01954_);
  or (_14831_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_14832_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_14833_, _14832_, _14831_);
  and (_14834_, _14833_, _02150_);
  or (_14835_, _14834_, _14830_);
  or (_14836_, _14835_, _02144_);
  or (_14837_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_14838_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_14839_, _14838_, _14837_);
  and (_14840_, _14839_, _01954_);
  or (_14841_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_14842_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_14843_, _14842_, _14841_);
  and (_14844_, _14843_, _02150_);
  or (_14845_, _14844_, _14840_);
  or (_14846_, _14845_, _02131_);
  and (_14847_, _14846_, _02077_);
  and (_14848_, _14847_, _14836_);
  or (_14849_, _14848_, _14826_);
  and (_14850_, _14849_, _02065_);
  and (_14851_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_14852_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_14853_, _14852_, _14851_);
  and (_14854_, _14853_, _01954_);
  and (_14855_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_14856_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_14857_, _14856_, _14855_);
  and (_14858_, _14857_, _02150_);
  or (_14859_, _14858_, _14854_);
  or (_14860_, _14859_, _02144_);
  and (_14861_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_14862_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_14863_, _14862_, _14861_);
  and (_14864_, _14863_, _01954_);
  and (_14865_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_14866_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_14867_, _14866_, _14865_);
  and (_14868_, _14867_, _02150_);
  or (_14869_, _14868_, _14864_);
  or (_14870_, _14869_, _02131_);
  and (_14871_, _14870_, _02157_);
  and (_14872_, _14871_, _14860_);
  or (_14873_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_14874_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_14875_, _14874_, _02150_);
  and (_14876_, _14875_, _14873_);
  or (_14877_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_14878_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_14879_, _14878_, _01954_);
  and (_14880_, _14879_, _14877_);
  or (_14881_, _14880_, _14876_);
  or (_14882_, _14881_, _02144_);
  or (_14883_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_14884_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_14885_, _14884_, _02150_);
  and (_14886_, _14885_, _14883_);
  or (_14887_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_14888_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_14889_, _14888_, _01954_);
  and (_14890_, _14889_, _14887_);
  or (_14891_, _14890_, _14886_);
  or (_14892_, _14891_, _02131_);
  and (_14893_, _14892_, _02077_);
  and (_14894_, _14893_, _14882_);
  or (_14895_, _14894_, _14872_);
  and (_14896_, _14895_, _02194_);
  or (_14897_, _14896_, _14850_);
  and (_14898_, _14897_, _02143_);
  and (_14899_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_14900_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_14901_, _14900_, _14899_);
  and (_14902_, _14901_, _01954_);
  and (_14903_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_14904_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_14905_, _14904_, _14903_);
  and (_14906_, _14905_, _02150_);
  or (_14907_, _14906_, _14902_);
  and (_14908_, _14907_, _02131_);
  and (_14909_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_14910_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_14911_, _14910_, _14909_);
  and (_14912_, _14911_, _01954_);
  and (_14913_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_14914_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_14915_, _14914_, _14913_);
  and (_14916_, _14915_, _02150_);
  or (_14917_, _14916_, _14912_);
  and (_14918_, _14917_, _02144_);
  or (_14919_, _14918_, _14908_);
  and (_14920_, _14919_, _02157_);
  or (_14921_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_14922_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_14923_, _14922_, _02150_);
  and (_14924_, _14923_, _14921_);
  or (_14925_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_14926_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and (_14927_, _14926_, _01954_);
  and (_14928_, _14927_, _14925_);
  or (_14929_, _14928_, _14924_);
  and (_14930_, _14929_, _02131_);
  or (_14931_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_14932_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and (_14933_, _14932_, _02150_);
  and (_14934_, _14933_, _14931_);
  or (_14935_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_14936_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_14937_, _14936_, _01954_);
  and (_14938_, _14937_, _14935_);
  or (_14939_, _14938_, _14934_);
  and (_14940_, _14939_, _02144_);
  or (_14941_, _14940_, _14930_);
  and (_14942_, _14941_, _02077_);
  or (_14943_, _14942_, _14920_);
  and (_14944_, _14943_, _02194_);
  and (_14945_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_14946_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_14947_, _14946_, _14945_);
  and (_14948_, _14947_, _01954_);
  and (_14949_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_14950_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_14951_, _14950_, _14949_);
  and (_14952_, _14951_, _02150_);
  or (_14953_, _14952_, _14948_);
  and (_14954_, _14953_, _02131_);
  and (_14955_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_14956_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_14957_, _14956_, _14955_);
  and (_14958_, _14957_, _01954_);
  and (_14959_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_14960_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_14961_, _14960_, _14959_);
  and (_14962_, _14961_, _02150_);
  or (_14963_, _14962_, _14958_);
  and (_14964_, _14963_, _02144_);
  or (_14965_, _14964_, _14954_);
  and (_14966_, _14965_, _02157_);
  or (_14967_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_14968_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_14969_, _14968_, _14967_);
  and (_14970_, _14969_, _01954_);
  or (_14971_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_14972_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_14973_, _14972_, _14971_);
  and (_14974_, _14973_, _02150_);
  or (_14975_, _14974_, _14970_);
  and (_14976_, _14975_, _02131_);
  or (_14977_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_14978_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_14979_, _14978_, _14977_);
  and (_14980_, _14979_, _01954_);
  or (_14981_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_14982_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_14983_, _14982_, _14981_);
  and (_14984_, _14983_, _02150_);
  or (_14985_, _14984_, _14980_);
  and (_14986_, _14985_, _02144_);
  or (_14987_, _14986_, _14976_);
  and (_14988_, _14987_, _02077_);
  or (_14989_, _14988_, _14966_);
  and (_14990_, _14989_, _02065_);
  or (_14991_, _14990_, _14944_);
  and (_14992_, _14991_, _02005_);
  or (_14993_, _14992_, _14898_);
  or (_14994_, _14993_, _02054_);
  and (_14995_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_14996_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_14997_, _14996_, _14995_);
  and (_14998_, _14997_, _01954_);
  and (_14999_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_15000_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_15001_, _15000_, _14999_);
  and (_15002_, _15001_, _02150_);
  or (_15003_, _15002_, _14998_);
  or (_15004_, _15003_, _02144_);
  and (_15005_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_15006_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_15007_, _15006_, _15005_);
  and (_15008_, _15007_, _01954_);
  and (_15009_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_15010_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_15011_, _15010_, _15009_);
  and (_15012_, _15011_, _02150_);
  or (_15013_, _15012_, _15008_);
  or (_15014_, _15013_, _02131_);
  and (_15015_, _15014_, _02157_);
  and (_15016_, _15015_, _15004_);
  or (_15017_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_15018_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_15019_, _15018_, _02150_);
  and (_15020_, _15019_, _15017_);
  or (_15021_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_15022_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_15023_, _15022_, _01954_);
  and (_15024_, _15023_, _15021_);
  or (_15025_, _15024_, _15020_);
  or (_15026_, _15025_, _02144_);
  or (_15027_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_15028_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_15029_, _15028_, _02150_);
  and (_15030_, _15029_, _15027_);
  or (_15031_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_15032_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_15033_, _15032_, _01954_);
  and (_15034_, _15033_, _15031_);
  or (_15035_, _15034_, _15030_);
  or (_15036_, _15035_, _02131_);
  and (_15037_, _15036_, _02077_);
  and (_15038_, _15037_, _15026_);
  or (_15039_, _15038_, _15016_);
  and (_15040_, _15039_, _02194_);
  and (_15041_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_15042_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_15043_, _15042_, _15041_);
  and (_15044_, _15043_, _01954_);
  and (_15045_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_15046_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_15047_, _15046_, _15045_);
  and (_15048_, _15047_, _02150_);
  or (_15049_, _15048_, _15044_);
  or (_15050_, _15049_, _02144_);
  and (_15051_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_15052_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_15053_, _15052_, _15051_);
  and (_15054_, _15053_, _01954_);
  and (_15055_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_15056_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_15057_, _15056_, _15055_);
  and (_15058_, _15057_, _02150_);
  or (_15059_, _15058_, _15054_);
  or (_15060_, _15059_, _02131_);
  and (_15061_, _15060_, _02157_);
  and (_15062_, _15061_, _15050_);
  or (_15063_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_15064_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_15065_, _15064_, _15063_);
  and (_15066_, _15065_, _01954_);
  or (_15067_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_15068_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_15069_, _15068_, _15067_);
  and (_15070_, _15069_, _02150_);
  or (_15071_, _15070_, _15066_);
  or (_15072_, _15071_, _02144_);
  or (_15073_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_15074_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_15075_, _15074_, _15073_);
  and (_15076_, _15075_, _01954_);
  or (_15077_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_15078_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_15079_, _15078_, _15077_);
  and (_15080_, _15079_, _02150_);
  or (_15081_, _15080_, _15076_);
  or (_15082_, _15081_, _02131_);
  and (_15083_, _15082_, _02077_);
  and (_15084_, _15083_, _15072_);
  or (_15085_, _15084_, _15062_);
  and (_15086_, _15085_, _02065_);
  or (_15087_, _15086_, _15040_);
  and (_15088_, _15087_, _02143_);
  or (_15089_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_15090_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_15091_, _15090_, _15089_);
  and (_15092_, _15091_, _01954_);
  or (_15093_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_15094_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_15095_, _15094_, _15093_);
  and (_15096_, _15095_, _02150_);
  or (_15097_, _15096_, _15092_);
  and (_15098_, _15097_, _02144_);
  or (_15099_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_15100_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_15101_, _15100_, _15099_);
  and (_15102_, _15101_, _01954_);
  or (_15103_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_15104_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_15105_, _15104_, _15103_);
  and (_15106_, _15105_, _02150_);
  or (_15107_, _15106_, _15102_);
  and (_15108_, _15107_, _02131_);
  or (_15109_, _15108_, _15098_);
  and (_15110_, _15109_, _02077_);
  and (_15111_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_15112_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_15113_, _15112_, _15111_);
  and (_15114_, _15113_, _01954_);
  and (_15115_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_15116_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_15117_, _15116_, _15115_);
  and (_15118_, _15117_, _02150_);
  or (_15119_, _15118_, _15114_);
  and (_15120_, _15119_, _02144_);
  and (_15121_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_15122_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_15123_, _15122_, _15121_);
  and (_15124_, _15123_, _01954_);
  and (_15125_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_15126_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_15127_, _15126_, _15125_);
  and (_15128_, _15127_, _02150_);
  or (_15129_, _15128_, _15124_);
  and (_15130_, _15129_, _02131_);
  or (_15131_, _15130_, _15120_);
  and (_15132_, _15131_, _02157_);
  or (_15133_, _15132_, _15110_);
  and (_15134_, _15133_, _02065_);
  or (_15135_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_15136_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_15137_, _15136_, _02150_);
  and (_15138_, _15137_, _15135_);
  or (_15139_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_15140_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_15141_, _15140_, _01954_);
  and (_15142_, _15141_, _15139_);
  or (_15143_, _15142_, _15138_);
  and (_15144_, _15143_, _02144_);
  or (_15145_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_15146_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_15147_, _15146_, _02150_);
  and (_15148_, _15147_, _15145_);
  or (_15149_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_15150_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_15151_, _15150_, _01954_);
  and (_15152_, _15151_, _15149_);
  or (_15153_, _15152_, _15148_);
  and (_15154_, _15153_, _02131_);
  or (_15155_, _15154_, _15144_);
  and (_15156_, _15155_, _02077_);
  and (_15157_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_15158_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_15159_, _15158_, _15157_);
  and (_15160_, _15159_, _01954_);
  and (_15161_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_15162_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_15163_, _15162_, _15161_);
  and (_15164_, _15163_, _02150_);
  or (_15165_, _15164_, _15160_);
  and (_15166_, _15165_, _02144_);
  and (_15167_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_15168_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_15169_, _15168_, _15167_);
  and (_15170_, _15169_, _01954_);
  and (_15171_, _02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_15172_, _01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_15173_, _15172_, _15171_);
  and (_15174_, _15173_, _02150_);
  or (_15175_, _15174_, _15170_);
  and (_15176_, _15175_, _02131_);
  or (_15177_, _15176_, _15166_);
  and (_15178_, _15177_, _02157_);
  or (_15179_, _15178_, _15156_);
  and (_15180_, _15179_, _02194_);
  or (_15181_, _15180_, _15134_);
  and (_15182_, _15181_, _02005_);
  or (_15183_, _15182_, _15088_);
  or (_15184_, _15183_, _02374_);
  and (_15185_, _15184_, _14994_);
  or (_15186_, _15185_, _01748_);
  and (_15187_, _15186_, _14804_);
  or (_15188_, _15187_, _02141_);
  or (_15189_, _02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_15190_, _15189_, _27355_);
  and (_15248_, _15190_, _15188_);
  and (pc_log_change, _25988_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  nor (_18890_, _26452_, rst);
  and (_15191_, _26350_, _26286_);
  and (_15192_, _15191_, _26269_);
  not (_15193_, _15192_);
  and (_15194_, _26335_, _26413_);
  and (_15195_, _26351_, _26155_);
  nor (_15196_, _15195_, _15194_);
  and (_15197_, _15196_, _15193_);
  and (_15198_, _26350_, _26181_);
  or (_15199_, _26286_, _26155_);
  nand (_15200_, _15199_, _15198_);
  and (_15201_, _15200_, _15197_);
  and (_15202_, _25987_, _27355_);
  not (_15203_, _15202_);
  or (_15204_, _15203_, _15194_);
  or (_18893_, _15204_, _15201_);
  not (_15205_, _26121_);
  nor (_15206_, _15205_, _26079_);
  and (_15207_, _15206_, _26149_);
  and (_15208_, _15207_, _26028_);
  nor (_15209_, _26259_, _26204_);
  not (_15210_, _26177_);
  nor (_15211_, _26232_, _15210_);
  and (_15212_, _15211_, _15209_);
  and (_15213_, _15212_, _15208_);
  and (_15214_, _26232_, _26177_);
  and (_15215_, _26259_, _26204_);
  and (_15216_, _15215_, _15214_);
  and (_15217_, _15216_, _15207_);
  nor (_15218_, _26149_, _26079_);
  and (_15219_, _15218_, _15205_);
  not (_15220_, _26204_);
  nor (_15221_, _26259_, _15220_);
  and (_15223_, _15221_, _15214_);
  and (_15224_, _15223_, _15219_);
  and (_15225_, _26149_, _15205_);
  or (_15226_, _15225_, _26079_);
  and (_15227_, _15226_, _15223_);
  or (_15228_, _15227_, _15224_);
  or (_15229_, _15228_, _15217_);
  or (_15230_, _15229_, _15213_);
  not (_15231_, _26232_);
  and (_15232_, _15209_, _15231_);
  and (_15233_, _15232_, _15208_);
  and (_15234_, _15233_, _15210_);
  and (_15235_, _15209_, _26232_);
  and (_15237_, _15235_, _15208_);
  and (_15239_, _15221_, _15231_);
  not (_15241_, _26028_);
  and (_15243_, _15207_, _15241_);
  and (_15245_, _15243_, _15239_);
  or (_15247_, _15245_, _15237_);
  or (_15249_, _15247_, _15234_);
  or (_15250_, _15249_, _15230_);
  and (_15251_, _26232_, _15210_);
  and (_15252_, _26259_, _15220_);
  and (_15253_, _15252_, _15251_);
  nor (_15254_, _15253_, _15241_);
  not (_15255_, _26149_);
  and (_15256_, _15206_, _15255_);
  not (_15257_, _15256_);
  nor (_15258_, _15257_, _15254_);
  not (_15259_, _15258_);
  and (_15260_, _15214_, _15209_);
  and (_15261_, _15255_, _26028_);
  and (_15262_, _15261_, _15206_);
  and (_15263_, _15262_, _15260_);
  nor (_15264_, _26232_, _26177_);
  and (_15265_, _15252_, _15264_);
  and (_15266_, _15265_, _15262_);
  nor (_15267_, _15266_, _15263_);
  and (_15268_, _15267_, _15259_);
  and (_15269_, _15252_, _15214_);
  and (_15270_, _15269_, _15243_);
  and (_15271_, _15215_, _15211_);
  and (_15272_, _15219_, _15241_);
  and (_15273_, _15272_, _15271_);
  or (_15274_, _15273_, _15270_);
  and (_15275_, _15252_, _26177_);
  and (_15276_, _15275_, _15262_);
  and (_15277_, _15215_, _26232_);
  and (_15278_, _15262_, _15277_);
  or (_15279_, _15278_, _15276_);
  or (_15280_, _15279_, _15274_);
  and (_15281_, _15251_, _15209_);
  or (_15282_, _15281_, _15212_);
  and (_15283_, _15282_, _15262_);
  and (_15284_, _15271_, _26079_);
  and (_15285_, _15251_, _15215_);
  and (_15286_, _15285_, _15207_);
  or (_15287_, _15286_, _15284_);
  or (_15288_, _15287_, _15283_);
  and (_15289_, _15219_, _26028_);
  and (_15290_, _15221_, _15210_);
  and (_15291_, _15290_, _15289_);
  and (_15292_, _15264_, _15221_);
  and (_15293_, _15262_, _15292_);
  or (_15294_, _15293_, _15291_);
  or (_15295_, _15294_, _15288_);
  nor (_15296_, _15295_, _15280_);
  nand (_15297_, _15296_, _15268_);
  or (_15298_, _15297_, _15250_);
  and (_15299_, _15298_, _25988_);
  not (_15300_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_15301_, _25986_, _23914_);
  and (_15302_, _15301_, _26370_);
  nor (_15303_, _15302_, _15300_);
  or (_15304_, _15303_, rst);
  or (_18896_, _15304_, _15299_);
  not (_15305_, _25982_);
  or (_15306_, _26204_, _15305_);
  or (_15307_, _25982_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_15308_, _15307_, _27355_);
  and (_18899_, _15308_, _15306_);
  and (_15309_, \oc8051_top_1.oc8051_sfr1.wait_data , _27355_);
  and (_15310_, _15309_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_15311_, _26272_, _26413_);
  or (_15312_, _26306_, _26274_);
  or (_15313_, _15312_, _15311_);
  and (_15314_, _26438_, _26351_);
  and (_15315_, _15194_, _26269_);
  or (_15316_, _15315_, _15314_);
  and (_15317_, _26336_, _26286_);
  nor (_15318_, _15317_, _26375_);
  not (_15319_, _15318_);
  or (_15320_, _15319_, _15316_);
  or (_15321_, _15320_, _15313_);
  or (_15322_, _15321_, _26318_);
  and (_15323_, _15322_, _15202_);
  or (_18902_, _15323_, _15310_);
  and (_15324_, _26359_, _26286_);
  or (_15325_, _15324_, _26414_);
  nor (_15326_, _26181_, _26087_);
  and (_15327_, _15326_, _26271_);
  or (_15328_, _15327_, _26405_);
  and (_15329_, _26277_, _26278_);
  and (_15330_, _15329_, _26272_);
  or (_15331_, _15330_, _15328_);
  or (_15332_, _15331_, _15325_);
  and (_15333_, _15332_, _25987_);
  and (_15334_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15335_, _26382_, _15300_);
  not (_15336_, _26441_);
  and (_15337_, _15336_, _15335_);
  or (_15338_, _15337_, _15334_);
  or (_15339_, _15338_, _15333_);
  and (_18905_, _15339_, _27355_);
  and (_15340_, _15309_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15341_, _26438_, _26320_);
  not (_15342_, _26280_);
  nor (_15343_, _26320_, _26289_);
  nor (_15344_, _15343_, _15342_);
  or (_15345_, _15344_, _15341_);
  and (_15346_, _15329_, _26294_);
  or (_15347_, _15346_, _15345_);
  not (_15348_, _26400_);
  nor (_15349_, _15343_, _26087_);
  nor (_15350_, _26269_, _26087_);
  and (_15351_, _15350_, _26293_);
  or (_15352_, _15351_, _15349_);
  or (_15353_, _15352_, _15348_);
  and (_15354_, _26438_, _26362_);
  and (_15355_, _15350_, _26265_);
  or (_15356_, _15355_, _15325_);
  or (_15357_, _15356_, _15354_);
  or (_15358_, _15357_, _15353_);
  or (_15359_, _15358_, _15347_);
  and (_15360_, _15359_, _15202_);
  or (_18908_, _15360_, _15340_);
  and (_15361_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15362_, _26357_, _25987_);
  or (_15363_, _15362_, _15361_);
  or (_15364_, _15363_, _15337_);
  and (_18911_, _15364_, _27355_);
  not (_15365_, _15197_);
  and (_15366_, _15365_, _15335_);
  or (_15367_, _15366_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15368_, _26279_, _26284_);
  and (_15369_, _15368_, _26181_);
  and (_15370_, _26087_, _26034_);
  and (_15371_, _15370_, _26154_);
  and (_15372_, _26294_, _15371_);
  or (_15373_, _15372_, _15369_);
  and (_15374_, _15373_, _26372_);
  or (_15375_, _15374_, _25983_);
  and (_15376_, _26293_, _26273_);
  nor (_15377_, _15376_, _15368_);
  nor (_15378_, _15377_, _26269_);
  or (_15379_, _15378_, _15315_);
  and (_15380_, _15379_, _15375_);
  or (_15381_, _15380_, _15367_);
  or (_15382_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _23914_);
  and (_15383_, _15382_, _27355_);
  and (_18914_, _15383_, _15381_);
  and (_15384_, _15309_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_15385_, _15327_, _26348_);
  or (_15386_, _26309_, _26306_);
  or (_15387_, _15386_, _26268_);
  or (_15388_, _15387_, _15385_);
  and (_15389_, _15350_, _26271_);
  or (_15390_, _15389_, _15351_);
  or (_15391_, _26414_, _26290_);
  or (_15392_, _15391_, _15390_);
  and (_15393_, _26326_, _26294_);
  and (_15394_, _26326_, _26272_);
  or (_15395_, _15394_, _15346_);
  or (_15396_, _15395_, _15393_);
  or (_15397_, _15396_, _15392_);
  or (_15398_, _15397_, _15388_);
  and (_15399_, _15398_, _15202_);
  or (_18917_, _15399_, _15384_);
  and (_15400_, _15309_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_15401_, _15329_, _26341_);
  and (_15402_, _26263_, _26208_);
  and (_15403_, _15402_, _26413_);
  or (_15404_, _15403_, _15330_);
  or (_15405_, _15404_, _15401_);
  or (_15406_, _15405_, _15352_);
  not (_15407_, _26302_);
  and (_15408_, _26438_, _26282_);
  or (_15409_, _15408_, _15407_);
  and (_15410_, _26326_, _26289_);
  not (_15411_, _26425_);
  and (_15412_, _26327_, _26270_);
  or (_15413_, _15412_, _15411_);
  or (_15414_, _15413_, _15410_);
  or (_15415_, _15414_, _15409_);
  or (_15416_, _15415_, _15406_);
  and (_15417_, _15326_, _26270_);
  and (_15418_, _15326_, _26298_);
  or (_15419_, _15418_, _15417_);
  nor (_15420_, _26399_, _26342_);
  not (_15421_, _15420_);
  or (_15422_, _15421_, _26288_);
  or (_15423_, _15422_, _15419_);
  or (_15424_, _15423_, _15347_);
  or (_15425_, _15424_, _15416_);
  and (_15426_, _15425_, _15202_);
  or (_18920_, _15426_, _15400_);
  and (_15427_, _15350_, _26335_);
  and (_15428_, _15329_, _26311_);
  or (_15429_, _15428_, _26403_);
  or (_15430_, _15429_, _15427_);
  not (_15431_, _26407_);
  and (_15432_, _26311_, _26322_);
  or (_15433_, _15432_, _15431_);
  or (_15434_, _15433_, _15430_);
  and (_15435_, _15329_, _26359_);
  or (_15436_, _15435_, _15434_);
  and (_15437_, _15436_, _25987_);
  nand (_15438_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_15439_, _15438_, _26449_);
  or (_15440_, _15439_, _15437_);
  and (_18923_, _15440_, _27355_);
  not (_15441_, _26361_);
  or (_15442_, _15441_, _26344_);
  or (_15443_, _15442_, _15344_);
  or (_15444_, _26348_, _26307_);
  and (_15445_, _26297_, _26181_);
  and (_15446_, _15445_, _26280_);
  or (_15447_, _15446_, _26301_);
  and (_15448_, _26294_, _26273_);
  or (_15449_, _15448_, _26295_);
  or (_15450_, _15449_, _15447_);
  or (_15451_, _15450_, _26275_);
  or (_15452_, _15451_, _15444_);
  or (_15453_, _15452_, _15443_);
  and (_15454_, _15350_, _26297_);
  or (_15455_, _15454_, _26323_);
  and (_15456_, _15326_, _26335_);
  or (_15457_, _15456_, _15369_);
  or (_15458_, _15457_, _15328_);
  or (_15459_, _15458_, _15455_);
  and (_15460_, _15445_, _26326_);
  nor (_15461_, _15460_, _26399_);
  nand (_15462_, _15461_, _26328_);
  or (_15463_, _26420_, _26334_);
  or (_15464_, _15463_, _15462_);
  or (_15465_, _15464_, _15459_);
  or (_15466_, _15465_, _15352_);
  or (_15467_, _15466_, _15453_);
  and (_15468_, _15467_, _25987_);
  and (_15469_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15470_, _26372_, _26316_);
  or (_15471_, _15374_, _15337_);
  or (_15472_, _15471_, _15470_);
  or (_15473_, _15472_, _15469_);
  or (_15474_, _15473_, _15468_);
  and (_18926_, _15474_, _27355_);
  nor (_18984_, _26434_, rst);
  and (_18986_, _26387_, _27355_);
  or (_18989_, _15203_, _15197_);
  nor (_15475_, _15194_, _15191_);
  or (_18992_, _15475_, _15203_);
  or (_15476_, _15291_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_15477_, _15476_, _15247_);
  and (_15478_, _15477_, _15302_);
  nor (_15479_, _15301_, _26370_);
  or (_15480_, _15479_, rst);
  or (_18995_, _15480_, _15478_);
  nand (_15481_, _26028_, _25982_);
  or (_15482_, _25982_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_15483_, _15482_, _27355_);
  and (_18998_, _15483_, _15481_);
  or (_15484_, _26149_, _15305_);
  or (_15485_, _25982_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_15486_, _15485_, _27355_);
  and (_19001_, _15486_, _15484_);
  nand (_15487_, _26121_, _25982_);
  or (_15488_, _25982_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_15489_, _15488_, _27355_);
  and (_19004_, _15489_, _15487_);
  or (_15490_, _26079_, _15305_);
  or (_15491_, _25982_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_15492_, _15491_, _27355_);
  and (_19007_, _15492_, _15490_);
  or (_15493_, _26177_, _15305_);
  or (_15494_, _25982_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_15495_, _15494_, _27355_);
  and (_19010_, _15495_, _15493_);
  or (_15496_, _26232_, _15305_);
  or (_15497_, _25982_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_15498_, _15497_, _27355_);
  and (_19013_, _15498_, _15496_);
  or (_15499_, _26259_, _15305_);
  or (_15500_, _25982_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_15501_, _15500_, _27355_);
  and (_19016_, _15501_, _15499_);
  or (_15502_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _23914_);
  and (_15503_, _15502_, _27355_);
  and (_15504_, _15503_, _15367_);
  and (_15505_, _26438_, _26294_);
  and (_15506_, _26438_, _26289_);
  or (_15507_, _15506_, _15505_);
  or (_15508_, _15507_, _15341_);
  and (_15509_, _15350_, _26281_);
  or (_15510_, _15509_, _15432_);
  and (_15511_, _15329_, _26282_);
  or (_15512_, _15511_, _15324_);
  or (_15513_, _15512_, _15510_);
  or (_15514_, _15513_, _15508_);
  nor (_15515_, _15418_, _15431_);
  nand (_15516_, _15515_, _26426_);
  or (_15517_, _15403_, _26414_);
  or (_15518_, _15517_, _15430_);
  or (_15519_, _15518_, _15516_);
  not (_15520_, _15326_);
  nor (_15521_, _26423_, _15520_);
  and (_15522_, _15329_, _26351_);
  or (_15523_, _15522_, _15521_);
  and (_15524_, _15198_, _26438_);
  and (_15525_, _26333_, _26326_);
  or (_15526_, _15525_, _15524_);
  or (_15527_, _15526_, _15523_);
  or (_15528_, _15435_, _15401_);
  and (_15529_, _26438_, _26299_);
  and (_15530_, _15329_, _26333_);
  or (_15531_, _15530_, _15529_);
  or (_15532_, _15531_, _15528_);
  or (_15533_, _15532_, _15527_);
  or (_15534_, _15533_, _15519_);
  or (_15535_, _15534_, _15514_);
  and (_15536_, _15535_, _15202_);
  or (_19019_, _15536_, _15504_);
  and (_15537_, _15309_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_15538_, _26438_, _26339_);
  nor (_15539_, _15355_, _26398_);
  or (_15540_, _26341_, _26282_);
  nand (_15541_, _15540_, _26273_);
  nand (_15542_, _15541_, _15539_);
  or (_15543_, _15542_, _15538_);
  or (_15544_, _15354_, _15316_);
  or (_15545_, _15512_, _15419_);
  or (_15546_, _15545_, _15544_);
  not (_15547_, _26349_);
  and (_15548_, _26438_, _26341_);
  or (_15549_, _15548_, _15547_);
  or (_15550_, _15549_, _15414_);
  or (_15551_, _15550_, _15546_);
  or (_15552_, _15551_, _15543_);
  and (_15553_, _15552_, _15202_);
  or (_23904_, _15553_, _15537_);
  or (_15554_, _15463_, _15457_);
  or (_15555_, _15554_, _15453_);
  and (_15556_, _15555_, _25987_);
  and (_15557_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15558_, _15557_, _15472_);
  or (_15559_, _15558_, _15556_);
  and (_23905_, _15559_, _27355_);
  and (_15560_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15561_, _15560_, _15471_);
  and (_15562_, _15561_, _27355_);
  and (_15563_, _26343_, _26269_);
  or (_15564_, _15563_, _26405_);
  or (_15565_, _15564_, _15378_);
  or (_15566_, _15565_, _15462_);
  and (_15567_, _15566_, _15202_);
  or (_23906_, _15567_, _15562_);
  and (_15568_, _26438_, _26272_);
  or (_15569_, _15435_, _15568_);
  or (_15570_, _15524_, _26439_);
  and (_15571_, _15329_, _26266_);
  or (_15572_, _15571_, _15314_);
  or (_15573_, _15572_, _15570_);
  or (_15574_, _15573_, _15508_);
  or (_15575_, _15574_, _15569_);
  or (_15576_, _15408_, _15431_);
  or (_15577_, _15529_, _15548_);
  or (_15578_, _15577_, _15576_);
  nor (_15579_, _15460_, _15454_);
  nand (_15580_, _15579_, _26417_);
  or (_15581_, _15580_, _15378_);
  or (_15582_, _15581_, _15578_);
  or (_15583_, _15194_, _26440_);
  and (_15584_, _15428_, _26181_);
  or (_15585_, _15584_, _15530_);
  or (_15586_, _15585_, _15583_);
  and (_15587_, _26333_, _26273_);
  and (_15588_, _15198_, _26280_);
  and (_15589_, _15428_, _26269_);
  or (_15590_, _15589_, _15588_);
  or (_15591_, _15590_, _15587_);
  or (_15592_, _15591_, _15586_);
  or (_15593_, _15427_, _26404_);
  or (_15594_, _15510_, _15403_);
  or (_15595_, _15594_, _15593_);
  or (_15596_, _15595_, _15592_);
  or (_15597_, _15596_, _15582_);
  or (_15598_, _15597_, _15575_);
  and (_15599_, _15598_, _25987_);
  and (_15600_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15601_, _15366_, _26450_);
  or (_15602_, _15601_, _15600_);
  or (_15603_, _15602_, _15599_);
  and (_23907_, _15603_, _27355_);
  and (_15604_, _15350_, _26350_);
  nor (_15605_, _15604_, _15446_);
  and (_15606_, _15605_, _26407_);
  nand (_15607_, _15606_, _26418_);
  and (_15608_, _15540_, _26413_);
  or (_15609_, _15608_, _26340_);
  or (_15610_, _15609_, _15607_);
  or (_15611_, _26440_, _26334_);
  and (_15612_, _15198_, _26326_);
  or (_15613_, _15612_, _15324_);
  or (_15614_, _15613_, _15611_);
  or (_15615_, _15614_, _15594_);
  or (_15616_, _15615_, _15593_);
  or (_15617_, _15616_, _15610_);
  or (_15618_, _15617_, _15575_);
  and (_15619_, _15618_, _25987_);
  and (_15620_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15621_, _15620_, _15601_);
  or (_15622_, _15621_, _15619_);
  and (_23908_, _15622_, _27355_);
  and (_15623_, _15309_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_15624_, _26312_, _26413_);
  or (_15625_, _15584_, _15624_);
  and (_15626_, _26397_, _26311_);
  and (_15627_, _15350_, _26264_);
  and (_15628_, _15627_, _26208_);
  or (_15629_, _15628_, _15626_);
  or (_15630_, _15629_, _15625_);
  or (_15631_, _15630_, _15392_);
  or (_15632_, _15435_, _01750_);
  or (_15633_, _15632_, _15444_);
  or (_15634_, _15633_, _15631_);
  or (_15635_, _15506_, _15346_);
  and (_15636_, _26289_, _26413_);
  and (_15637_, _26294_, _26413_);
  or (_15638_, _15637_, _15636_);
  or (_15639_, _15427_, _15327_);
  or (_15640_, _15639_, _15638_);
  or (_15641_, _15640_, _15635_);
  nand (_15642_, _26407_, _26360_);
  or (_15643_, _15394_, _15393_);
  or (_15644_, _15643_, _15642_);
  and (_15645_, _26266_, _26413_);
  or (_15646_, _15645_, _01753_);
  or (_15647_, _15646_, _15644_);
  or (_15648_, _15647_, _15641_);
  or (_15649_, _15648_, _15634_);
  and (_15650_, _15649_, _15202_);
  or (_23909_, _15650_, _15623_);
  or (_15651_, _15589_, _15410_);
  or (_15652_, _15651_, _15637_);
  or (_15653_, _15652_, _15409_);
  or (_15654_, _15653_, _15586_);
  or (_15655_, _15506_, _15624_);
  not (_15656_, _26338_);
  or (_15657_, _15510_, _15656_);
  or (_15658_, _15657_, _15655_);
  not (_15659_, _26417_);
  or (_15660_, _15659_, _26283_);
  or (_15661_, _15412_, _15330_);
  or (_15662_, _15661_, _15660_);
  or (_15663_, _15417_, _26414_);
  or (_15664_, _15663_, _26404_);
  or (_15665_, _15664_, _15662_);
  or (_15666_, _15665_, _15658_);
  or (_15667_, _15666_, _15654_);
  and (_15668_, _15667_, _15202_);
  and (_15669_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15670_, _26440_, _26393_);
  or (_15671_, _15670_, _15669_);
  and (_15672_, _15671_, _27355_);
  or (_23910_, _15672_, _15668_);
  nor (_15673_, _15530_, _15656_);
  or (_15674_, _15435_, _15314_);
  or (_15675_, _15674_, _15571_);
  and (_15676_, _26311_, _26413_);
  or (_15677_, _15676_, _01752_);
  or (_15678_, _15355_, _15330_);
  or (_15679_, _15678_, _15677_);
  nor (_15680_, _15679_, _15675_);
  nand (_15681_, _15680_, _15673_);
  or (_15682_, _15639_, _26409_);
  or (_15683_, _15524_, _26267_);
  or (_15684_, _15509_, _26402_);
  or (_15685_, _15684_, _15683_);
  or (_15686_, _15685_, _15682_);
  or (_15687_, _15686_, _15353_);
  or (_15688_, _15687_, _15347_);
  or (_15689_, _15688_, _15681_);
  and (_15690_, _15689_, _25987_);
  and (_15691_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15692_, _15691_, _26447_);
  or (_15693_, _15692_, _15690_);
  and (_23911_, _15693_, _27355_);
  or (_15694_, _15683_, _15635_);
  or (_15695_, _15694_, _15684_);
  and (_15696_, _26293_, _26413_);
  or (_15697_, _26405_, _26399_);
  or (_15698_, _15697_, _15696_);
  or (_15699_, _15530_, _26334_);
  or (_15700_, _15699_, _15698_);
  or (_15701_, _15385_, _01750_);
  or (_15702_, _15701_, _15700_);
  or (_15703_, _15352_, _15345_);
  or (_15704_, _15703_, _15702_);
  or (_15705_, _15704_, _15695_);
  and (_15706_, _15705_, _25987_);
  and (_15707_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15708_, _15707_, _26448_);
  or (_15709_, _15708_, _15706_);
  and (_23912_, _15709_, _27355_);
  and (_15710_, _15309_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_15711_, _15655_, _15638_);
  or (_15712_, _15711_, _15646_);
  not (_15713_, _26284_);
  and (_15714_, _26266_, _15713_);
  or (_15715_, _15311_, _26309_);
  or (_15716_, _15715_, _15714_);
  or (_15717_, _15716_, _15434_);
  or (_15718_, _15717_, _15632_);
  or (_15719_, _15718_, _15712_);
  and (_15720_, _15719_, _15202_);
  or (_23913_, _15720_, _15710_);
  and (_24306_, _26204_, _27355_);
  nor (_24307_, _01743_, rst);
  and (_15721_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_15722_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_15723_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_15724_, _26002_, _26193_);
  nor (_15725_, _15724_, _15723_);
  nor (_15726_, _25996_, _01735_);
  and (_15727_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_15728_, _15727_, _15726_);
  not (_15729_, _26009_);
  and (_15730_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_15731_, _26018_, _26190_);
  nor (_15732_, _15731_, _15730_);
  and (_15733_, _15732_, _15728_);
  and (_15734_, _15733_, _15725_);
  nor (_15735_, _15734_, _25992_);
  nor (_15736_, _15735_, _15722_);
  nor (_15737_, _15736_, _01726_);
  nor (_15738_, _15737_, _15721_);
  nor (_24308_, _15738_, rst);
  nor (_24320_, _26028_, rst);
  and (_24321_, _26149_, _27355_);
  nor (_24322_, _26121_, rst);
  and (_24323_, _26079_, _27355_);
  and (_24324_, _26177_, _27355_);
  and (_24325_, _26232_, _27355_);
  and (_24327_, _26259_, _27355_);
  nor (_24328_, _01847_, rst);
  nor (_24329_, _01947_, rst);
  nor (_24330_, _02124_, rst);
  nor (_24331_, _01806_, rst);
  nor (_24333_, _01902_, rst);
  nor (_24334_, _01980_, rst);
  nor (_24335_, _02047_, rst);
  and (_15739_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_15740_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_15741_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor (_15742_, _26002_, _25994_);
  nor (_15743_, _15742_, _15741_);
  nor (_15744_, _25996_, _01841_);
  and (_15745_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_15746_, _15745_, _15744_);
  and (_15747_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_15748_, _26018_, _26008_);
  nor (_15749_, _15748_, _15747_);
  and (_15750_, _15749_, _15746_);
  and (_15751_, _15750_, _15743_);
  nor (_15752_, _15751_, _25992_);
  nor (_15753_, _15752_, _15740_);
  nor (_15754_, _15753_, _01726_);
  nor (_15755_, _15754_, _15739_);
  nor (_24336_, _15755_, rst);
  and (_15756_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_15757_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  nor (_15758_, _25996_, _01935_);
  nor (_15759_, _26002_, _26129_);
  nor (_15760_, _15759_, _15758_);
  and (_15761_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor (_15762_, _26018_, _26127_);
  nor (_15763_, _15762_, _15761_);
  and (_15764_, _15763_, _15760_);
  and (_15765_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_15766_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_15767_, _15766_, _15765_);
  and (_15768_, _15767_, _15764_);
  nor (_15769_, _15768_, _25992_);
  nor (_15770_, _15769_, _15757_);
  nor (_15771_, _15770_, _01726_);
  nor (_15772_, _15771_, _15756_);
  nor (_24337_, _15772_, rst);
  and (_15773_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_15774_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  nor (_15775_, _25996_, _02112_);
  nor (_15776_, _26002_, _26111_);
  nor (_15777_, _15776_, _15775_);
  and (_15778_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_15779_, _26018_, _26105_);
  nor (_15780_, _15779_, _15778_);
  and (_15781_, _15780_, _15777_);
  and (_15782_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_15783_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_15784_, _15783_, _15782_);
  and (_15785_, _15784_, _15781_);
  nor (_15786_, _15785_, _25992_);
  nor (_15787_, _15786_, _15774_);
  nor (_15788_, _15787_, _01726_);
  nor (_15789_, _15788_, _15773_);
  nor (_24339_, _15789_, rst);
  and (_15790_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_15791_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_15792_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor (_15793_, _26002_, _26057_);
  nor (_15794_, _15793_, _15792_);
  nor (_15795_, _25996_, _01794_);
  and (_15796_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_15797_, _15796_, _15795_);
  and (_15798_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_15799_, _26018_, _26051_);
  nor (_15800_, _15799_, _15798_);
  and (_15801_, _15800_, _15797_);
  and (_15802_, _15801_, _15794_);
  nor (_15803_, _15802_, _25992_);
  nor (_15804_, _15803_, _15791_);
  nor (_15805_, _15804_, _01726_);
  nor (_15806_, _15805_, _15790_);
  nor (_24340_, _15806_, rst);
  and (_15807_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_15808_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  nor (_15809_, _25996_, _01892_);
  nor (_15810_, _26002_, _26159_);
  nor (_15811_, _15810_, _15809_);
  and (_15812_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_15813_, _26018_, _26157_);
  nor (_15814_, _15813_, _15812_);
  and (_15815_, _15814_, _15811_);
  and (_15816_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_15817_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_15818_, _15817_, _15816_);
  and (_15819_, _15818_, _15815_);
  nor (_15820_, _15819_, _25992_);
  nor (_15821_, _15820_, _15808_);
  nor (_15822_, _15821_, _01726_);
  nor (_15823_, _15822_, _15807_);
  nor (_24341_, _15823_, rst);
  and (_15824_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_15825_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_15826_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_15827_, _26002_, _26212_);
  nor (_15828_, _15827_, _15826_);
  nor (_15829_, _25996_, _01971_);
  and (_15830_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_15831_, _15830_, _15829_);
  and (_15832_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_15833_, _26018_, _26218_);
  nor (_15834_, _15833_, _15832_);
  and (_15835_, _15834_, _15831_);
  and (_15836_, _15835_, _15828_);
  nor (_15837_, _15836_, _25992_);
  nor (_15838_, _15837_, _15825_);
  nor (_15839_, _15838_, _01726_);
  nor (_15840_, _15839_, _15824_);
  nor (_24342_, _15840_, rst);
  and (_15841_, _01726_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_15842_, _25992_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_15843_, _15729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_15844_, _26013_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_15845_, _15844_, _15843_);
  and (_15846_, _26006_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor (_15847_, _26018_, _26251_);
  nor (_15848_, _15847_, _15846_);
  nor (_15849_, _26002_, _26245_);
  nor (_15850_, _25996_, _02035_);
  nor (_15851_, _15850_, _15849_);
  and (_15852_, _15851_, _15848_);
  and (_15853_, _15852_, _15845_);
  nor (_15854_, _15853_, _25992_);
  nor (_15855_, _15854_, _15842_);
  nor (_15856_, _15855_, _01726_);
  nor (_15857_, _15856_, _15841_);
  nor (_24343_, _15857_, rst);
  and (_15858_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_15859_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_15860_, pc_log_change, _15859_);
  or (_15861_, _15860_, _15858_);
  and (_24370_, _15861_, _27355_);
  or (_15862_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand (_15863_, pc_log_change, _15859_);
  and (_15864_, _15863_, _27355_);
  and (_24372_, _15864_, _15862_);
  nor (_24404_, _01748_, rst);
  nor (_24405_, _01639_, rst);
  and (_24406_, _01721_, _27355_);
  and (_15865_, _26383_, _26353_);
  not (_15866_, _15865_);
  nor (_15867_, _02004_, _26922_);
  and (_15868_, _02004_, _26922_);
  nor (_15869_, _15868_, _15867_);
  nor (_15870_, _01907_, _01637_);
  and (_15871_, _01907_, _01637_);
  nor (_15872_, _15871_, _15870_);
  and (_15873_, _15872_, _15869_);
  nor (_15874_, _01811_, _25116_);
  and (_15875_, _01811_, _25116_);
  nor (_15876_, _15875_, _15874_);
  nor (_15877_, _02053_, _26458_);
  and (_15878_, _02053_, _26458_);
  nor (_15879_, _15878_, _15877_);
  and (_15880_, _15879_, _02062_);
  and (_15881_, _15880_, _15876_);
  and (_15882_, _15881_, _15873_);
  nor (_15883_, _01854_, _25053_);
  and (_15884_, _01854_, _25053_);
  nor (_15885_, _15884_, _15883_);
  nor (_15886_, _15885_, _27160_);
  and (_15887_, _01952_, _25714_);
  nor (_15888_, _01952_, _25714_);
  or (_15889_, _15888_, _15887_);
  nor (_15890_, _02129_, _25020_);
  and (_15891_, _02129_, _25020_);
  nor (_15892_, _15891_, _15890_);
  nor (_15893_, _15892_, _15889_);
  and (_15894_, _15893_, _15886_);
  and (_15895_, _15894_, _15882_);
  nor (_15896_, _25101_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_15897_, _15896_, _15895_);
  not (_15898_, _15897_);
  nor (_15899_, _26319_, _26382_);
  nor (_15900_, _25517_, _27575_);
  and (_15901_, _15900_, _15882_);
  and (_15902_, _15901_, _15899_);
  nor (_15903_, _15377_, _26393_);
  nor (_15904_, _15865_, _26372_);
  and (_15905_, _26311_, _15371_);
  or (_15906_, _15317_, _15659_);
  and (_15907_, _15899_, _25193_);
  not (_15908_, _15907_);
  nor (_15909_, _15899_, _26446_);
  and (_15910_, _25675_, _25530_);
  nand (_15911_, _15910_, _25760_);
  nor (_15912_, _15911_, _25792_);
  and (_15913_, _15912_, _25857_);
  and (_15914_, _15913_, _25335_);
  and (_15915_, _15914_, _25918_);
  and (_15916_, _15915_, _15909_);
  and (_15917_, _15916_, _25351_);
  and (_15918_, _26376_, _26291_);
  and (_15919_, _15918_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_15920_, _15919_, _15917_);
  nor (_15921_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_15922_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_15923_, _15922_, _15921_);
  nor (_15924_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_15925_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_15926_, _15925_, _15924_);
  and (_15927_, _15926_, _15923_);
  nand (_15928_, _15927_, _26432_);
  and (_15929_, _15928_, _15920_);
  and (_15930_, _15929_, _15908_);
  not (_15931_, _26286_);
  or (_15932_, _26312_, _26299_);
  nor (_15933_, _15932_, _26333_);
  nor (_15934_, _15933_, _15931_);
  not (_15935_, _15934_);
  or (_15936_, _15571_, _26290_);
  nor (_15937_, _15936_, _15389_);
  and (_15938_, _15937_, _15539_);
  and (_15939_, _15938_, _15935_);
  not (_15940_, _15939_);
  and (_15941_, _15940_, _15930_);
  and (_15942_, _26375_, _26269_);
  nor (_15943_, _15942_, _26317_);
  nor (_15944_, _15943_, _15930_);
  or (_15945_, _15944_, _15941_);
  or (_15946_, _15945_, _15906_);
  nor (_15947_, _15946_, _15905_);
  nor (_15948_, _15947_, _15904_);
  nor (_15949_, _15948_, _15903_);
  not (_15950_, _26446_);
  nor (_15951_, _15899_, _26281_);
  nor (_15952_, _15951_, _15950_);
  nor (_15953_, _26942_, _26933_);
  and (_15954_, _15953_, _26998_);
  not (_15955_, _15954_);
  and (_15956_, _15955_, _15952_);
  and (_15957_, _26446_, _26236_);
  not (_15958_, _27102_);
  and (_15959_, _15958_, _15957_);
  nor (_15960_, _15959_, _15956_);
  not (_15961_, _15960_);
  nor (_15962_, _15961_, _15949_);
  not (_15963_, _15962_);
  nor (_15964_, _15963_, _15902_);
  and (_15965_, _15964_, _15898_);
  and (_15966_, _15965_, _15866_);
  and (_24410_, _15966_, _27355_);
  and (_24411_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _27355_);
  and (_24412_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _27355_);
  and (_15967_, _25995_, _25999_);
  nor (_15968_, _15967_, _01726_);
  nor (_15969_, _15968_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_15970_, _15969_);
  and (_15971_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_15972_, _15971_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_15973_, _15972_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_15974_, _15973_, _15970_);
  and (_15975_, _15974_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_15976_, _15975_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_15977_, _15976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_15978_, _15977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_15979_, _15978_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_15980_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_15981_, _15980_, _15979_);
  and (_15982_, _15981_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_15983_, _15982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_15984_, _15983_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_15985_, _15983_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_15986_, _15985_, _15984_);
  or (_15987_, _15986_, _15965_);
  and (_15988_, _15987_, _27355_);
  and (_15989_, _26286_, _25983_);
  and (_15990_, _15989_, _26311_);
  not (_15991_, _15990_);
  nand (_15992_, _15539_, _26319_);
  or (_15993_, _15992_, _15936_);
  nand (_15994_, _15993_, _26372_);
  and (_15995_, _26383_, _15905_);
  and (_15996_, _26293_, _15371_);
  and (_15997_, _15996_, _25983_);
  nor (_15998_, _15997_, _15995_);
  and (_15999_, _15998_, _15994_);
  and (_16000_, _15999_, _15991_);
  and (_16001_, _16000_, _01743_);
  nand (_16002_, _15999_, _15991_);
  and (_16003_, _16002_, _15738_);
  nor (_16004_, _16003_, _16001_);
  and (_16005_, _16004_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_16006_, _16005_);
  nor (_16007_, _16004_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_16008_, _16007_, _16005_);
  not (_16009_, _16008_);
  and (_16010_, _16000_, _02047_);
  and (_16011_, _16002_, _15857_);
  nor (_16012_, _16011_, _16010_);
  and (_16013_, _16012_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_16014_, _16013_);
  nor (_16015_, _16012_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_16016_, _16015_, _16013_);
  and (_16017_, _16000_, _01980_);
  and (_16018_, _16002_, _15840_);
  nor (_16019_, _16018_, _16017_);
  nor (_16020_, _16019_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_16021_, _16019_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_16022_, _16000_, _01902_);
  and (_16023_, _16002_, _15823_);
  nor (_16024_, _16023_, _16022_);
  nand (_16025_, _16024_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_16026_, _16000_, _01806_);
  and (_16027_, _16002_, _15806_);
  nor (_16028_, _16027_, _16026_);
  nor (_16029_, _16028_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_16030_, _16028_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_16031_, _16002_, _02125_);
  not (_16032_, _15789_);
  or (_16033_, _16000_, _16032_);
  and (_16034_, _16033_, _16031_);
  and (_16035_, _16034_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_16036_, _16002_, _01948_);
  not (_16037_, _15772_);
  or (_16038_, _16000_, _16037_);
  and (_16039_, _16038_, _16036_);
  nand (_16040_, _16039_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_16041_, _16040_);
  or (_16042_, _16002_, _01848_);
  not (_16043_, _15755_);
  or (_16044_, _16000_, _16043_);
  and (_16045_, _16044_, _16042_);
  and (_16046_, _16045_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_16047_, _16039_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_16048_, _16047_, _16040_);
  and (_16049_, _16048_, _16046_);
  or (_16050_, _16049_, _16041_);
  not (_16051_, _16035_);
  or (_16052_, _16034_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_16053_, _16052_, _16051_);
  and (_16054_, _16053_, _16050_);
  or (_16055_, _16054_, _16035_);
  nor (_16056_, _16055_, _16030_);
  nor (_16057_, _16056_, _16029_);
  or (_16058_, _16024_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_16059_, _16058_, _16025_);
  nand (_16060_, _16059_, _16057_);
  nand (_16061_, _16060_, _16025_);
  nor (_16062_, _16061_, _16021_);
  nor (_16063_, _16062_, _16020_);
  nand (_16064_, _16063_, _16016_);
  and (_16065_, _16064_, _16014_);
  or (_16066_, _16065_, _16009_);
  and (_16067_, _16066_, _16006_);
  nand (_16068_, _16067_, _24240_);
  or (_16069_, _16068_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_16070_, _16069_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_16071_, _16070_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_16072_, _16071_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_16073_, _16072_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_16074_, _16073_, _24129_);
  nand (_16075_, _16074_, _16004_);
  not (_16076_, _16004_);
  nor (_16077_, _16067_, _24240_);
  and (_16078_, _16077_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_16079_, _16078_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_16080_, _16079_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_16081_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_16082_, _16081_, _16080_);
  nand (_16083_, _16082_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_16084_, _16083_, _16076_);
  nand (_16085_, _16084_, _16075_);
  nand (_16086_, _16085_, _24158_);
  or (_16087_, _16085_, _24158_);
  and (_16088_, _16087_, _16086_);
  not (_16089_, _26372_);
  not (_16090_, _15992_);
  and (_16091_, _15318_, _26417_);
  and (_16092_, _16091_, _15937_);
  and (_16093_, _16092_, _16090_);
  nor (_16094_, _16093_, _16089_);
  nor (_16095_, _16094_, _15990_);
  nor (_16096_, _26417_, _16089_);
  nor (_16097_, _16096_, _15903_);
  not (_16098_, _16097_);
  and (_16099_, _16098_, _16000_);
  nor (_16100_, _16099_, _16095_);
  and (_16101_, _16100_, _16088_);
  and (_16102_, _15895_, _25102_);
  and (_16103_, _16102_, _25444_);
  nor (_16104_, _16103_, _15902_);
  and (_16105_, _15958_, _26432_);
  not (_16106_, _16105_);
  and (_16107_, _15955_, _15918_);
  nor (_16108_, _16107_, _15949_);
  and (_16109_, _16108_, _16106_);
  and (_16110_, _16109_, _16104_);
  and (_16111_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_16112_, _16111_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_16113_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_16114_, _16113_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_16115_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_16116_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_16117_, _16116_, _16115_);
  and (_16118_, _16117_, _16114_);
  and (_16119_, _16118_, _16112_);
  and (_16120_, _16119_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_16121_, _16120_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_16122_, _16121_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_16123_, _16122_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_16124_, _16123_, _24158_);
  or (_16125_, _16123_, _24158_);
  and (_16126_, _16125_, _16124_);
  and (_16127_, _15999_, _15903_);
  and (_16128_, _16127_, _16126_);
  and (_16129_, _15995_, _25441_);
  and (_16130_, _16096_, _26678_);
  and (_16131_, _16097_, _15999_);
  and (_16132_, _16131_, _16095_);
  and (_16133_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_16134_, _15376_, _25983_);
  and (_16135_, _16134_, _01744_);
  or (_16136_, _16135_, _16133_);
  or (_16137_, _16136_, _16130_);
  or (_16138_, _16137_, _16129_);
  nor (_16139_, _16138_, _16128_);
  nand (_16140_, _16139_, _16110_);
  or (_16141_, _16140_, _16101_);
  and (_24414_, _16141_, _15988_);
  and (_16142_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _27355_);
  and (_16143_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_16144_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_16145_, _25987_, _16144_);
  not (_16146_, _16145_);
  not (_16147_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_16148_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_16149_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_16150_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_16151_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_16152_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_16153_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_16154_, _16153_, _16151_);
  and (_16155_, _16154_, _16152_);
  nor (_16156_, _16155_, _16151_);
  nor (_16157_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_16158_, _16157_, _16150_);
  not (_16159_, _16158_);
  nor (_16160_, _16159_, _16156_);
  nor (_16161_, _16160_, _16150_);
  not (_16162_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_16163_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_16164_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_16165_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_16166_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_16167_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_16168_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_16169_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_16170_, _16169_, _16168_);
  and (_16171_, _16170_, _16167_);
  and (_16172_, _16171_, _16166_);
  and (_16173_, _16172_, _16165_);
  and (_16174_, _16173_, _16164_);
  and (_16175_, _16174_, _16163_);
  and (_16176_, _16175_, _16162_);
  and (_16177_, _16176_, _16161_);
  and (_16178_, _16177_, _16149_);
  and (_16179_, _16178_, _16148_);
  and (_16180_, _16179_, _16147_);
  nor (_16181_, _16180_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_16182_, _16180_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_16183_, _16182_, _16181_);
  nor (_16184_, _16179_, _16147_);
  nor (_16185_, _16184_, _16180_);
  not (_16186_, _16185_);
  nor (_16187_, _16178_, _16148_);
  nor (_16188_, _16187_, _16179_);
  not (_16189_, _16188_);
  nor (_16190_, _16177_, _16149_);
  nor (_16191_, _16190_, _16178_);
  not (_16192_, _16191_);
  and (_16193_, _16161_, _16175_);
  nor (_16194_, _16193_, _16162_);
  nor (_16195_, _16194_, _16177_);
  not (_16196_, _16195_);
  and (_16197_, _16161_, _16173_);
  and (_16198_, _16197_, _16164_);
  nor (_16199_, _16198_, _16163_);
  or (_16200_, _16199_, _16193_);
  nor (_16201_, _16197_, _16164_);
  nor (_16202_, _16201_, _16198_);
  not (_16203_, _16202_);
  and (_16204_, _16161_, _16171_);
  nor (_16205_, _16204_, _16166_);
  and (_16206_, _16161_, _16172_);
  or (_16207_, _16206_, _16205_);
  and (_16208_, _16161_, _16170_);
  nor (_16209_, _16208_, _16167_);
  nor (_16210_, _16209_, _16204_);
  not (_16211_, _16210_);
  and (_16212_, _16161_, _16169_);
  nor (_16213_, _16212_, _16168_);
  nor (_16214_, _16213_, _16208_);
  not (_16215_, _16214_);
  not (_16216_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_16217_, _16161_, _16216_);
  nor (_16218_, _16161_, _16216_);
  nor (_16219_, _16218_, _16217_);
  not (_16220_, _16219_);
  and (_16221_, _15265_, _15243_);
  and (_16222_, _15221_, _15211_);
  and (_16223_, _15262_, _16222_);
  and (_16224_, _15262_, _15223_);
  or (_16225_, _16224_, _16223_);
  nor (_16226_, _16225_, _16221_);
  and (_16227_, _15289_, _15281_);
  and (_16228_, _15272_, _15235_);
  nor (_16229_, _16228_, _16227_);
  and (_16230_, _16229_, _16226_);
  nor (_16231_, _15293_, _15276_);
  not (_16232_, _26079_);
  and (_16233_, _15251_, _15221_);
  nor (_16234_, _16233_, _15269_);
  nor (_16235_, _16234_, _16232_);
  not (_16236_, _15272_);
  nor (_16237_, _15269_, _15292_);
  nor (_16238_, _16237_, _16236_);
  nor (_16239_, _16238_, _16235_);
  and (_16240_, _16239_, _16231_);
  and (_16241_, _16240_, _16230_);
  not (_16242_, _15262_);
  and (_16243_, _15215_, _15231_);
  nor (_16244_, _16233_, _16243_);
  nor (_16245_, _16244_, _16242_);
  not (_16246_, _16245_);
  and (_16247_, _15285_, _15272_);
  not (_16248_, _15208_);
  nor (_16249_, _15271_, _15269_);
  nor (_16250_, _16249_, _16248_);
  nor (_16251_, _16250_, _16247_);
  and (_16252_, _16251_, _16246_);
  and (_16253_, _16252_, _15268_);
  and (_16254_, _16253_, _16241_);
  not (_16255_, _15292_);
  nor (_16256_, _15208_, _26079_);
  nor (_16257_, _16256_, _16255_);
  not (_16258_, _16257_);
  and (_16259_, _15264_, _15215_);
  nor (_16260_, _16259_, _16222_);
  nor (_16261_, _15265_, _15216_);
  and (_16262_, _16261_, _16260_);
  nor (_16263_, _16262_, _16236_);
  not (_16264_, _15232_);
  nor (_16265_, _15272_, _15208_);
  nor (_16266_, _16265_, _16264_);
  nor (_16267_, _16266_, _16263_);
  and (_16268_, _16267_, _16258_);
  or (_16269_, _16233_, _16222_);
  not (_16270_, _16269_);
  nor (_16271_, _16259_, _15223_);
  and (_16272_, _16271_, _16270_);
  nor (_16273_, _16272_, _16248_);
  and (_16274_, _15225_, _16232_);
  and (_16275_, _15290_, _16274_);
  not (_16276_, _16275_);
  nor (_16277_, _15284_, _15227_);
  and (_16278_, _16277_, _16276_);
  not (_16279_, _16278_);
  nor (_16280_, _16279_, _16273_);
  and (_16281_, _15252_, _15211_);
  not (_16282_, _16281_);
  nor (_16283_, _15219_, _15208_);
  nor (_16284_, _16283_, _16282_);
  nor (_16285_, _15219_, _15207_);
  and (_16286_, _15265_, _26028_);
  nor (_16287_, _16286_, _15253_);
  nor (_16288_, _16287_, _16285_);
  nor (_16289_, _16288_, _16284_);
  and (_16290_, _16289_, _16280_);
  and (_16291_, _16290_, _16268_);
  nor (_16292_, _15283_, _15273_);
  nand (_16293_, _15224_, _15241_);
  and (_16294_, _15289_, _15223_);
  and (_16295_, _16281_, _15243_);
  nor (_16296_, _16295_, _16294_);
  and (_16297_, _16296_, _16293_);
  and (_16298_, _16297_, _16292_);
  not (_16299_, _16298_);
  nor (_16300_, _15289_, _16274_);
  not (_16301_, _15289_);
  nor (_16302_, _16222_, _15260_);
  nor (_16303_, _16302_, _16301_);
  nor (_16304_, _16303_, _15269_);
  nor (_16305_, _16304_, _16300_);
  nor (_16306_, _16305_, _16299_);
  and (_16307_, _16306_, _16291_);
  and (_16308_, _16307_, _16254_);
  nor (_16309_, _16154_, _16152_);
  nor (_16310_, _16309_, _16155_);
  not (_16311_, _16310_);
  nor (_16312_, _16311_, _16308_);
  not (_16313_, _16312_);
  and (_16314_, _15253_, _15243_);
  or (_16315_, _16223_, _16221_);
  or (_16316_, _16315_, _16314_);
  or (_16317_, _15263_, _15227_);
  or (_16318_, _16238_, _15233_);
  or (_16319_, _16318_, _16317_);
  or (_16320_, _16319_, _16316_);
  or (_16321_, _16320_, _16299_);
  nor (_16322_, _16321_, _16308_);
  not (_16323_, _16322_);
  nor (_16324_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_16325_, _16324_, _16152_);
  and (_16326_, _16325_, _16323_);
  and (_16327_, _16311_, _16308_);
  nor (_16328_, _16327_, _16312_);
  nand (_16329_, _16328_, _16326_);
  and (_16330_, _16329_, _16313_);
  not (_16331_, _16330_);
  and (_16332_, _16159_, _16156_);
  nor (_16333_, _16332_, _16160_);
  and (_16334_, _16333_, _16331_);
  and (_16335_, _16334_, _16220_);
  not (_16336_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_16337_, _16217_, _16336_);
  or (_16338_, _16337_, _16212_);
  and (_16339_, _16338_, _16335_);
  and (_16340_, _16339_, _16215_);
  and (_16341_, _16340_, _16211_);
  and (_16342_, _16341_, _16207_);
  nor (_16343_, _16206_, _16165_);
  or (_16344_, _16343_, _16197_);
  and (_16345_, _16344_, _16342_);
  and (_16346_, _16345_, _16203_);
  and (_16347_, _16346_, _16200_);
  and (_16348_, _16347_, _16196_);
  and (_16349_, _16348_, _16192_);
  and (_16350_, _16349_, _16189_);
  and (_16351_, _16350_, _16186_);
  or (_16352_, _16351_, _16183_);
  nand (_16353_, _16351_, _16183_);
  and (_16354_, _16353_, _16352_);
  or (_16355_, _16354_, _16146_);
  or (_16356_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_16357_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_16358_, _16357_, _16356_);
  and (_16359_, _16358_, _16355_);
  or (_24415_, _16359_, _16143_);
  nor (_16360_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_24416_, _16360_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_24417_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _27355_);
  nor (_16361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_16362_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_16363_, _16362_, _16361_);
  nor (_16364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_16365_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_16366_, _16365_, _16364_);
  and (_16367_, _16366_, _16363_);
  nor (_16368_, _16367_, rst);
  and (_16369_, \oc8051_top_1.oc8051_rom1.ea_int , _25984_);
  nand (_16370_, _16369_, _25987_);
  and (_16371_, _16370_, _24417_);
  or (_24418_, _16371_, _16368_);
  and (_16372_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_16373_, _16372_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_24419_, _16373_, _27355_);
  nor (_16374_, _15969_, _01726_);
  nor (_16375_, _16308_, _26000_);
  not (_16376_, _16375_);
  nor (_16377_, _16322_, _26016_);
  and (_16378_, _16308_, _26000_);
  nor (_16379_, _16378_, _16375_);
  nand (_16380_, _16379_, _16377_);
  and (_16381_, _16380_, _16376_);
  nor (_16382_, _16381_, _01726_);
  and (_16383_, _16382_, _25999_);
  nor (_16384_, _16382_, _25999_);
  nor (_16385_, _16384_, _16383_);
  nor (_16386_, _16385_, _16374_);
  and (_16387_, _26001_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_16388_, _16387_, _16374_);
  and (_16389_, _16388_, _16321_);
  or (_16390_, _16389_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_16391_, _16390_, _16386_);
  and (_24420_, _16391_, _27355_);
  and (_16392_, _26200_, _26023_);
  and (_16393_, _16392_, _26071_);
  and (_16394_, _26255_, _26142_);
  and (_16395_, _16394_, _26115_);
  and (_16396_, _25988_, _27355_);
  and (_16397_, _16396_, _26171_);
  and (_16398_, _16397_, _26227_);
  and (_16399_, _16398_, _16395_);
  and (_24423_, _16399_, _16393_);
  nor (_16400_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_16401_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_16402_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_24426_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _27355_);
  and (_16403_, _24426_, _16402_);
  or (_24424_, _16403_, _16401_);
  not (_16404_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_16405_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_16406_, _16405_, _16404_);
  and (_16407_, _16405_, _16404_);
  nor (_16408_, _16407_, _16406_);
  not (_16409_, _16408_);
  and (_16410_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_16411_, _16410_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_16412_, _16410_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_16413_, _16412_, _16411_);
  or (_16414_, _16413_, _16405_);
  and (_16415_, _16414_, _16409_);
  nor (_16416_, _16406_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_16417_, _16406_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_16418_, _16417_, _16416_);
  or (_16419_, _16411_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_24428_, _16419_, _27355_);
  and (_16420_, _24428_, _16418_);
  and (_24427_, _16420_, _16415_);
  not (_16421_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_16422_, _15969_, _16421_);
  and (_16423_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_16424_, _16422_);
  and (_16425_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_16426_, _16425_, _16423_);
  and (_24429_, _16426_, _27355_);
  and (_16427_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_16428_, _16422_, _26193_);
  or (_16429_, _16428_, _16427_);
  and (_24430_, _16429_, _27355_);
  and (_16430_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_16431_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16432_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _16431_);
  and (_16433_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_16434_, _16433_, _16430_);
  and (_24431_, _16434_, _27355_);
  and (_16435_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  or (_16436_, _16435_, _16432_);
  and (_24433_, _16436_, _27355_);
  or (_16437_, _16431_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_24434_, _16437_, _27355_);
  not (_16438_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_16439_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_16440_, _16439_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_16441_, _16431_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_16442_, _16441_, _27355_);
  and (_24435_, _16442_, _16440_);
  or (_16443_, _16431_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_24436_, _16443_, _27355_);
  nor (_16444_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_16445_, _16444_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16446_, _16445_, _27355_);
  and (_16447_, _24426_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_24437_, _16447_, _16446_);
  and (_16448_, _16421_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_16449_, _16448_, _16445_);
  and (_24438_, _16449_, _27355_);
  not (_16450_, _16445_);
  or (_16451_, _16450_, _26678_);
  or (_16452_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_16453_, _16452_, _27355_);
  and (_24439_, _16453_, _16451_);
  and (_16454_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_16455_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_16456_, pc_log_change, _16455_);
  or (_16457_, _16456_, _16454_);
  and (_24470_, _16457_, _27355_);
  and (_16458_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_16459_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_16460_, pc_log_change, _16459_);
  or (_16461_, _16460_, _16458_);
  and (_24472_, _16461_, _27355_);
  and (_16462_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_16463_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_16464_, pc_log_change, _16463_);
  or (_16465_, _16464_, _16462_);
  and (_24473_, _16465_, _27355_);
  and (_16466_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_16467_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_16468_, pc_log_change, _16467_);
  or (_16469_, _16468_, _16466_);
  and (_24474_, _16469_, _27355_);
  and (_16470_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_16471_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_16472_, pc_log_change, _16471_);
  or (_16473_, _16472_, _16470_);
  and (_24475_, _16473_, _27355_);
  and (_16474_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_16475_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_16476_, pc_log_change, _16475_);
  or (_16477_, _16476_, _16474_);
  and (_24476_, _16477_, _27355_);
  and (_16478_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_16479_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_16480_, pc_log_change, _16479_);
  or (_16481_, _16480_, _16478_);
  and (_24477_, _16481_, _27355_);
  and (_16482_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_16483_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_16484_, pc_log_change, _16483_);
  or (_16485_, _16484_, _16482_);
  and (_24478_, _16485_, _27355_);
  and (_16486_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_16487_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_16488_, pc_log_change, _16487_);
  or (_16489_, _16488_, _16486_);
  and (_24479_, _16489_, _27355_);
  and (_16490_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_16491_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_16492_, pc_log_change, _16491_);
  or (_16493_, _16492_, _16490_);
  and (_24480_, _16493_, _27355_);
  and (_16494_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_16495_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_16496_, pc_log_change, _16495_);
  or (_16497_, _16496_, _16494_);
  and (_24481_, _16497_, _27355_);
  and (_16498_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_16499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_16500_, pc_log_change, _16499_);
  or (_16501_, _16500_, _16498_);
  and (_24483_, _16501_, _27355_);
  and (_16502_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_16503_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_16504_, pc_log_change, _16503_);
  or (_16505_, _16504_, _16502_);
  and (_24484_, _16505_, _27355_);
  and (_16506_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_16507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_16508_, pc_log_change, _16507_);
  or (_16509_, _16508_, _16506_);
  and (_24485_, _16509_, _27355_);
  and (_16510_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_16511_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_16512_, pc_log_change, _16511_);
  or (_16513_, _16512_, _16510_);
  and (_24486_, _16513_, _27355_);
  and (_16514_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_16515_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_16516_, pc_log_change, _16515_);
  or (_16517_, _16516_, _16514_);
  and (_24490_, _16517_, _27355_);
  and (_16518_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_16519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_16520_, pc_log_change, _16519_);
  or (_16521_, _16520_, _16518_);
  and (_24491_, _16521_, _27355_);
  and (_16522_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_16523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_16524_, pc_log_change, _16523_);
  or (_16525_, _16524_, _16522_);
  and (_24492_, _16525_, _27355_);
  and (_16526_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_16527_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_16528_, pc_log_change, _16527_);
  or (_16529_, _16528_, _16526_);
  and (_24493_, _16529_, _27355_);
  or (_16530_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand (_16531_, pc_log_change, _16471_);
  and (_16532_, _16531_, _27355_);
  and (_24494_, _16532_, _16530_);
  or (_16533_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand (_16534_, pc_log_change, _16475_);
  and (_16535_, _16534_, _27355_);
  and (_24495_, _16535_, _16533_);
  or (_16536_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand (_16537_, pc_log_change, _16479_);
  and (_16538_, _16537_, _27355_);
  and (_24497_, _16538_, _16536_);
  and (_16539_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_16540_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_16541_, pc_log_change, _16540_);
  or (_16542_, _16541_, _16539_);
  and (_24498_, _16542_, _27355_);
  or (_16543_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand (_16544_, pc_log_change, _16487_);
  and (_16545_, _16544_, _27355_);
  and (_24499_, _16545_, _16543_);
  and (_16546_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not (_16547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_16548_, pc_log_change, _16547_);
  or (_16549_, _16548_, _16546_);
  and (_24500_, _16549_, _27355_);
  and (_16550_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not (_16551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_16552_, pc_log_change, _16551_);
  or (_16553_, _16552_, _16550_);
  and (_24501_, _16553_, _27355_);
  or (_16554_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nand (_16555_, pc_log_change, _16499_);
  and (_16556_, _16555_, _27355_);
  and (_24502_, _16556_, _16554_);
  and (_16557_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  not (_16558_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_16559_, pc_log_change, _16558_);
  or (_16560_, _16559_, _16557_);
  and (_24503_, _16560_, _27355_);
  or (_16561_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nand (_16562_, pc_log_change, _16507_);
  and (_16563_, _16562_, _27355_);
  and (_24504_, _16563_, _16561_);
  or (_16564_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand (_16565_, pc_log_change, _16511_);
  and (_16566_, _16565_, _27355_);
  and (_24505_, _16566_, _16564_);
  and (_24692_, _26033_, _27355_);
  and (_24693_, _26153_, _27355_);
  and (_24695_, _26125_, _27355_);
  nor (_24696_, _01632_, rst);
  nor (_16567_, _16422_, _26008_);
  and (_16568_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_16569_, _16568_, _16422_);
  or (_16570_, _16569_, _16567_);
  and (_24697_, _16570_, _27355_);
  nor (_16571_, _16422_, _26127_);
  and (_16572_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_16573_, _16572_, _16422_);
  or (_16574_, _16573_, _16571_);
  and (_24698_, _16574_, _27355_);
  nor (_16575_, _16422_, _26105_);
  and (_16576_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_16577_, _16576_, _16575_);
  and (_24699_, _16577_, _27355_);
  nor (_16578_, _16422_, _26051_);
  and (_16579_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_16580_, _16579_, _16578_);
  and (_24700_, _16580_, _27355_);
  nor (_16581_, _16422_, _26157_);
  and (_16582_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_16583_, _16582_, _16581_);
  and (_24701_, _16583_, _27355_);
  nor (_16584_, _16422_, _26218_);
  and (_16585_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_16586_, _16585_, _16422_);
  or (_16587_, _16586_, _16584_);
  and (_24702_, _16587_, _27355_);
  nor (_16588_, _16422_, _26251_);
  and (_16589_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_16590_, _16589_, _16588_);
  and (_24703_, _16590_, _27355_);
  nor (_16591_, _16422_, _26190_);
  and (_16592_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_16593_, _16592_, _16591_);
  and (_24704_, _16593_, _27355_);
  and (_16594_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nor (_16595_, _16422_, _01841_);
  or (_16596_, _16595_, _16594_);
  and (_24706_, _16596_, _27355_);
  and (_16597_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nor (_16598_, _16422_, _01935_);
  or (_16599_, _16598_, _16597_);
  and (_24707_, _16599_, _27355_);
  and (_16600_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nor (_16601_, _16422_, _02112_);
  or (_16602_, _16601_, _16600_);
  and (_24708_, _16602_, _27355_);
  and (_16603_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nor (_16604_, _16422_, _01794_);
  or (_16605_, _16604_, _16603_);
  and (_24709_, _16605_, _27355_);
  and (_16606_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nor (_16607_, _16422_, _01892_);
  or (_16608_, _16607_, _16606_);
  and (_24710_, _16608_, _27355_);
  and (_16609_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nor (_16610_, _16422_, _01971_);
  or (_16611_, _16610_, _16609_);
  and (_24711_, _16611_, _27355_);
  and (_16612_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nor (_16613_, _16422_, _02035_);
  or (_16614_, _16613_, _16612_);
  and (_24712_, _16614_, _27355_);
  and (_16615_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nor (_16616_, _16422_, _01735_);
  or (_16617_, _16616_, _16615_);
  and (_24713_, _16617_, _27355_);
  and (_16618_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_16619_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_16620_, _16619_, _16618_);
  and (_24714_, _16620_, _27355_);
  and (_16621_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_16622_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_16623_, _16622_, _16621_);
  and (_24715_, _16623_, _27355_);
  and (_16624_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_16625_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_16626_, _16625_, _16624_);
  and (_24717_, _16626_, _27355_);
  and (_16627_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_16628_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_16629_, _16628_, _16627_);
  and (_24718_, _16629_, _27355_);
  and (_16630_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_16631_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_16632_, _16631_, _16630_);
  and (_24719_, _16632_, _27355_);
  and (_16633_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_16634_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_16635_, _16634_, _16633_);
  and (_24720_, _16635_, _27355_);
  and (_16636_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_16637_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_16638_, _16637_, _16636_);
  and (_24721_, _16638_, _27355_);
  and (_16639_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_16640_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_16641_, _16640_, _16639_);
  and (_24722_, _16641_, _27355_);
  and (_16642_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_16643_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_16644_, _16643_, _16642_);
  and (_24723_, _16644_, _27355_);
  and (_16645_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_16646_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_16647_, _16646_, _16645_);
  and (_24724_, _16647_, _27355_);
  and (_16648_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_16649_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_16650_, _16649_, _16648_);
  and (_24725_, _16650_, _27355_);
  and (_16651_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_16652_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_16653_, _16652_, _16651_);
  and (_24726_, _16653_, _27355_);
  and (_16654_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_16655_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_16656_, _16655_, _16654_);
  and (_24728_, _16656_, _27355_);
  and (_16657_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_16658_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_16659_, _16658_, _16657_);
  and (_24729_, _16659_, _27355_);
  and (_16660_, _16422_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_16661_, _16424_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_16662_, _16661_, _16660_);
  and (_24730_, _16662_, _27355_);
  and (_24731_, _01830_, _27355_);
  and (_24732_, _01926_, _27355_);
  and (_24733_, _02104_, _27355_);
  and (_24735_, _01784_, _27355_);
  and (_24736_, _01880_, _27355_);
  and (_24737_, _02000_, _27355_);
  and (_24738_, _02029_, _27355_);
  and (_24755_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _27355_);
  and (_24756_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _27355_);
  and (_24757_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _27355_);
  and (_24758_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _27355_);
  and (_24759_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _27355_);
  and (_24760_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _27355_);
  and (_24761_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _27355_);
  not (_16663_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_16664_, _15966_, _16663_);
  or (_16665_, _16132_, _16096_);
  and (_16666_, _16665_, _25563_);
  or (_16667_, _16045_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_16668_, _16046_);
  and (_16669_, _26311_, _25983_);
  and (_16670_, _16669_, _26286_);
  nor (_16671_, _16094_, _16670_);
  not (_16672_, _16670_);
  nor (_16673_, _16134_, _15865_);
  and (_16674_, _16673_, _15994_);
  and (_16675_, _16674_, _16672_);
  and (_16676_, _16098_, _16675_);
  nor (_16677_, _16676_, _16671_);
  and (_16678_, _16677_, _16668_);
  and (_16679_, _16678_, _16667_);
  and (_16680_, _16134_, _16043_);
  not (_16681_, _16094_);
  and (_16682_, _16676_, _16681_);
  and (_16683_, _16682_, _01848_);
  or (_16684_, _16683_, _16680_);
  or (_16685_, _16684_, _16679_);
  or (_16686_, _16685_, _16666_);
  and (_16687_, _16686_, _16110_);
  or (_16688_, _16687_, _16664_);
  and (_24762_, _16688_, _27355_);
  not (_16689_, _15965_);
  and (_16690_, _16689_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_16691_, _16665_, _25639_);
  or (_16692_, _16048_, _16046_);
  not (_16693_, _16049_);
  and (_16694_, _16677_, _16693_);
  and (_16695_, _16694_, _16692_);
  and (_16696_, _16682_, _01948_);
  and (_16697_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_16698_, _16134_, _16037_);
  or (_16699_, _16698_, _16697_);
  or (_16700_, _16699_, _16696_);
  or (_16701_, _16700_, _16695_);
  or (_16702_, _16701_, _16691_);
  and (_16703_, _16702_, _15965_);
  or (_16704_, _16703_, _16690_);
  and (_24763_, _16704_, _27355_);
  not (_16705_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_16706_, _15969_, _16705_);
  and (_16707_, _15969_, _16705_);
  nor (_16708_, _16707_, _16706_);
  and (_16709_, _16708_, _16689_);
  and (_16710_, _16665_, _25705_);
  or (_16711_, _16053_, _16050_);
  not (_16712_, _16054_);
  and (_16713_, _16677_, _16712_);
  and (_16714_, _16713_, _16711_);
  and (_16715_, _16682_, _02125_);
  and (_16716_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_16717_, _16134_, _16032_);
  or (_16718_, _16717_, _16716_);
  or (_16719_, _16718_, _16715_);
  or (_16720_, _16719_, _16714_);
  or (_16721_, _16720_, _16710_);
  and (_16722_, _16721_, _15965_);
  or (_16723_, _16722_, _16709_);
  and (_24765_, _16723_, _27355_);
  and (_16724_, _16706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_16725_, _16706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_16726_, _16725_, _16724_);
  or (_16727_, _16726_, _15965_);
  and (_16728_, _16727_, _27355_);
  and (_16729_, _16665_, _25770_);
  and (_16730_, _15995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not (_16731_, _15806_);
  and (_16732_, _15997_, _16731_);
  and (_16733_, _16127_, _01807_);
  or (_16734_, _16733_, _16732_);
  or (_16735_, _16734_, _16730_);
  or (_16736_, _16029_, _16030_);
  and (_16737_, _16736_, _16055_);
  nor (_16738_, _16736_, _16055_);
  or (_16739_, _16738_, _16737_);
  and (_16740_, _16739_, _16100_);
  or (_16741_, _16740_, _16735_);
  nor (_16742_, _16741_, _16729_);
  nand (_16743_, _16742_, _16110_);
  and (_24766_, _16743_, _16728_);
  and (_16744_, _15972_, _15970_);
  nor (_16745_, _16724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_16746_, _16745_, _16744_);
  or (_16747_, _16746_, _15965_);
  and (_16748_, _16747_, _27355_);
  and (_16749_, _16665_, _25830_);
  or (_16750_, _16059_, _16057_);
  and (_16751_, _16677_, _16060_);
  and (_16752_, _16751_, _16750_);
  and (_16753_, _16682_, _01903_);
  and (_16754_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  not (_16755_, _15823_);
  and (_16756_, _16134_, _16755_);
  or (_16757_, _16756_, _16754_);
  or (_16758_, _16757_, _16753_);
  nor (_16759_, _16758_, _16752_);
  nand (_16760_, _16759_, _15965_);
  or (_16761_, _16760_, _16749_);
  and (_24767_, _16761_, _16748_);
  nor (_16762_, _16744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_16763_, _16762_, _15974_);
  nor (_16764_, _16763_, _15965_);
  and (_16765_, _16665_, _25898_);
  not (_16766_, _16061_);
  or (_16767_, _16021_, _16020_);
  nand (_16768_, _16767_, _16766_);
  or (_16769_, _16767_, _16766_);
  and (_16770_, _16769_, _16677_);
  and (_16771_, _16770_, _16768_);
  and (_16772_, _16682_, _01981_);
  and (_16773_, _15865_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_16774_, _15840_);
  and (_16775_, _16134_, _16774_);
  or (_16776_, _16775_, _16773_);
  or (_16777_, _16776_, _16772_);
  or (_16778_, _16777_, _16771_);
  or (_16779_, _16778_, _16765_);
  and (_16780_, _16779_, _15965_);
  or (_16781_, _16780_, _16764_);
  and (_24768_, _16781_, _27355_);
  nor (_16782_, _15974_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_16783_, _16782_, _15975_);
  or (_16784_, _16783_, _15965_);
  and (_16785_, _16784_, _27355_);
  or (_16786_, _16063_, _16016_);
  and (_16787_, _16786_, _16064_);
  and (_16788_, _16787_, _16100_);
  and (_16789_, _16665_, _25964_);
  and (_16790_, _15995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_16791_, _15857_);
  and (_16792_, _15997_, _16791_);
  and (_16793_, _16127_, _02048_);
  or (_16794_, _16793_, _16792_);
  or (_16795_, _16794_, _16790_);
  or (_16796_, _16795_, _16789_);
  nor (_16797_, _16796_, _16788_);
  nand (_16798_, _16797_, _16110_);
  and (_24769_, _16798_, _16785_);
  nor (_16799_, _15975_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_16800_, _16799_, _15976_);
  or (_16801_, _16800_, _15965_);
  and (_16802_, _16801_, _27355_);
  and (_16803_, _16665_, _25441_);
  and (_16804_, _15995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_16805_, _15738_);
  and (_16806_, _15997_, _16805_);
  and (_16807_, _16127_, _01744_);
  or (_16808_, _16807_, _16806_);
  or (_16809_, _16808_, _16804_);
  nand (_16810_, _16065_, _16009_);
  and (_16811_, _16100_, _16066_);
  and (_16812_, _16811_, _16810_);
  or (_16813_, _16812_, _16809_);
  nor (_16814_, _16813_, _16803_);
  nand (_16815_, _16814_, _16110_);
  and (_24770_, _16815_, _16802_);
  nor (_16816_, _15976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_16817_, _16816_, _15977_);
  or (_16818_, _16817_, _15965_);
  and (_16819_, _16818_, _27355_);
  nor (_16820_, _16067_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_16821_, _16067_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_16822_, _16821_, _16820_);
  nor (_16823_, _16822_, _16004_);
  and (_16824_, _16822_, _16004_);
  or (_16825_, _16824_, _16823_);
  and (_16826_, _16825_, _16677_);
  nor (_16827_, _15866_, _25562_);
  and (_16828_, _16096_, _26713_);
  and (_16829_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_16830_, _16134_, _01848_);
  or (_16831_, _16830_, _16829_);
  and (_16832_, _16682_, _26232_);
  nor (_16833_, _16832_, _16831_);
  nand (_16834_, _16833_, _15965_);
  or (_16835_, _16834_, _16828_);
  or (_16836_, _16835_, _16827_);
  or (_16837_, _16836_, _16826_);
  and (_24771_, _16837_, _16819_);
  nor (_16838_, _15977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_16839_, _16838_, _15978_);
  or (_16840_, _16839_, _15965_);
  and (_16841_, _16840_, _27355_);
  nor (_16842_, _16068_, _16076_);
  and (_16843_, _16077_, _16076_);
  nor (_16844_, _16843_, _16842_);
  nand (_16845_, _16844_, _24188_);
  or (_16846_, _16844_, _24188_);
  and (_16847_, _16846_, _16845_);
  and (_16848_, _16847_, _16100_);
  and (_16849_, _16127_, _26259_);
  and (_16850_, _15995_, _25639_);
  not (_16851_, _16096_);
  nor (_16852_, _16851_, _26745_);
  and (_16853_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_16854_, _16134_, _01948_);
  or (_16855_, _16854_, _16853_);
  or (_16856_, _16855_, _16852_);
  or (_16857_, _16856_, _16850_);
  nor (_16858_, _16857_, _16849_);
  nand (_16859_, _16858_, _16110_);
  or (_16860_, _16859_, _16848_);
  and (_24772_, _16860_, _16841_);
  nor (_16861_, _15978_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_16862_, _16861_, _15979_);
  or (_16863_, _16862_, _15965_);
  and (_16864_, _16863_, _27355_);
  and (_16865_, _16842_, _24188_);
  and (_16866_, _16078_, _16076_);
  nor (_16867_, _16866_, _16865_);
  nand (_16868_, _16867_, _24204_);
  or (_16869_, _16867_, _24204_);
  and (_16870_, _16869_, _16677_);
  and (_16871_, _16870_, _16868_);
  nor (_16872_, _15866_, _25704_);
  nor (_16873_, _16851_, _26775_);
  and (_16874_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_16875_, _16134_, _02125_);
  or (_16876_, _16875_, _16874_);
  and (_16877_, _16127_, _26204_);
  or (_16878_, _16877_, _16876_);
  nor (_16879_, _16878_, _16873_);
  nand (_16880_, _16879_, _15965_);
  or (_16881_, _16880_, _16872_);
  or (_16882_, _16881_, _16871_);
  and (_24773_, _16882_, _16864_);
  nor (_16883_, _15979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_16884_, _15979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_16885_, _16884_, _16883_);
  or (_16886_, _16885_, _15965_);
  and (_16887_, _16886_, _27355_);
  nand (_16888_, _16079_, _16076_);
  or (_16889_, _16070_, _16076_);
  nand (_16890_, _16889_, _16888_);
  nand (_16891_, _16890_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_16892_, _16890_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_16893_, _16892_, _16677_);
  and (_16894_, _16893_, _16891_);
  nor (_16895_, _15866_, _25769_);
  nor (_16896_, _16851_, _26808_);
  and (_16897_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_16898_, _16134_, _01807_);
  or (_16899_, _16898_, _16897_);
  nor (_16900_, _16119_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_16901_, _16900_, _16120_);
  and (_16902_, _16901_, _16682_);
  or (_16903_, _16902_, _16899_);
  nor (_16904_, _16903_, _16896_);
  nand (_16905_, _16904_, _15965_);
  or (_16906_, _16905_, _16895_);
  or (_16907_, _16906_, _16894_);
  and (_24774_, _16907_, _16887_);
  nor (_16908_, _16884_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_16909_, _16908_, _15981_);
  or (_16910_, _16909_, _15965_);
  and (_16911_, _16910_, _27355_);
  nor (_16912_, _16071_, _16076_);
  and (_16913_, _16080_, _16076_);
  nor (_16914_, _16913_, _16912_);
  nand (_16915_, _16914_, _23940_);
  or (_16916_, _16914_, _23940_);
  and (_16917_, _16916_, _16915_);
  and (_16918_, _16917_, _16100_);
  nor (_16919_, _16120_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_16920_, _16919_, _16121_);
  and (_16921_, _16920_, _16127_);
  and (_16922_, _15995_, _25830_);
  and (_16923_, _16096_, _26837_);
  and (_16924_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_16925_, _16134_, _01903_);
  or (_16926_, _16925_, _16924_);
  or (_16927_, _16926_, _16923_);
  or (_16928_, _16927_, _16922_);
  nor (_16929_, _16928_, _16921_);
  nand (_16930_, _16929_, _16110_);
  or (_16931_, _16930_, _16918_);
  and (_24776_, _16931_, _16911_);
  not (_16932_, _16110_);
  or (_16933_, _16072_, _16076_);
  nand (_16934_, _16913_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_16935_, _16934_, _16933_);
  nor (_16936_, _16935_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_16937_, _16935_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_16938_, _16937_, _16936_);
  and (_16939_, _16938_, _16677_);
  and (_16940_, _15865_, _25898_);
  and (_16941_, _16096_, _26867_);
  and (_16942_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_16943_, _16134_, _01981_);
  or (_16944_, _16943_, _16942_);
  nor (_16945_, _16121_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_16946_, _16945_, _16122_);
  and (_16947_, _16946_, _16682_);
  or (_16948_, _16947_, _16944_);
  or (_16949_, _16948_, _16941_);
  or (_16950_, _16949_, _16940_);
  or (_16951_, _16950_, _16939_);
  or (_16952_, _16951_, _16932_);
  nor (_16953_, _15981_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_16954_, _16953_, _15982_);
  or (_16955_, _16954_, _16110_);
  and (_16956_, _16955_, _27355_);
  and (_24777_, _16956_, _16952_);
  or (_16957_, _16082_, _16004_);
  or (_16958_, _16073_, _16076_);
  and (_16959_, _16958_, _16957_);
  nor (_16960_, _16959_, _24129_);
  and (_16961_, _16959_, _24129_);
  or (_16962_, _16961_, _16960_);
  and (_16963_, _16962_, _16677_);
  nor (_16964_, _15866_, _25963_);
  nor (_16965_, _16851_, _26898_);
  and (_16966_, _16132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_16967_, _16134_, _02048_);
  or (_16968_, _16967_, _16966_);
  or (_16969_, _16122_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_16970_, _16969_, _16123_);
  and (_16971_, _16970_, _16682_);
  or (_16972_, _16971_, _16968_);
  or (_16973_, _16972_, _16965_);
  or (_16974_, _16973_, _16964_);
  or (_16975_, _16974_, _16963_);
  or (_16976_, _16975_, _16932_);
  nor (_16977_, _15982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_16978_, _16977_, _15983_);
  or (_16979_, _16978_, _16110_);
  and (_16980_, _16979_, _27355_);
  and (_24778_, _16980_, _16976_);
  and (_16981_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_16982_, _16325_, _16323_);
  nor (_16983_, _16982_, _16326_);
  or (_16984_, _16983_, _16146_);
  or (_16985_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_16986_, _16985_, _16357_);
  and (_16987_, _16986_, _16984_);
  or (_24779_, _16987_, _16981_);
  or (_16988_, _16328_, _16326_);
  and (_16989_, _16988_, _16329_);
  or (_16990_, _16989_, _16146_);
  or (_16991_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_16992_, _16991_, _16357_);
  and (_16993_, _16992_, _16990_);
  and (_16994_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_24780_, _16994_, _16993_);
  nor (_16995_, _16333_, _16331_);
  nor (_16996_, _16995_, _16334_);
  or (_16997_, _16996_, _16146_);
  or (_16998_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_16999_, _16998_, _16357_);
  and (_17000_, _16999_, _16997_);
  and (_17001_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_24781_, _17001_, _17000_);
  nor (_17002_, _16334_, _16220_);
  nor (_17003_, _17002_, _16335_);
  or (_17004_, _17003_, _16146_);
  or (_17005_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_17006_, _17005_, _16357_);
  and (_17007_, _17006_, _17004_);
  and (_17008_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_24782_, _17008_, _17007_);
  and (_17009_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_17010_, _16338_, _16335_);
  nor (_17011_, _17010_, _16339_);
  or (_17012_, _17011_, _16146_);
  or (_17013_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_17014_, _17013_, _16357_);
  and (_17015_, _17014_, _17012_);
  or (_24783_, _17015_, _17009_);
  and (_17016_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_17017_, _16339_, _16215_);
  nor (_17018_, _17017_, _16340_);
  or (_17019_, _17018_, _16146_);
  or (_17020_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_17021_, _17020_, _16357_);
  and (_17022_, _17021_, _17019_);
  or (_24784_, _17022_, _17016_);
  and (_17023_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_17024_, _16340_, _16211_);
  nor (_17025_, _17024_, _16341_);
  or (_17026_, _17025_, _16146_);
  or (_17027_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_17028_, _17027_, _16357_);
  and (_17029_, _17028_, _17026_);
  or (_24785_, _17029_, _17023_);
  or (_17030_, _16341_, _16207_);
  nor (_17031_, _16342_, _16146_);
  and (_17032_, _17031_, _17030_);
  nor (_17033_, _16145_, _24160_);
  or (_17034_, _17033_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_17035_, _17034_, _17032_);
  or (_17036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _25984_);
  and (_17037_, _17036_, _27355_);
  and (_24787_, _17037_, _17035_);
  nor (_17038_, _16344_, _16342_);
  nor (_17039_, _17038_, _16345_);
  or (_17040_, _17039_, _16146_);
  or (_17041_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_17042_, _17041_, _16357_);
  and (_17043_, _17042_, _17040_);
  and (_17044_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_24788_, _17044_, _17043_);
  nor (_17045_, _16345_, _16203_);
  nor (_17046_, _17045_, _16346_);
  or (_17047_, _17046_, _16146_);
  or (_17048_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_17049_, _17048_, _16357_);
  and (_17050_, _17049_, _17047_);
  and (_17051_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_24789_, _17051_, _17050_);
  nor (_17052_, _16346_, _16200_);
  nor (_17053_, _17052_, _16347_);
  or (_17054_, _17053_, _16146_);
  or (_17055_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_17056_, _17055_, _16357_);
  and (_17057_, _17056_, _17054_);
  and (_17058_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_24790_, _17058_, _17057_);
  nor (_17059_, _16347_, _16196_);
  nor (_17060_, _17059_, _16348_);
  or (_17061_, _17060_, _16146_);
  or (_17062_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_17063_, _17062_, _16357_);
  and (_17064_, _17063_, _17061_);
  and (_17065_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_24791_, _17065_, _17064_);
  nor (_17066_, _16348_, _16192_);
  nor (_17067_, _17066_, _16349_);
  or (_17068_, _17067_, _16146_);
  or (_17069_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_17070_, _17069_, _16357_);
  and (_17071_, _17070_, _17068_);
  and (_17072_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_24792_, _17072_, _17071_);
  nor (_17073_, _16349_, _16189_);
  nor (_17074_, _17073_, _16350_);
  or (_17075_, _17074_, _16146_);
  or (_17076_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_17077_, _17076_, _16357_);
  and (_17078_, _17077_, _17075_);
  and (_17079_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_24793_, _17079_, _17078_);
  and (_17080_, _16142_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_17081_, _16350_, _16186_);
  nor (_17082_, _17081_, _16351_);
  or (_17083_, _17082_, _16146_);
  or (_17084_, _16145_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_17085_, _17084_, _16357_);
  and (_17086_, _17085_, _17083_);
  or (_24794_, _17086_, _17080_);
  and (_17087_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_17088_, _17087_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_24795_, _17088_, _27355_);
  and (_17089_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_17090_, _17089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_24796_, _17090_, _27355_);
  and (_17091_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_17092_, _17091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_24798_, _17092_, _27355_);
  and (_17093_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_17094_, _17093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_24799_, _17094_, _27355_);
  and (_17095_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_17096_, _17095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_24800_, _17096_, _27355_);
  and (_17097_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_17098_, _17097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_24801_, _17098_, _27355_);
  and (_17099_, _16367_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_17100_, _17099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_24802_, _17100_, _27355_);
  nor (_17101_, _16322_, _01726_);
  nand (_17102_, _17101_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_17103_, _17101_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_17104_, _17103_, _16357_);
  and (_24803_, _17104_, _17102_);
  or (_17105_, _16379_, _16377_);
  and (_17106_, _17105_, _16380_);
  or (_17107_, _17106_, _01726_);
  or (_17108_, _25987_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_17109_, _17108_, _16357_);
  and (_24804_, _17109_, _17107_);
  and (_17110_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_17111_, _16568_, _24426_);
  or (_24821_, _17111_, _17110_);
  and (_17112_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_17113_, _16572_, _24426_);
  or (_24822_, _17113_, _17112_);
  and (_17114_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_17115_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_17116_, _17115_, _24426_);
  or (_24823_, _17116_, _17114_);
  and (_17117_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_17118_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_17119_, _17118_, _24426_);
  or (_24824_, _17119_, _17117_);
  and (_17120_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_17121_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_17122_, _17121_, _24426_);
  or (_24825_, _17122_, _17120_);
  and (_17123_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_17124_, _16585_, _24426_);
  or (_24826_, _17124_, _17123_);
  and (_17125_, _16400_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_17126_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_17127_, _17126_, _24426_);
  or (_24827_, _17127_, _17125_);
  and (_24828_, _16408_, _27355_);
  nor (_24829_, _16418_, rst);
  and (_24831_, _16414_, _27355_);
  or (_17128_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand (_17129_, _16422_, _26008_);
  and (_17130_, _17129_, _27355_);
  and (_24832_, _17130_, _17128_);
  or (_17131_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nand (_17132_, _16422_, _26127_);
  and (_17133_, _17132_, _27355_);
  and (_24833_, _17133_, _17131_);
  or (_17134_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_17135_, _16422_, _26105_);
  and (_17136_, _17135_, _27355_);
  and (_24834_, _17136_, _17134_);
  or (_17137_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_17138_, _16422_, _26051_);
  and (_17139_, _17138_, _27355_);
  and (_24835_, _17139_, _17137_);
  or (_17140_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand (_17141_, _16422_, _26157_);
  and (_17142_, _17141_, _27355_);
  and (_24836_, _17142_, _17140_);
  or (_17143_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_17144_, _16422_, _26218_);
  and (_17145_, _17144_, _27355_);
  and (_24837_, _17145_, _17143_);
  or (_17146_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_17147_, _16422_, _26251_);
  and (_17148_, _17147_, _27355_);
  and (_24838_, _17148_, _17146_);
  or (_17149_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_17150_, _16422_, _26190_);
  and (_17151_, _17150_, _27355_);
  and (_24839_, _17151_, _17149_);
  and (_17152_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_17153_, _16422_, _25998_);
  or (_17154_, _17153_, _17152_);
  and (_24840_, _17154_, _27355_);
  and (_17155_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_17156_, _16422_, _26135_);
  or (_17157_, _17156_, _17155_);
  and (_24842_, _17157_, _27355_);
  and (_17158_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_17159_, _16422_, _26093_);
  or (_17160_, _17159_, _17158_);
  and (_24843_, _17160_, _27355_);
  and (_17161_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_17162_, _16422_, _26061_);
  or (_17163_, _17162_, _17161_);
  and (_24844_, _17163_, _27355_);
  and (_17164_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_17165_, _16422_, _26163_);
  or (_17166_, _17165_, _17164_);
  and (_24845_, _17166_, _27355_);
  and (_17167_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_17168_, _16422_, _26214_);
  or (_17169_, _17168_, _17167_);
  and (_24846_, _17169_, _27355_);
  and (_17170_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_17171_, _16422_, _26242_);
  or (_17172_, _17171_, _17170_);
  and (_24847_, _17172_, _27355_);
  and (_17173_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_17174_, _16422_, _26195_);
  or (_17175_, _17174_, _17173_);
  and (_24848_, _17175_, _27355_);
  and (_17176_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_17177_, _16422_, _26015_);
  or (_17178_, _17177_, _17176_);
  and (_24849_, _17178_, _27355_);
  and (_17179_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor (_17180_, _16422_, _26132_);
  or (_17181_, _17180_, _17179_);
  and (_24850_, _17181_, _27355_);
  and (_17182_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_17183_, _16422_, _26097_);
  or (_17184_, _17183_, _17182_);
  and (_24851_, _17184_, _27355_);
  and (_17185_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_17186_, _16422_, _26043_);
  or (_17187_, _17186_, _17185_);
  and (_24853_, _17187_, _27355_);
  and (_17188_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_17189_, _16422_, _26167_);
  or (_17190_, _17189_, _17188_);
  and (_24854_, _17190_, _27355_);
  and (_17191_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_17192_, _16422_, _26222_);
  or (_17193_, _17192_, _17191_);
  and (_24855_, _17193_, _27355_);
  and (_17194_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_17195_, _16422_, _26247_);
  or (_17196_, _17195_, _17194_);
  and (_24856_, _17196_, _27355_);
  and (_17197_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_17198_, _16422_, _26186_);
  or (_17199_, _17198_, _17197_);
  and (_24857_, _17199_, _27355_);
  and (_17200_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor (_17201_, _16422_, _25994_);
  or (_17202_, _17201_, _17200_);
  and (_24858_, _17202_, _27355_);
  and (_17203_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor (_17204_, _16422_, _26129_);
  or (_17205_, _17204_, _17203_);
  and (_24859_, _17205_, _27355_);
  and (_17206_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor (_17207_, _16422_, _26111_);
  or (_17208_, _17207_, _17206_);
  and (_24860_, _17208_, _27355_);
  and (_17209_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor (_17210_, _16422_, _26057_);
  or (_17211_, _17210_, _17209_);
  and (_24861_, _17211_, _27355_);
  and (_17212_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor (_17213_, _16422_, _26159_);
  or (_17214_, _17213_, _17212_);
  and (_24862_, _17214_, _27355_);
  and (_17215_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_17216_, _16422_, _26212_);
  or (_17217_, _17216_, _17215_);
  and (_24864_, _17217_, _27355_);
  and (_17218_, _16422_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor (_17219_, _16422_, _26245_);
  or (_17220_, _17219_, _17218_);
  and (_24865_, _17220_, _27355_);
  and (_17221_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_17222_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_17223_, _17222_, _17221_);
  and (_24866_, _17223_, _27355_);
  and (_17224_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_17225_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_17226_, _17225_, _17224_);
  and (_24867_, _17226_, _27355_);
  and (_17227_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_17228_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_17229_, _17228_, _17227_);
  and (_24868_, _17229_, _27355_);
  and (_17230_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_17231_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_17232_, _17231_, _17230_);
  and (_24869_, _17232_, _27355_);
  and (_17233_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_17234_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_17235_, _17234_, _17233_);
  and (_24870_, _17235_, _27355_);
  and (_17236_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_17237_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_17238_, _17237_, _17236_);
  and (_24871_, _17238_, _27355_);
  and (_17239_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_17240_, _16432_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_17241_, _17240_, _17239_);
  and (_24872_, _17241_, _27355_);
  and (_17242_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17243_, _01830_, _16438_);
  or (_17244_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_17245_, _17244_, _16431_);
  and (_17246_, _17245_, _17243_);
  or (_17247_, _17246_, _17242_);
  and (_24873_, _17247_, _27355_);
  and (_17248_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17249_, _01926_, _16438_);
  or (_17250_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_17251_, _17250_, _16431_);
  and (_17252_, _17251_, _17249_);
  or (_17253_, _17252_, _17248_);
  and (_24875_, _17253_, _27355_);
  and (_17254_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17255_, _02104_, _16438_);
  or (_17256_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_17257_, _17256_, _16431_);
  and (_17258_, _17257_, _17255_);
  or (_17259_, _17258_, _17254_);
  and (_24876_, _17259_, _27355_);
  and (_17260_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17261_, _01784_, _16438_);
  or (_17262_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_17263_, _17262_, _16431_);
  and (_17264_, _17263_, _17261_);
  or (_17265_, _17264_, _17260_);
  and (_24877_, _17265_, _27355_);
  and (_17266_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17267_, _01880_, _16438_);
  or (_17268_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_17269_, _17268_, _16431_);
  and (_17270_, _17269_, _17267_);
  or (_17271_, _17270_, _17266_);
  and (_24878_, _17271_, _27355_);
  and (_17272_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17273_, _02000_, _16438_);
  or (_17274_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_17275_, _17274_, _16431_);
  and (_17276_, _17275_, _17273_);
  or (_17277_, _17276_, _17272_);
  and (_24879_, _17277_, _27355_);
  and (_17278_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17279_, _02029_, _16438_);
  or (_17280_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_17281_, _17280_, _16431_);
  and (_17282_, _17281_, _17279_);
  or (_17283_, _17282_, _17278_);
  and (_24880_, _17283_, _27355_);
  and (_17284_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17285_, _01721_, _16438_);
  or (_17286_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_17287_, _17286_, _16431_);
  and (_17289_, _17287_, _17285_);
  or (_17290_, _17289_, _17284_);
  and (_24881_, _17290_, _27355_);
  and (_17291_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_17292_, _17291_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17293_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _16431_);
  and (_17294_, _17293_, _27355_);
  and (_24882_, _17294_, _17292_);
  and (_17295_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_17296_, _17295_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17298_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _16431_);
  and (_17299_, _17298_, _27355_);
  and (_24883_, _17299_, _17296_);
  and (_17300_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_17301_, _17300_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17302_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _16431_);
  and (_17303_, _17302_, _27355_);
  and (_24884_, _17303_, _17301_);
  and (_17304_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_17305_, _17304_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17307_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _16431_);
  and (_17308_, _17307_, _27355_);
  and (_24886_, _17308_, _17305_);
  and (_17309_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_17310_, _17309_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17311_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _16431_);
  and (_17312_, _17311_, _27355_);
  and (_24887_, _17312_, _17310_);
  and (_17313_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_17314_, _17313_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17316_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _16431_);
  and (_17317_, _17316_, _27355_);
  and (_24888_, _17317_, _17314_);
  and (_17318_, _16438_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_17319_, _17318_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17320_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _16431_);
  and (_17321_, _17320_, _27355_);
  and (_24889_, _17321_, _17319_);
  nand (_17322_, _16445_, _25562_);
  or (_17323_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_17325_, _17323_, _27355_);
  and (_24890_, _17325_, _17322_);
  or (_17326_, _16450_, _25639_);
  or (_17327_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_17328_, _17327_, _27355_);
  and (_24891_, _17328_, _17326_);
  nand (_17329_, _16445_, _25704_);
  or (_17330_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_17331_, _17330_, _27355_);
  and (_24892_, _17331_, _17329_);
  nand (_17333_, _16445_, _25769_);
  or (_17334_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_17335_, _17334_, _27355_);
  and (_24893_, _17335_, _17333_);
  or (_17336_, _16450_, _25830_);
  or (_17337_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_17338_, _17337_, _27355_);
  and (_24894_, _17338_, _17336_);
  or (_17339_, _16450_, _25898_);
  or (_17340_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_17341_, _17340_, _27355_);
  and (_24895_, _17341_, _17339_);
  nand (_17342_, _16445_, _25963_);
  or (_17343_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_17344_, _17343_, _27355_);
  and (_24897_, _17344_, _17342_);
  or (_17345_, _16450_, _25441_);
  or (_17346_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_17347_, _17346_, _27355_);
  and (_24898_, _17347_, _17345_);
  or (_17348_, _16450_, _26713_);
  or (_17349_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_17350_, _17349_, _27355_);
  and (_24899_, _17350_, _17348_);
  nand (_17351_, _16445_, _26745_);
  or (_17352_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_17353_, _17352_, _27355_);
  and (_24900_, _17353_, _17351_);
  nand (_17354_, _16445_, _26775_);
  or (_17355_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_17356_, _17355_, _27355_);
  and (_24901_, _17356_, _17354_);
  nand (_17357_, _16445_, _26808_);
  or (_17358_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_17359_, _17358_, _27355_);
  and (_24902_, _17359_, _17357_);
  or (_17360_, _16450_, _26837_);
  or (_17361_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_17362_, _17361_, _27355_);
  and (_24903_, _17362_, _17360_);
  or (_17363_, _16450_, _26867_);
  or (_17364_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_17365_, _17364_, _27355_);
  and (_24904_, _17365_, _17363_);
  nand (_17366_, _16445_, _26898_);
  or (_17367_, _16445_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_17368_, _17367_, _27355_);
  and (_24905_, _17368_, _17366_);
  nor (_25154_, _01762_, rst);
  and (_17369_, _01671_, _01654_);
  nand (_17370_, _17369_, _26543_);
  or (_17371_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_17372_, _17371_, _27355_);
  and (_25156_, _17372_, _17370_);
  not (_17373_, _01672_);
  nor (_17374_, _17373_, _26543_);
  and (_17375_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_17376_, _17375_, _01656_);
  or (_17377_, _17376_, _17374_);
  or (_17378_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_17379_, _17378_, _27355_);
  and (_25157_, _17379_, _17377_);
  and (_17380_, _01668_, _01654_);
  not (_17381_, _17380_);
  nor (_17382_, _17381_, _26543_);
  and (_17383_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_17384_, _17383_, _17382_);
  and (_25158_, _17384_, _27355_);
  and (_17385_, _01676_, _01654_);
  not (_17386_, _17385_);
  and (_17387_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_17388_, _17386_, _26543_);
  or (_17389_, _17388_, _17387_);
  and (_25159_, _17389_, _27355_);
  and (_17390_, _01678_, _01654_);
  not (_17391_, _17390_);
  nor (_17392_, _17391_, _26543_);
  and (_17393_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or (_17394_, _17393_, _17392_);
  and (_25160_, _17394_, _27355_);
  nand (_17395_, _01673_, _01654_);
  or (_17396_, _17395_, _01682_);
  or (_17397_, _01676_, _01668_);
  or (_17398_, _17397_, _01678_);
  and (_17399_, _17398_, _01654_);
  or (_17400_, _17399_, _17396_);
  and (_17401_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  not (_17402_, _26543_);
  and (_17403_, _01679_, _01654_);
  and (_17404_, _17403_, _17402_);
  or (_17405_, _17404_, _17401_);
  and (_25161_, _17405_, _27355_);
  and (_17406_, _01663_, _01654_);
  not (_17407_, _17406_);
  and (_17408_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_17409_, _17407_, _26543_);
  or (_17410_, _17409_, _17408_);
  and (_25162_, _17410_, _27355_);
  and (_17411_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  not (_17412_, _01651_);
  nor (_17413_, _17412_, _00755_);
  and (_17414_, _17413_, _01654_);
  not (_17415_, _17414_);
  nor (_17416_, _17415_, _26543_);
  or (_17417_, _17416_, _17411_);
  and (_25163_, _17417_, _27355_);
  nand (_17418_, _17369_, _26521_);
  or (_17419_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_17420_, _17419_, _17418_);
  and (_25261_, _17420_, _27355_);
  nand (_17421_, _17369_, _26512_);
  or (_17422_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_17423_, _17422_, _27355_);
  and (_25262_, _17423_, _17421_);
  nand (_17424_, _17369_, _26505_);
  or (_17425_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_17426_, _17425_, _27355_);
  and (_25263_, _17426_, _17424_);
  nand (_17427_, _17369_, _26497_);
  or (_17428_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_17429_, _17428_, _27355_);
  and (_25264_, _17429_, _17427_);
  nand (_17430_, _17369_, _26489_);
  or (_17431_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_17432_, _17431_, _27355_);
  and (_25265_, _17432_, _17430_);
  nand (_17433_, _17369_, _26482_);
  or (_17434_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_17435_, _17434_, _27355_);
  and (_25267_, _17435_, _17433_);
  nand (_17436_, _17369_, _26475_);
  or (_17437_, _17369_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_17438_, _17437_, _27355_);
  and (_25268_, _17438_, _17436_);
  nor (_17439_, _01656_, _26521_);
  and (_17440_, _17439_, _01672_);
  nand (_17441_, _01672_, _01654_);
  and (_17442_, _17441_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_17443_, _17442_, _17440_);
  and (_25269_, _17443_, _27355_);
  nor (_17444_, _17373_, _26512_);
  and (_17445_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_17446_, _17445_, _01656_);
  or (_17447_, _17446_, _17444_);
  or (_17448_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_17449_, _17448_, _27355_);
  and (_25270_, _17449_, _17447_);
  nor (_17450_, _17373_, _26505_);
  and (_17451_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_17452_, _17451_, _01656_);
  or (_17453_, _17452_, _17450_);
  or (_17454_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_17455_, _17454_, _27355_);
  and (_25271_, _17455_, _17453_);
  nor (_17456_, _17373_, _26497_);
  and (_17457_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_17458_, _17457_, _01656_);
  or (_17459_, _17458_, _17456_);
  or (_17460_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_17461_, _17460_, _27355_);
  and (_25272_, _17461_, _17459_);
  nor (_17462_, _17373_, _26489_);
  and (_17463_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_17464_, _17463_, _01656_);
  or (_17465_, _17464_, _17462_);
  or (_17466_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_17467_, _17466_, _27355_);
  and (_25273_, _17467_, _17465_);
  nor (_17468_, _17373_, _26482_);
  and (_17469_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_17470_, _17469_, _01656_);
  or (_17471_, _17470_, _17468_);
  or (_17472_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_17473_, _17472_, _27355_);
  and (_25274_, _17473_, _17471_);
  nor (_17474_, _17373_, _26475_);
  and (_17475_, _17373_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_17476_, _17475_, _01656_);
  or (_17477_, _17476_, _17474_);
  or (_17478_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_17479_, _17478_, _27355_);
  and (_25275_, _17479_, _17477_);
  or (_17480_, _01674_, _01656_);
  and (_17481_, _17480_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand (_17482_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_17483_, _17482_, _01673_);
  and (_17484_, _17380_, _26522_);
  or (_17485_, _17484_, _17483_);
  or (_17486_, _17485_, _17481_);
  and (_25276_, _17486_, _27355_);
  nor (_17487_, _17381_, _26512_);
  and (_17488_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_17489_, _17488_, _17487_);
  and (_25278_, _17489_, _27355_);
  and (_17490_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_17491_, _17381_, _26505_);
  or (_17492_, _17491_, _17490_);
  and (_25279_, _17492_, _27355_);
  nor (_17493_, _17381_, _26497_);
  and (_17494_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_17495_, _17494_, _17493_);
  and (_25280_, _17495_, _27355_);
  and (_17496_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_17497_, _17381_, _26489_);
  or (_17498_, _17497_, _17496_);
  and (_25281_, _17498_, _27355_);
  nor (_17499_, _17381_, _26482_);
  and (_17500_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_17501_, _17500_, _17499_);
  and (_25282_, _17501_, _27355_);
  nor (_17502_, _17381_, _26475_);
  and (_17503_, _17381_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_17504_, _17503_, _17502_);
  and (_25283_, _17504_, _27355_);
  and (_17505_, _17439_, _01676_);
  and (_17506_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_17507_, _17506_, _17505_);
  and (_25284_, _17507_, _27355_);
  nor (_17508_, _17386_, _26512_);
  and (_17509_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_17510_, _17509_, _17508_);
  and (_25285_, _17510_, _27355_);
  nor (_17511_, _17386_, _26505_);
  and (_17512_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_17513_, _17512_, _17511_);
  and (_25286_, _17513_, _27355_);
  nor (_17514_, _17386_, _26497_);
  and (_17515_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_17516_, _17515_, _17514_);
  and (_25287_, _17516_, _27355_);
  nor (_17517_, _17386_, _26489_);
  and (_17518_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_17519_, _17518_, _17517_);
  and (_25289_, _17519_, _27355_);
  nor (_17520_, _17386_, _26482_);
  and (_17521_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_17522_, _17521_, _17520_);
  and (_25290_, _17522_, _27355_);
  nor (_17523_, _17386_, _26475_);
  and (_17524_, _17386_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_17525_, _17524_, _17523_);
  and (_25291_, _17525_, _27355_);
  and (_17526_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_17527_, _17439_, _01678_);
  or (_17528_, _17527_, _17526_);
  and (_25292_, _17528_, _27355_);
  and (_17529_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_17530_, _17391_, _26512_);
  or (_17531_, _17530_, _17529_);
  and (_25293_, _17531_, _27355_);
  and (_17532_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_17533_, _17391_, _26505_);
  or (_17534_, _17533_, _17532_);
  and (_25294_, _17534_, _27355_);
  nor (_17535_, _17391_, _26497_);
  and (_17536_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_17537_, _17536_, _17535_);
  and (_25295_, _17537_, _27355_);
  nor (_17538_, _17391_, _26489_);
  and (_17539_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or (_17540_, _17539_, _17538_);
  and (_25296_, _17540_, _27355_);
  nor (_17541_, _17391_, _26482_);
  and (_17542_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_17543_, _17542_, _17541_);
  and (_25297_, _17543_, _27355_);
  nor (_17544_, _17391_, _26475_);
  and (_17545_, _17391_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_17546_, _17545_, _17544_);
  and (_25298_, _17546_, _27355_);
  and (_17547_, _17396_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_17548_, _17439_, _01679_);
  and (_17549_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_17550_, _17549_, _17398_);
  or (_17551_, _17550_, _17548_);
  or (_17552_, _17551_, _17547_);
  and (_25300_, _17552_, _27355_);
  and (_17553_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  not (_17554_, _26512_);
  and (_17555_, _17403_, _17554_);
  or (_17556_, _17555_, _17553_);
  and (_25301_, _17556_, _27355_);
  and (_17557_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_17558_, _17403_, _27805_);
  or (_17559_, _17558_, _17557_);
  and (_25302_, _17559_, _27355_);
  and (_17560_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_17561_, _17403_, _27827_);
  or (_17562_, _17561_, _17560_);
  and (_25303_, _17562_, _27355_);
  and (_17563_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_17564_, _17403_, _27829_);
  or (_17565_, _17564_, _17563_);
  and (_25304_, _17565_, _27355_);
  and (_17566_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_17567_, _17403_, _27840_);
  or (_17568_, _17567_, _17566_);
  and (_25305_, _17568_, _27355_);
  and (_17569_, _17400_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_17570_, _17403_, _27852_);
  or (_17571_, _17570_, _17569_);
  and (_25306_, _17571_, _27355_);
  and (_17572_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_17573_, _17439_, _01663_);
  or (_17574_, _17573_, _17572_);
  and (_25307_, _17574_, _27355_);
  not (_17575_, _01674_);
  or (_17576_, _01684_, _17575_);
  and (_17577_, _17576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_17578_, _17407_, _26512_);
  nand (_17579_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_17580_, _17579_, _01681_);
  or (_17581_, _17580_, _17578_);
  or (_17582_, _17581_, _17577_);
  and (_25308_, _17582_, _27355_);
  and (_17583_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_17584_, _17407_, _26505_);
  or (_17585_, _17584_, _17583_);
  and (_25309_, _17585_, _27355_);
  nor (_17586_, _17407_, _26497_);
  nor (_17587_, _01681_, _01656_);
  or (_17588_, _17587_, _17576_);
  and (_17589_, _17588_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or (_17590_, _17589_, _17586_);
  and (_25311_, _17590_, _27355_);
  and (_17591_, _17407_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_17592_, _17407_, _26489_);
  or (_17593_, _17592_, _17591_);
  and (_25312_, _17593_, _27355_);
  nor (_17594_, _17407_, _26482_);
  and (_17595_, _17588_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_17596_, _17595_, _17594_);
  and (_25313_, _17596_, _27355_);
  nor (_17597_, _17407_, _26475_);
  and (_17598_, _17588_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_17599_, _17598_, _17597_);
  and (_25314_, _17599_, _27355_);
  nand (_17600_, _01677_, _01674_);
  or (_17601_, _01685_, _17600_);
  and (_17602_, _17601_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_17603_, _01660_, _26521_);
  nand (_17604_, _01680_, _01665_);
  and (_17605_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_17606_, _17605_, _17604_);
  or (_17607_, _17606_, _17603_);
  or (_17608_, _17607_, _17602_);
  and (_25315_, _17608_, _27355_);
  and (_17609_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_17610_, _17415_, _26512_);
  or (_17611_, _17610_, _17609_);
  and (_25316_, _17611_, _27355_);
  nor (_17612_, _01660_, _26505_);
  and (_17613_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_17614_, _17613_, _17612_);
  and (_25317_, _17614_, _27355_);
  and (_17615_, _17601_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_17616_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_17617_, _17616_, _17604_);
  nor (_17618_, _01660_, _26497_);
  or (_17619_, _17618_, _17617_);
  or (_17620_, _17619_, _17615_);
  and (_25318_, _17620_, _27355_);
  nor (_17621_, _01660_, _26489_);
  and (_17622_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_17623_, _17622_, _17621_);
  and (_25319_, _17623_, _27355_);
  and (_17624_, _01660_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_17625_, _17415_, _26482_);
  or (_17626_, _17625_, _17624_);
  and (_25320_, _17626_, _27355_);
  and (_17627_, _17601_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_17628_, _01654_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_17629_, _17628_, _17604_);
  nor (_17630_, _01660_, _26475_);
  or (_17631_, _17630_, _17629_);
  or (_17632_, _17631_, _17627_);
  and (_25322_, _17632_, _27355_);
  not (_17633_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_17634_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_17635_, _17634_, _17633_);
  and (_17636_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _27355_);
  and (_25387_, _17636_, _17635_);
  nor (_17637_, _17635_, rst);
  nand (_17638_, _17634_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_17639_, _17634_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_17640_, _17639_, _17638_);
  and (_25388_, _17640_, _17637_);
  nor (_17641_, _02004_, _02053_);
  and (_17642_, _01811_, _02142_);
  and (_17643_, _17642_, _01907_);
  and (_17644_, _17643_, _17641_);
  and (_17645_, _17644_, _27034_);
  nor (_17646_, _17645_, _15901_);
  not (_17647_, _01854_);
  and (_17648_, _01952_, _17647_);
  and (_17649_, _17648_, _27840_);
  or (_17650_, _17649_, _02129_);
  nor (_17651_, _01952_, _01854_);
  and (_17652_, _17651_, _17402_);
  and (_17653_, _01952_, _01854_);
  and (_17654_, _17653_, _27829_);
  not (_17655_, _01952_);
  and (_17656_, _17655_, _01854_);
  and (_17657_, _17656_, _27852_);
  or (_17658_, _17657_, _17654_);
  or (_17659_, _17658_, _17652_);
  or (_17660_, _17659_, _17650_);
  not (_17661_, _02129_);
  and (_17662_, _17648_, _17554_);
  or (_17663_, _17662_, _17661_);
  and (_17664_, _17651_, _27827_);
  and (_17665_, _17653_, _26522_);
  and (_17666_, _17656_, _27805_);
  or (_17667_, _17666_, _17665_);
  or (_17668_, _17667_, _17664_);
  or (_17669_, _17668_, _17663_);
  nand (_17670_, _17669_, _17660_);
  nor (_17671_, _17670_, _17646_);
  not (_17672_, _02053_);
  and (_17673_, _02004_, _17672_);
  not (_17674_, _01907_);
  and (_17675_, _17642_, _17674_);
  and (_17676_, _17675_, _17673_);
  or (_17677_, _27115_, _27100_);
  nand (_17678_, _27115_, _27100_);
  nand (_17679_, _17678_, _17677_);
  nand (_17680_, _27071_, _27070_);
  nand (_17681_, _27088_, _17680_);
  or (_17682_, _27088_, _17680_);
  and (_17683_, _17682_, _17681_);
  nand (_17684_, _17683_, _17679_);
  or (_17685_, _17683_, _17679_);
  nand (_17686_, _17685_, _17684_);
  or (_17687_, _27135_, _27125_);
  nand (_17688_, _27135_, _27125_);
  nand (_17689_, _17688_, _17687_);
  nand (_17690_, _27146_, _27060_);
  or (_17691_, _27146_, _27060_);
  and (_17692_, _17691_, _17690_);
  nand (_17693_, _17692_, _17689_);
  or (_17694_, _17692_, _17689_);
  nand (_17695_, _17694_, _17693_);
  nand (_17696_, _17695_, _17686_);
  or (_17697_, _17695_, _17686_);
  nand (_17698_, _17697_, _17696_);
  nand (_17699_, _17698_, _02129_);
  or (_17700_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_17701_, _17700_, _17653_);
  and (_17702_, _17701_, _17699_);
  and (_17703_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_17704_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_17705_, _17704_, _17703_);
  and (_17706_, _17705_, _17661_);
  and (_17707_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_17708_, _02129_, _26928_);
  or (_17709_, _17708_, _17707_);
  and (_17710_, _17709_, _17651_);
  and (_17711_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_17712_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_17713_, _17712_, _17711_);
  and (_17714_, _17713_, _02129_);
  or (_17715_, _17714_, _17710_);
  or (_17716_, _17715_, _17706_);
  or (_17717_, _17716_, _17702_);
  and (_17718_, _17717_, _17676_);
  not (_17719_, _17642_);
  and (_17720_, _17673_, _01907_);
  or (_17721_, _17720_, _17719_);
  nor (_17722_, _01811_, _01748_);
  and (_17723_, _17722_, _01907_);
  and (_17724_, _17723_, _17673_);
  not (_17725_, _01811_);
  and (_17726_, _02053_, _02142_);
  nand (_17727_, _17726_, _17725_);
  nand (_17728_, _17727_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_17729_, _17728_, _17724_);
  and (_17730_, _17729_, _17721_);
  and (_17731_, _17675_, _17641_);
  and (_17732_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_17733_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_17734_, _17733_, _17732_);
  and (_17735_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_17736_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_17737_, _17736_, _17735_);
  or (_17738_, _17737_, _17734_);
  and (_17739_, _17738_, _17731_);
  and (_17740_, _17722_, _17674_);
  nor (_17741_, _02004_, _17672_);
  and (_17742_, _17741_, _17740_);
  and (_17743_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_17744_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_17745_, _17744_, _17743_);
  and (_17746_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_17747_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_17748_, _17747_, _17746_);
  or (_17749_, _17748_, _17745_);
  and (_17750_, _17749_, _17742_);
  or (_17751_, _17750_, _17739_);
  and (_17752_, _17751_, _02129_);
  or (_17753_, _17752_, _17730_);
  and (_17754_, _15895_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  nor (_17755_, _15349_, _26307_);
  and (_17756_, _17755_, _15420_);
  nor (_17757_, _15418_, _26402_);
  and (_17758_, _26327_, _26374_);
  not (_17759_, _17758_);
  and (_17760_, _17759_, _17757_);
  and (_17761_, _26281_, _26322_);
  nor (_17762_, _17761_, _26347_);
  not (_17763_, _15351_);
  and (_17764_, _17763_, _26321_);
  and (_17765_, _17764_, _17762_);
  and (_17766_, _17765_, _17760_);
  and (_17767_, _17766_, _15673_);
  and (_17768_, _17767_, _17756_);
  and (_17769_, _17768_, _26305_);
  nor (_17770_, _17769_, _26393_);
  or (_17771_, _17770_, p2_in[4]);
  not (_17772_, _17770_);
  or (_17773_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_17774_, _17773_, _17771_);
  and (_17775_, _17774_, _17653_);
  or (_17776_, _17775_, _02129_);
  or (_17777_, _17770_, p2_in[7]);
  or (_17778_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_17779_, _17778_, _17777_);
  and (_17780_, _17779_, _17651_);
  or (_17781_, _17770_, p2_in[5]);
  or (_17782_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_17783_, _17782_, _17781_);
  and (_17784_, _17783_, _17648_);
  or (_17785_, _17770_, p2_in[6]);
  or (_17786_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_17787_, _17786_, _17785_);
  and (_17788_, _17787_, _17656_);
  or (_17789_, _17788_, _17784_);
  or (_17790_, _17789_, _17780_);
  or (_17791_, _17790_, _17776_);
  and (_17792_, _17741_, _17643_);
  nor (_17793_, _17770_, p2_in[0]);
  and (_17794_, _17770_, _27415_);
  nor (_17795_, _17794_, _17793_);
  and (_17796_, _17795_, _17653_);
  or (_17797_, _17796_, _17661_);
  or (_17798_, _17770_, p2_in[2]);
  or (_17799_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_17800_, _17799_, _17798_);
  and (_17801_, _17800_, _17656_);
  or (_17802_, _17770_, p2_in[1]);
  or (_17803_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_17804_, _17803_, _17802_);
  and (_17805_, _17804_, _17648_);
  or (_17806_, _17770_, p2_in[3]);
  or (_17807_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_17808_, _17807_, _17806_);
  and (_17809_, _17808_, _17651_);
  or (_17810_, _17809_, _17805_);
  or (_17811_, _17810_, _17801_);
  or (_17812_, _17811_, _17797_);
  and (_17813_, _17812_, _17792_);
  and (_17814_, _17813_, _17791_);
  or (_17815_, _17814_, _17754_);
  and (_17816_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_17817_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_17818_, _17817_, _17816_);
  and (_17819_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_17820_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_17821_, _17820_, _17819_);
  or (_17822_, _17821_, _17818_);
  and (_17823_, _17822_, _17742_);
  and (_17825_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_17826_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_17827_, _17826_, _17825_);
  and (_17828_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_17829_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_17830_, _17829_, _17828_);
  or (_17831_, _17830_, _17827_);
  and (_17832_, _17831_, _17731_);
  or (_17833_, _17832_, _17823_);
  and (_17834_, _17833_, _17661_);
  and (_17835_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_17836_, _17835_, _02129_);
  and (_17837_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_17838_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_17839_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_17840_, _17839_, _17838_);
  or (_17841_, _17840_, _17837_);
  or (_17842_, _17841_, _17836_);
  and (_17843_, _02004_, _02053_);
  and (_17844_, _17740_, _17843_);
  and (_17845_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_17846_, _17845_, _17661_);
  and (_17847_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_17848_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_17849_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_17850_, _17849_, _17848_);
  or (_17851_, _17850_, _17847_);
  or (_17852_, _17851_, _17846_);
  and (_17853_, _17852_, _17844_);
  and (_17854_, _17853_, _17842_);
  or (_17855_, _17854_, _17834_);
  or (_17856_, _17855_, _17815_);
  or (_17857_, _17856_, _17753_);
  or (_17858_, _17770_, p0_in[2]);
  or (_17859_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_17860_, _17859_, _17858_);
  and (_17861_, _17860_, _17656_);
  nor (_17862_, _17770_, p0_in[0]);
  and (_17863_, _17770_, _27220_);
  nor (_17864_, _17863_, _17862_);
  and (_17865_, _17864_, _17653_);
  or (_17866_, _17865_, _17861_);
  or (_17867_, _17770_, p0_in[3]);
  or (_17868_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_17869_, _17868_, _17867_);
  and (_17870_, _17869_, _17651_);
  or (_17871_, _17770_, p0_in[1]);
  or (_17872_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_17873_, _17872_, _17871_);
  and (_17874_, _17873_, _17648_);
  or (_17875_, _17874_, _17870_);
  or (_17876_, _17875_, _17866_);
  and (_17877_, _17876_, _17643_);
  or (_17878_, _17770_, p1_in[3]);
  or (_17879_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_17880_, _17879_, _17878_);
  and (_17881_, _17880_, _17651_);
  or (_17882_, _17770_, p1_in[1]);
  or (_17883_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_17884_, _17883_, _17882_);
  and (_17885_, _17884_, _17648_);
  or (_17886_, _17885_, _17881_);
  or (_17887_, _17770_, p1_in[2]);
  or (_17888_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_17889_, _17888_, _17887_);
  and (_17890_, _17889_, _17656_);
  nor (_17891_, _17770_, p1_in[0]);
  and (_17892_, _17770_, _27321_);
  nor (_17893_, _17892_, _17891_);
  and (_17894_, _17893_, _17653_);
  or (_17895_, _17894_, _17890_);
  or (_17896_, _17895_, _17886_);
  and (_17897_, _17896_, _17675_);
  or (_17898_, _17897_, _17877_);
  and (_17899_, _17898_, _02129_);
  or (_17900_, _17770_, p1_in[6]);
  or (_17901_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_17902_, _17901_, _17900_);
  and (_17903_, _17902_, _17656_);
  or (_17904_, _17770_, p1_in[4]);
  or (_17905_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_17906_, _17905_, _17904_);
  and (_17907_, _17906_, _17653_);
  or (_17908_, _17907_, _17903_);
  or (_17909_, _17770_, p1_in[7]);
  or (_17910_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_17911_, _17910_, _17909_);
  and (_17912_, _17911_, _17651_);
  or (_17913_, _17770_, p1_in[5]);
  or (_17914_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_17915_, _17914_, _17913_);
  and (_17916_, _17915_, _17648_);
  or (_17917_, _17916_, _17912_);
  or (_17918_, _17917_, _17908_);
  and (_17919_, _17918_, _17675_);
  or (_17920_, _17770_, p0_in[6]);
  or (_17921_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_17922_, _17921_, _17920_);
  and (_17923_, _17922_, _17656_);
  or (_17924_, _17770_, p0_in[4]);
  or (_17925_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_17926_, _17925_, _17924_);
  and (_17927_, _17926_, _17653_);
  or (_17928_, _17927_, _17923_);
  or (_17929_, _17770_, p0_in[7]);
  or (_17930_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_17931_, _17930_, _17929_);
  and (_17932_, _17931_, _17651_);
  or (_17933_, _17770_, p0_in[5]);
  or (_17934_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_17935_, _17934_, _17933_);
  and (_17936_, _17935_, _17648_);
  or (_17937_, _17936_, _17932_);
  or (_17938_, _17937_, _17928_);
  and (_17939_, _17938_, _17643_);
  or (_17940_, _17939_, _17919_);
  and (_17941_, _17940_, _17661_);
  or (_17942_, _17941_, _17899_);
  and (_17943_, _17942_, _17843_);
  and (_17944_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_17945_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_17946_, _17945_, _17944_);
  and (_17947_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_17948_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_17949_, _17948_, _17947_);
  or (_17950_, _17949_, _17946_);
  and (_17951_, _17950_, _17741_);
  and (_17952_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_17953_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_17954_, _17953_, _17952_);
  and (_17955_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_17956_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_17957_, _17956_, _17955_);
  or (_17958_, _17957_, _17954_);
  and (_17959_, _17958_, _17843_);
  or (_17960_, _17959_, _17951_);
  and (_17961_, _17960_, _02129_);
  and (_17962_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_17963_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_17964_, _17963_, _17962_);
  and (_17965_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_17966_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_17967_, _17966_, _17965_);
  or (_17968_, _17967_, _17964_);
  and (_17969_, _17968_, _17843_);
  and (_17970_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_17971_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_17972_, _17971_, _17970_);
  and (_17973_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_17974_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_17975_, _17974_, _17973_);
  or (_17976_, _17975_, _17972_);
  and (_17977_, _17976_, _17741_);
  or (_17978_, _17977_, _17969_);
  and (_17979_, _17978_, _17661_);
  or (_17980_, _17979_, _17961_);
  and (_17981_, _17980_, _17723_);
  nor (_17982_, _17770_, p3_in[0]);
  and (_17983_, _17770_, _27499_);
  nor (_17984_, _17983_, _17982_);
  and (_17985_, _17984_, _17653_);
  or (_17986_, _17985_, _17661_);
  or (_17987_, _17770_, p3_in[2]);
  or (_17988_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_17989_, _17988_, _17987_);
  and (_17990_, _17989_, _17656_);
  or (_17991_, _17770_, p3_in[3]);
  or (_17992_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_17993_, _17992_, _17991_);
  and (_17994_, _17993_, _17651_);
  or (_17995_, _17770_, p3_in[1]);
  or (_17996_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_17997_, _17996_, _17995_);
  and (_17998_, _17997_, _17648_);
  or (_17999_, _17998_, _17994_);
  or (_18000_, _17999_, _17990_);
  or (_18001_, _18000_, _17986_);
  and (_18002_, _17741_, _17675_);
  or (_18003_, _17770_, p3_in[4]);
  or (_18004_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_18005_, _18004_, _18003_);
  and (_18006_, _18005_, _17653_);
  or (_18007_, _18006_, _02129_);
  or (_18008_, _17770_, p3_in[6]);
  or (_18009_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_18010_, _18009_, _18008_);
  and (_18011_, _18010_, _17656_);
  or (_18012_, _17770_, p3_in[7]);
  or (_18013_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_18014_, _18013_, _18012_);
  and (_18015_, _18014_, _17651_);
  or (_18016_, _17770_, p3_in[5]);
  or (_18017_, _17772_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_18018_, _18017_, _18016_);
  and (_18019_, _18018_, _17648_);
  or (_18020_, _18019_, _18015_);
  or (_18021_, _18020_, _18011_);
  or (_18022_, _18021_, _18007_);
  and (_18023_, _18022_, _18002_);
  and (_18024_, _18023_, _18001_);
  and (_18025_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_18026_, _18025_, _02129_);
  and (_18027_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_18028_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_18029_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_18030_, _18029_, _18028_);
  or (_18031_, _18030_, _18027_);
  or (_18032_, _18031_, _18026_);
  and (_18033_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_18034_, _18033_, _17661_);
  and (_18035_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_18036_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_18037_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_18038_, _18037_, _18036_);
  or (_18039_, _18038_, _18035_);
  or (_18040_, _18039_, _18034_);
  and (_18041_, _18040_, _17724_);
  and (_18042_, _18041_, _18032_);
  and (_18043_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_18044_, _18043_, _02129_);
  and (_18045_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_18046_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_18047_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_18048_, _18047_, _18046_);
  or (_18049_, _18048_, _18045_);
  or (_18050_, _18049_, _18044_);
  and (_18051_, _17656_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_18052_, _18051_, _17661_);
  and (_18053_, _17648_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_18054_, _17653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_18055_, _17651_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_18056_, _18055_, _18054_);
  or (_18057_, _18056_, _18053_);
  or (_18058_, _18057_, _18052_);
  and (_18059_, _18058_, _17644_);
  and (_18060_, _18059_, _18050_);
  or (_18061_, _18060_, _18042_);
  or (_18062_, _18061_, _18024_);
  or (_18063_, _18062_, _17981_);
  or (_18064_, _18063_, _17943_);
  or (_18065_, _18064_, _17857_);
  or (_18066_, _18065_, _17718_);
  nand (_18067_, _17754_, _25514_);
  and (_18068_, _18067_, _17646_);
  and (_18069_, _18068_, _18066_);
  or (_18070_, _18069_, _17671_);
  and (_25389_, _18070_, _27355_);
  and (_18071_, _02129_, _01811_);
  and (_18072_, _18071_, _17653_);
  and (_18073_, _01907_, _02142_);
  and (_18074_, _18073_, _17641_);
  and (_18075_, _18074_, _18072_);
  and (_18076_, _18075_, _27034_);
  and (_18077_, _17651_, _17661_);
  not (_18078_, _18077_);
  and (_18079_, _18078_, _27048_);
  and (_18080_, _18079_, _15882_);
  nor (_18081_, _18080_, _18076_);
  and (_18082_, _18081_, _15898_);
  and (_18083_, _17843_, _18073_);
  and (_18084_, _18071_, _17651_);
  and (_18085_, _18084_, _18083_);
  and (_18086_, _18085_, _26591_);
  and (_18087_, _17674_, _02004_);
  and (_18088_, _18072_, _02142_);
  and (_18089_, _18088_, _17672_);
  and (_18090_, _18089_, _18087_);
  and (_18091_, _18090_, _26933_);
  and (_18092_, _18075_, _27044_);
  or (_18093_, _18092_, _18091_);
  nor (_18094_, _18093_, _18086_);
  nor (_18095_, _18094_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_18096_, _18095_);
  and (_18097_, _18096_, _18082_);
  and (_18098_, _18071_, _17656_);
  and (_18099_, _18098_, _18083_);
  and (_18100_, _18099_, _26591_);
  or (_18101_, _18100_, rst);
  nor (_25391_, _18101_, _18097_);
  not (_18102_, _18100_);
  not (_18103_, _18090_);
  and (_18104_, _02129_, _17725_);
  and (_18105_, _18104_, _17651_);
  and (_18106_, _18105_, _18083_);
  and (_18107_, _18104_, _17653_);
  and (_18108_, _18087_, _17726_);
  and (_18109_, _18108_, _18107_);
  nor (_18110_, _18109_, _18106_);
  and (_18111_, _18107_, _18083_);
  nor (_18112_, _02129_, _01811_);
  and (_18113_, _18112_, _17653_);
  and (_18114_, _18113_, _18083_);
  nor (_18115_, _18114_, _18111_);
  and (_18116_, _18115_, _18110_);
  and (_18117_, _17741_, _18073_);
  and (_18118_, _18117_, _18107_);
  and (_18119_, _18112_, _17648_);
  and (_18120_, _18119_, _18083_);
  nor (_18121_, _18120_, _18118_);
  and (_18122_, _18104_, _17656_);
  and (_18123_, _18122_, _18083_);
  and (_18124_, _18104_, _17648_);
  and (_18125_, _18124_, _18108_);
  nor (_18126_, _18125_, _18123_);
  and (_18127_, _18126_, _18121_);
  and (_18128_, _18127_, _18116_);
  and (_18129_, _18128_, _18103_);
  and (_18130_, _17673_, _18073_);
  and (_18131_, _18130_, _18113_);
  and (_18132_, _18130_, _18105_);
  and (_18133_, _18077_, _01811_);
  and (_18134_, _18133_, _18083_);
  or (_18135_, _18134_, _18132_);
  nor (_18136_, _18135_, _18131_);
  and (_18137_, _18130_, _18119_);
  and (_18138_, _18130_, _18122_);
  nor (_18139_, _18138_, _18137_);
  nor (_18140_, _01907_, _02004_);
  and (_18141_, _18140_, _17726_);
  nand (_18142_, _18141_, _18133_);
  not (_18143_, _18071_);
  nand (_18144_, _18083_, _17648_);
  or (_18145_, _18144_, _18143_);
  and (_18146_, _18145_, _18142_);
  and (_18147_, _18146_, _18139_);
  not (_18148_, _18104_);
  or (_18149_, _18144_, _18148_);
  nor (_18150_, _18099_, _18085_);
  and (_18151_, _18150_, _18149_);
  and (_18152_, _18130_, _18107_);
  not (_18153_, _17673_);
  and (_18154_, _18088_, _18153_);
  nor (_18155_, _18154_, _18152_);
  and (_18156_, _18155_, _18151_);
  and (_18157_, _18156_, _18147_);
  and (_18158_, _18157_, _18136_);
  and (_18159_, _18158_, _18129_);
  not (_18160_, _18159_);
  nand (_18161_, _18160_, _18097_);
  and (_18162_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_18163_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_18164_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_18165_, _18164_, _18163_);
  and (_18166_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_18167_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_18168_, _18167_, _18166_);
  or (_18169_, _18168_, _18165_);
  and (_18170_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_18171_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_18172_, _18171_, _18170_);
  and (_18173_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_18174_, _18141_, _18133_);
  and (_18175_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_18176_, _18175_, _18173_);
  or (_18177_, _18176_, _18172_);
  or (_18178_, _18177_, _18169_);
  and (_18179_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_18180_, _18124_, _18083_);
  and (_18181_, _18180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_18182_, _18181_, _18179_);
  and (_18183_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_18184_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_18185_, _18184_, _18183_);
  or (_18186_, _18185_, _18182_);
  and (_18187_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_18188_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_18189_, _18188_, _18187_);
  and (_18190_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_18191_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_18192_, _18191_, _18190_);
  or (_18193_, _18192_, _18189_);
  or (_18194_, _18193_, _18186_);
  or (_18195_, _18194_, _18178_);
  and (_18196_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_18197_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_18198_, _18197_, _18196_);
  and (_18199_, _18140_, _18089_);
  and (_18200_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_18201_, _18071_, _17648_);
  and (_18202_, _18201_, _18083_);
  and (_18203_, _18202_, _26545_);
  or (_18204_, _18203_, _18200_);
  or (_18205_, _18204_, _18198_);
  and (_18206_, _18083_, _18072_);
  and (_18207_, _18206_, _17931_);
  and (_18208_, _18108_, _18072_);
  and (_18209_, _18208_, _17911_);
  or (_18210_, _18209_, _18207_);
  and (_18211_, _18141_, _18072_);
  and (_18212_, _18211_, _18014_);
  and (_18213_, _18117_, _18072_);
  and (_18214_, _18213_, _17779_);
  or (_18215_, _18214_, _18212_);
  or (_18216_, _18215_, _18210_);
  or (_18217_, _18216_, _18205_);
  and (_18218_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_18219_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_18220_, _18219_, _18218_);
  or (_18221_, _18220_, _18217_);
  or (_18222_, _18221_, _18195_);
  and (_18223_, _18222_, _18097_);
  or (_18224_, _18223_, _18162_);
  and (_18225_, _18224_, _18102_);
  and (_18226_, _18100_, _25441_);
  or (_18227_, _18226_, _18225_);
  and (_25392_, _18227_, _27355_);
  nor (_25485_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_18228_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_18229_, _17634_, rst);
  and (_25486_, _18229_, _18228_);
  nor (_18230_, _17634_, _17633_);
  or (_18231_, _18230_, _17635_);
  and (_18232_, _17638_, _27355_);
  and (_25487_, _18232_, _18231_);
  or (_18233_, _18103_, _17698_);
  nand (_18234_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_18235_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_18236_, _18235_, _18234_);
  nand (_18237_, _18206_, _17864_);
  nand (_18238_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_18239_, _18238_, _18237_);
  and (_18240_, _18239_, _18236_);
  nand (_18241_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand (_18242_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_18243_, _18242_, _18241_);
  nand (_18244_, _18211_, _17984_);
  nand (_18245_, _18213_, _17795_);
  and (_18246_, _18245_, _18244_);
  and (_18247_, _18246_, _18243_);
  and (_18248_, _18247_, _18240_);
  nand (_18249_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_18250_, _18208_, _17893_);
  nand (_18251_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_18252_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_18253_, _18252_, _18251_);
  and (_18254_, _18253_, _18250_);
  and (_18255_, _18254_, _18249_);
  and (_18256_, _18255_, _18248_);
  nand (_18257_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand (_18258_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_18259_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_18260_, _18259_, _18258_);
  and (_18261_, _18260_, _18257_);
  nand (_18262_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_18263_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_18264_, _18263_, _18262_);
  nand (_18265_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_18266_, _18145_, _26553_);
  and (_18267_, _18266_, _18265_);
  and (_18268_, _18267_, _18264_);
  nand (_18269_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_18270_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_18271_, _18270_, _18269_);
  nand (_18272_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_18273_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_18274_, _18273_, _18272_);
  and (_18275_, _18274_, _18271_);
  nand (_18276_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_18277_, _18149_, _27720_);
  and (_18278_, _18277_, _18276_);
  and (_18279_, _18278_, _18275_);
  and (_18280_, _18279_, _18268_);
  and (_18281_, _18280_, _18261_);
  and (_18282_, _18281_, _18256_);
  nand (_18283_, _18282_, _18233_);
  and (_18284_, _18283_, _18097_);
  and (_18285_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_18286_, _18285_, _18100_);
  or (_18287_, _18286_, _18284_);
  nand (_18288_, _18100_, _25562_);
  and (_18289_, _18288_, _27355_);
  and (_25488_, _18289_, _18287_);
  and (_18290_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_18291_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_18292_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_18293_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_18294_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_18295_, _18294_, _18293_);
  or (_18296_, _18295_, _18292_);
  or (_18297_, _18296_, _18291_);
  or (_18298_, _18297_, _18290_);
  and (_18299_, _18213_, _17804_);
  and (_18300_, _18211_, _17997_);
  or (_18301_, _18300_, _18299_);
  and (_18302_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_18303_, _18208_, _17884_);
  or (_18304_, _18303_, _18302_);
  or (_18305_, _18304_, _18301_);
  and (_18306_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_18307_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_18308_, _18307_, _18306_);
  or (_18309_, _18308_, _18305_);
  and (_18310_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_18311_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_18312_, _18311_, _18310_);
  and (_18313_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_18314_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_18315_, _18314_, _18313_);
  or (_18316_, _18315_, _18312_);
  and (_18317_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_18318_, _18206_, _17873_);
  or (_18319_, _18318_, _18317_);
  and (_18320_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_18321_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_18322_, _18321_, _18320_);
  or (_18323_, _18322_, _18319_);
  or (_18324_, _18323_, _18316_);
  or (_18325_, _18324_, _18309_);
  and (_18326_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_18327_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_18328_, _18149_, _27701_);
  or (_18329_, _18328_, _18327_);
  or (_18330_, _18329_, _18326_);
  and (_18331_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_18332_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_18333_, _18332_, _18331_);
  and (_18334_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_18335_, _18145_, _26559_);
  or (_18336_, _18335_, _18334_);
  or (_18337_, _18336_, _18333_);
  or (_18338_, _18337_, _18330_);
  or (_18339_, _18338_, _18325_);
  or (_18340_, _18339_, _18298_);
  and (_18341_, _18340_, _18097_);
  and (_18342_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_18343_, _18342_, _18341_);
  or (_18344_, _18343_, _18100_);
  or (_18345_, _18102_, _25639_);
  and (_18346_, _18345_, _27355_);
  and (_25489_, _18346_, _18344_);
  and (_18347_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_18348_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_18349_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_18350_, _18349_, _18348_);
  and (_18351_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_18352_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_18353_, _18352_, _18351_);
  or (_18354_, _18353_, _18350_);
  and (_18355_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_18356_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_18357_, _18356_, _18355_);
  and (_18358_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_18359_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_18360_, _18359_, _18358_);
  or (_18361_, _18360_, _18357_);
  or (_18362_, _18361_, _18354_);
  and (_18363_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_18364_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_18365_, _18364_, _18363_);
  and (_18366_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_18367_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_18368_, _18367_, _18366_);
  or (_18369_, _18368_, _18365_);
  and (_18370_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_18371_, _18180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_18372_, _18371_, _18370_);
  and (_18373_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_18374_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_18375_, _18374_, _18373_);
  or (_18376_, _18375_, _18372_);
  or (_18377_, _18376_, _18369_);
  or (_18378_, _18377_, _18362_);
  and (_18379_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_18380_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_18381_, _18380_, _18379_);
  and (_18382_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_18383_, _18202_, _02108_);
  or (_18384_, _18383_, _18382_);
  or (_18385_, _18384_, _18381_);
  and (_18386_, _18211_, _17989_);
  and (_18387_, _18213_, _17800_);
  or (_18388_, _18387_, _18386_);
  and (_18389_, _18206_, _17860_);
  and (_18390_, _18208_, _17889_);
  or (_18391_, _18390_, _18389_);
  or (_18392_, _18391_, _18388_);
  or (_18393_, _18392_, _18385_);
  and (_18394_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_18395_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_18396_, _18395_, _18394_);
  or (_18397_, _18396_, _18393_);
  or (_18398_, _18397_, _18378_);
  and (_18399_, _18398_, _18097_);
  or (_18400_, _18399_, _18100_);
  or (_18401_, _18400_, _18347_);
  nand (_18402_, _18100_, _25704_);
  and (_18403_, _18402_, _27355_);
  and (_25490_, _18403_, _18401_);
  and (_18404_, _18208_, _17880_);
  and (_18405_, _18206_, _17869_);
  and (_18406_, _18213_, _17808_);
  or (_18407_, _18406_, _18405_);
  or (_18408_, _18407_, _18404_);
  and (_18409_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_18410_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_18411_, _18410_, _18409_);
  and (_18412_, _18211_, _17993_);
  nor (_18413_, _18145_, _26571_);
  or (_18414_, _18413_, _18412_);
  or (_18415_, _18414_, _18411_);
  or (_18416_, _18415_, _18408_);
  and (_18417_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_18418_, _18180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_18419_, _18418_, _18417_);
  and (_18420_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_18421_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_18422_, _18421_, _18420_);
  or (_18423_, _18422_, _18419_);
  and (_18424_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_18425_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_18426_, _18425_, _18424_);
  and (_18427_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_18428_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_18429_, _18428_, _18427_);
  or (_18430_, _18429_, _18426_);
  or (_18431_, _18430_, _18423_);
  and (_18432_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_18433_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_18434_, _18433_, _18432_);
  and (_18435_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_18436_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_18437_, _18436_, _18435_);
  or (_18438_, _18437_, _18434_);
  and (_18439_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_18440_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_18441_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_18442_, _18441_, _18440_);
  or (_18443_, _18442_, _18439_);
  and (_18444_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_18445_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_18446_, _18445_, _18444_);
  and (_18447_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_18448_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_18449_, _18448_, _18447_);
  or (_18450_, _18449_, _18446_);
  or (_18451_, _18450_, _18443_);
  or (_18452_, _18451_, _18438_);
  or (_18453_, _18452_, _18431_);
  or (_18454_, _18453_, _18416_);
  and (_18455_, _18454_, _18097_);
  and (_18456_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_18457_, _18456_, _18455_);
  or (_18458_, _18457_, _18100_);
  nand (_18459_, _18100_, _25769_);
  and (_18460_, _18459_, _27355_);
  and (_25492_, _18460_, _18458_);
  and (_18461_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_18462_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_18463_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_18464_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_18465_, _18464_, _18463_);
  and (_18466_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_18467_, _18466_, _18465_);
  or (_18468_, _18467_, _18462_);
  or (_18469_, _18468_, _18461_);
  and (_18470_, _18208_, _17906_);
  and (_18471_, _18206_, _17926_);
  or (_18472_, _18471_, _18470_);
  and (_18473_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_18474_, _18213_, _17774_);
  or (_18475_, _18474_, _18473_);
  or (_18476_, _18475_, _18472_);
  and (_18477_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_18478_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_18479_, _18478_, _18477_);
  or (_18480_, _18479_, _18476_);
  and (_18481_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_18482_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_18483_, _18482_, _18481_);
  and (_18484_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_18485_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_18486_, _18485_, _18484_);
  or (_18487_, _18486_, _18483_);
  and (_18488_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_18489_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_18490_, _18489_, _18488_);
  and (_18491_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_18492_, _18211_, _18005_);
  or (_18493_, _18492_, _18491_);
  or (_18494_, _18493_, _18490_);
  or (_18495_, _18494_, _18487_);
  or (_18496_, _18495_, _18480_);
  nor (_18497_, _18149_, _27580_);
  and (_18498_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_18499_, _18145_, _26577_);
  or (_18500_, _18499_, _18498_);
  or (_18501_, _18500_, _18497_);
  and (_18502_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_18503_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_18504_, _18503_, _18502_);
  and (_18505_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_18506_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_18507_, _18506_, _18505_);
  or (_18508_, _18507_, _18504_);
  or (_18509_, _18508_, _18501_);
  or (_18510_, _18509_, _18496_);
  or (_18511_, _18510_, _18469_);
  and (_18512_, _18511_, _18097_);
  and (_18513_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_18514_, _18513_, _18512_);
  or (_18515_, _18514_, _18100_);
  or (_18516_, _18102_, _25830_);
  and (_18517_, _18516_, _27355_);
  and (_25493_, _18517_, _18515_);
  and (_18518_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18519_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_18520_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_18521_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_18522_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_18523_, _18522_, _18521_);
  or (_18524_, _18523_, _18520_);
  or (_18525_, _18524_, _18519_);
  or (_18526_, _18525_, _18518_);
  and (_18527_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_18528_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_18529_, _18528_, _18527_);
  and (_18530_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_18531_, _18208_, _17915_);
  or (_18532_, _18531_, _18530_);
  or (_18533_, _18532_, _18529_);
  and (_18534_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_18535_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_18536_, _18535_, _18534_);
  or (_18537_, _18536_, _18533_);
  and (_18538_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_18539_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_18540_, _18539_, _18538_);
  and (_18541_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_18542_, _18211_, _18018_);
  or (_18543_, _18542_, _18541_);
  or (_18544_, _18543_, _18540_);
  and (_18545_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_18546_, _18213_, _17783_);
  or (_18547_, _18546_, _18545_);
  and (_18548_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_18549_, _18206_, _17935_);
  or (_18550_, _18549_, _18548_);
  or (_18551_, _18550_, _18547_);
  or (_18552_, _18551_, _18544_);
  or (_18553_, _18552_, _18537_);
  and (_18554_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_18555_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_18556_, _18145_, _26583_);
  or (_18557_, _18556_, _18555_);
  or (_18558_, _18557_, _18554_);
  and (_18559_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_18560_, _18149_, _27582_);
  or (_18561_, _18560_, _18559_);
  and (_18562_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_18563_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_18564_, _18563_, _18562_);
  or (_18565_, _18564_, _18561_);
  or (_18566_, _18565_, _18558_);
  or (_18567_, _18566_, _18553_);
  or (_18568_, _18567_, _18526_);
  and (_18569_, _18568_, _18097_);
  and (_18570_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_18571_, _18570_, _18569_);
  or (_18572_, _18571_, _18100_);
  or (_18573_, _18102_, _25898_);
  and (_18574_, _18573_, _27355_);
  and (_25494_, _18574_, _18572_);
  nand (_18575_, _18100_, _25963_);
  and (_18576_, _18575_, _27355_);
  and (_18577_, _18161_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_18578_, _18090_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_18579_, _18199_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_18580_, _18114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_18581_, _18125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_18582_, _18099_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_18583_, _18582_, _18581_);
  or (_18584_, _18583_, _18580_);
  or (_18585_, _18584_, _18579_);
  or (_18586_, _18585_, _18578_);
  and (_18587_, _18118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_18588_, _18211_, _18010_);
  or (_18589_, _18588_, _18587_);
  and (_18590_, _18123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_18591_, _18208_, _17902_);
  or (_18592_, _18591_, _18590_);
  or (_18593_, _18592_, _18589_);
  and (_18594_, _18152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_18595_, _18134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_18596_, _18595_, _18594_);
  or (_18597_, _18596_, _18593_);
  and (_18598_, _18120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_18599_, _18109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_18600_, _18599_, _18598_);
  and (_18601_, _18111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_18602_, _18075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_18603_, _18602_, _18601_);
  or (_18604_, _18603_, _18600_);
  and (_18605_, _18085_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_18606_, _18213_, _17787_);
  or (_18607_, _18606_, _18605_);
  and (_18608_, _18106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_18609_, _18206_, _17922_);
  or (_18610_, _18609_, _18608_);
  or (_18611_, _18610_, _18607_);
  or (_18612_, _18611_, _18604_);
  or (_18613_, _18612_, _18597_);
  and (_18614_, _18174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_18615_, _18132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_18616_, _18145_, _26589_);
  or (_18617_, _18616_, _18615_);
  or (_18618_, _18617_, _18614_);
  and (_18619_, _18131_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_18620_, _18138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_18621_, _18620_, _18619_);
  and (_18622_, _18137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_18623_, _18149_, _27591_);
  or (_18624_, _18623_, _18622_);
  or (_18625_, _18624_, _18621_);
  or (_18626_, _18625_, _18618_);
  or (_18627_, _18626_, _18613_);
  or (_18628_, _18627_, _18586_);
  and (_18629_, _18628_, _18097_);
  or (_18630_, _18629_, _18577_);
  or (_18631_, _18630_, _18100_);
  and (_25495_, _18631_, _18576_);
  and (_25567_, _02141_, _27355_);
  and (_25568_, _03058_, _27355_);
  nor (_25571_, _02129_, rst);
  and (_25586_, _02983_, _27355_);
  and (_25587_, _02997_, _27355_);
  and (_25588_, _03007_, _27355_);
  and (_25589_, _03016_, _27355_);
  and (_25590_, _03026_, _27355_);
  and (_25591_, _03036_, _27355_);
  and (_25592_, _03047_, _27355_);
  nor (_25593_, _01854_, rst);
  nor (_25594_, _01952_, rst);
  nor (_18632_, _16708_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_18633_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18634_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _18633_);
  nor (_18635_, _18634_, _18632_);
  not (_18636_, _18635_);
  nor (_18637_, _16726_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18638_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _18633_);
  nor (_18639_, _18638_, _18637_);
  nor (_18640_, _18639_, _18636_);
  and (_18641_, _18640_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_18642_, _18639_, _18635_);
  and (_18643_, _18642_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_18644_, _18643_, _18641_);
  and (_18645_, _18639_, _18636_);
  and (_18646_, _18645_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_18647_, _18639_, _18635_);
  and (_18648_, _18647_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_18649_, _18648_, _18646_);
  and (_18650_, _18649_, _18644_);
  nor (_18651_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _18633_);
  nor (_18653_, _18652_, _18651_);
  nor (_18654_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18655_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _18633_);
  nor (_18656_, _18655_, _18654_);
  nor (_18657_, _18656_, _18653_);
  not (_18658_, _18657_);
  nor (_18659_, _18658_, _18650_);
  and (_18660_, _18642_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_18661_, _18647_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_18662_, _18661_, _18660_);
  and (_18663_, _18645_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_18664_, _18640_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_18665_, _18664_, _18663_);
  and (_18666_, _18665_, _18662_);
  and (_18667_, _18656_, _18653_);
  not (_18668_, _18667_);
  nor (_18669_, _18668_, _18666_);
  nor (_18670_, _18669_, _18659_);
  and (_18671_, _18642_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_18672_, _18647_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_18673_, _18672_, _18671_);
  and (_18674_, _18645_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_18675_, _18640_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_18676_, _18675_, _18674_);
  and (_18677_, _18676_, _18673_);
  not (_18678_, _18653_);
  and (_18679_, _18656_, _18678_);
  not (_18680_, _18679_);
  nor (_18681_, _18680_, _18677_);
  and (_18682_, _18640_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_18683_, _18647_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_18684_, _18683_, _18682_);
  and (_18685_, _18645_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_18686_, _18642_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_18687_, _18686_, _18685_);
  and (_18688_, _18687_, _18684_);
  not (_18689_, _18656_);
  and (_18690_, _18689_, _18653_);
  not (_18691_, _18690_);
  nor (_18692_, _18691_, _18688_);
  nor (_18693_, _18692_, _18681_);
  and (_18694_, _18693_, _18670_);
  not (_18695_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_18696_, _18653_, _18695_);
  or (_18697_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_18698_, _18697_, _18696_);
  not (_18699_, _18639_);
  and (_18700_, _18656_, _18635_);
  and (_18701_, _18700_, _18699_);
  and (_18702_, _18701_, _18698_);
  not (_18703_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_18704_, _18653_, _18703_);
  or (_18705_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_18706_, _18705_, _18704_);
  and (_18707_, _18700_, _18639_);
  and (_18708_, _18707_, _18706_);
  or (_18709_, _18708_, _18702_);
  and (_18710_, _18689_, _18635_);
  not (_18711_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_18712_, _18653_, _18711_);
  or (_18713_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_18714_, _18713_, _18712_);
  and (_18715_, _18714_, _18639_);
  not (_18716_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_18717_, _18653_, _18716_);
  or (_18718_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_18719_, _18718_, _18717_);
  and (_18720_, _18719_, _18699_);
  or (_18721_, _18720_, _18715_);
  and (_18722_, _18721_, _18710_);
  not (_18723_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_18724_, _18653_, _18723_);
  or (_18725_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_18726_, _18725_, _18724_);
  and (_18727_, _18726_, _18656_);
  not (_18728_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_18729_, _18653_, _18728_);
  or (_18730_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_18731_, _18730_, _18729_);
  and (_18732_, _18731_, _18689_);
  or (_18733_, _18732_, _18727_);
  and (_18734_, _18733_, _18639_);
  not (_18735_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_18736_, _18653_, _18735_);
  or (_18737_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_18738_, _18737_, _18736_);
  and (_18739_, _18738_, _18656_);
  not (_18740_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_18741_, _18653_, _18740_);
  or (_18742_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_18743_, _18742_, _18741_);
  and (_18744_, _18743_, _18689_);
  nor (_18745_, _18744_, _18739_);
  nor (_18746_, _18745_, _18639_);
  or (_18747_, _18746_, _18734_);
  and (_18748_, _18747_, _18636_);
  or (_18749_, _18748_, _18722_);
  nor (_18750_, _18749_, _18709_);
  nor (_18751_, _18750_, _18694_);
  and (_18752_, _18694_, word_in[7]);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _18752_, _18751_);
  and (_18753_, _18667_, _18635_);
  nor (_18754_, _18753_, _18699_);
  and (_18755_, _18667_, _18640_);
  nor (_18756_, _18755_, _18754_);
  nor (_18757_, _18667_, _18635_);
  nor (_18758_, _18757_, _18753_);
  not (_18759_, _18758_);
  and (_18760_, _18759_, _18756_);
  and (_18761_, _18760_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_18762_, _18761_);
  not (_18763_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand (_18764_, _18756_, _18763_);
  nor (_18765_, _18756_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_18766_, _18765_, _18759_);
  and (_18767_, _18766_, _18764_);
  nor (_18768_, _18758_, _18756_);
  and (_18769_, _18768_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_18770_, _18769_, _18767_);
  and (_18771_, _18770_, _18762_);
  nor (_18772_, _18771_, _18658_);
  and (_18773_, _18760_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_18774_, _18773_);
  not (_18775_, _18756_);
  or (_18776_, _18775_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_18777_, _18756_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_18778_, _18777_, _18759_);
  and (_18779_, _18778_, _18776_);
  and (_18780_, _18768_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_18781_, _18780_, _18779_);
  and (_18782_, _18781_, _18774_);
  nor (_18783_, _18782_, _18680_);
  nor (_18784_, _18783_, _18772_);
  and (_18785_, _18760_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_18786_, _18785_);
  not (_18787_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand (_18788_, _18756_, _18787_);
  nor (_18789_, _18756_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_18790_, _18789_, _18759_);
  and (_18791_, _18790_, _18788_);
  and (_18792_, _18768_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_18793_, _18792_, _18791_);
  and (_18794_, _18793_, _18786_);
  nor (_18795_, _18794_, _18668_);
  and (_18796_, _18760_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_18797_, _18796_);
  not (_18798_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand (_18799_, _18756_, _18798_);
  nor (_18800_, _18756_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_18801_, _18800_, _18759_);
  and (_18802_, _18801_, _18799_);
  and (_18803_, _18768_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_18804_, _18803_, _18802_);
  and (_18805_, _18804_, _18797_);
  nor (_18806_, _18805_, _18691_);
  nor (_18807_, _18806_, _18795_);
  and (_18808_, _18807_, _18784_);
  or (_18809_, _18667_, _18657_);
  not (_18810_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_18811_, _18653_, _18810_);
  or (_18812_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_18813_, _18812_, _18811_);
  and (_18814_, _18813_, _18809_);
  not (_18815_, _18809_);
  and (_18816_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor (_18817_, _18653_, _18735_);
  or (_18818_, _18817_, _18816_);
  and (_18819_, _18818_, _18815_);
  or (_18820_, _18819_, _18814_);
  or (_18821_, _18820_, _18758_);
  not (_18822_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_18823_, _18653_, _18822_);
  or (_18824_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_18825_, _18824_, _18823_);
  and (_18826_, _18825_, _18809_);
  not (_18827_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_18828_, _18653_, _18827_);
  or (_18829_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_18830_, _18829_, _18828_);
  and (_18831_, _18830_, _18815_);
  nor (_18832_, _18831_, _18826_);
  nand (_18833_, _18832_, _18758_);
  and (_18834_, _18833_, _18756_);
  and (_18835_, _18834_, _18821_);
  not (_18836_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_18837_, _18653_, _18836_);
  or (_18838_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_18839_, _18838_, _18837_);
  and (_18840_, _18839_, _18809_);
  not (_18841_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_18842_, _18653_, _18841_);
  or (_18843_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_18844_, _18843_, _18842_);
  and (_18845_, _18844_, _18815_);
  or (_18846_, _18845_, _18840_);
  or (_18847_, _18846_, _18758_);
  not (_18848_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_18849_, _18653_, _18848_);
  or (_18850_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_18851_, _18850_, _18849_);
  and (_18852_, _18851_, _18809_);
  not (_18853_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_18854_, _18653_, _18853_);
  or (_18855_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_18856_, _18855_, _18854_);
  and (_18857_, _18856_, _18815_);
  nor (_18858_, _18857_, _18852_);
  nand (_18859_, _18858_, _18758_);
  nand (_18860_, _18859_, _18847_);
  nor (_18861_, _18860_, _18756_);
  nor (_18862_, _18861_, _18835_);
  nor (_18863_, _18862_, _18808_);
  and (_18864_, _18808_, word_in[15]);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _18864_, _18863_);
  not (_18865_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_18866_, _18701_);
  or (_18867_, _18700_, _18699_);
  and (_18868_, _18867_, _18866_);
  and (_18869_, _18868_, _18865_);
  and (_18870_, _18689_, _18642_);
  nor (_18871_, _18707_, _18870_);
  not (_18872_, _18871_);
  nor (_18873_, _18689_, _18635_);
  nor (_18874_, _18873_, _18710_);
  and (_18875_, _18874_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_18876_, _18875_, _18872_);
  nor (_18877_, _18876_, _18869_);
  and (_18878_, _18868_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_18879_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_18880_, _18868_, _18879_);
  nor (_18881_, _18880_, _18878_);
  nor (_18882_, _18881_, _18636_);
  nor (_18883_, _18882_, _18877_);
  nor (_18884_, _18883_, _18656_);
  and (_18885_, _18868_, _18763_);
  not (_18886_, _18873_);
  not (_18887_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_18888_, _18639_, _18887_);
  nor (_18889_, _18888_, _18886_);
  not (_18891_, _18889_);
  nor (_18892_, _18891_, _18885_);
  not (_18894_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_18895_, _18868_, _18894_);
  and (_18897_, _18700_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_18898_, _18897_, _18707_);
  nor (_18900_, _18898_, _18895_);
  or (_18901_, _18900_, _18678_);
  or (_18903_, _18901_, _18892_);
  nor (_18904_, _18903_, _18884_);
  not (_18906_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_18907_, _18868_, _18906_);
  and (_18909_, _18874_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_18910_, _18909_, _18872_);
  nor (_18912_, _18910_, _18907_);
  and (_18913_, _18868_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_18915_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_18916_, _18868_, _18915_);
  nor (_18918_, _18916_, _18913_);
  nor (_18919_, _18918_, _18636_);
  nor (_18921_, _18919_, _18912_);
  nor (_18922_, _18921_, _18656_);
  and (_18924_, _18868_, _18787_);
  not (_18925_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_18927_, _18639_, _18925_);
  nor (_18928_, _18927_, _18886_);
  not (_18929_, _18928_);
  nor (_18930_, _18929_, _18924_);
  not (_18931_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_18932_, _18868_, _18931_);
  and (_18933_, _18700_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_18934_, _18933_, _18707_);
  nor (_18935_, _18934_, _18932_);
  or (_18936_, _18935_, _18653_);
  or (_18937_, _18936_, _18930_);
  nor (_18938_, _18937_, _18922_);
  nor (_18939_, _18938_, _18904_);
  or (_18940_, _18738_, _18656_);
  or (_18941_, _18743_, _18689_);
  and (_18942_, _18941_, _18940_);
  and (_18943_, _18942_, _18874_);
  and (_18944_, _18710_, _18698_);
  and (_18945_, _18719_, _18873_);
  or (_18946_, _18945_, _18944_);
  or (_18947_, _18946_, _18943_);
  and (_18948_, _18947_, _18868_);
  or (_18949_, _18726_, _18656_);
  or (_18950_, _18731_, _18689_);
  and (_18951_, _18950_, _18949_);
  and (_18952_, _18951_, _18874_);
  and (_18953_, _18710_, _18706_);
  and (_18954_, _18714_, _18873_);
  or (_18955_, _18954_, _18953_);
  nor (_18956_, _18955_, _18952_);
  nor (_18957_, _18956_, _18868_);
  or (_18958_, _18957_, _18948_);
  and (_18959_, _18958_, _18939_);
  not (_18960_, _18939_);
  and (_18961_, _18960_, word_in[23]);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _18961_, _18959_);
  and (_18962_, _18658_, _18635_);
  nor (_18963_, _18658_, _18635_);
  nor (_18964_, _18963_, _18962_);
  and (_18965_, _18962_, _18639_);
  nor (_18966_, _18962_, _18639_);
  nor (_18967_, _18966_, _18965_);
  nor (_18968_, _18967_, _18865_);
  and (_18969_, _18967_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_18970_, _18969_, _18968_);
  nor (_18971_, _18970_, _18964_);
  nand (_18972_, _18967_, _18879_);
  not (_18973_, _18964_);
  nor (_18974_, _18967_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_18975_, _18974_, _18973_);
  and (_18976_, _18975_, _18972_);
  nor (_18977_, _18976_, _18971_);
  nor (_18978_, _18977_, _18658_);
  nor (_18979_, _18967_, \oc8051_symbolic_cxrom1.regvalid [5]);
  not (_18980_, _18979_);
  nor (_18981_, _18973_, _18888_);
  and (_18982_, _18981_, _18980_);
  nor (_18983_, _18967_, _18894_);
  and (_18985_, _18967_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_18987_, _18985_, _18983_);
  nor (_18988_, _18987_, _18964_);
  nor (_18990_, _18988_, _18982_);
  nor (_18991_, _18990_, _18680_);
  nor (_18993_, _18991_, _18978_);
  nor (_18994_, _18967_, _18906_);
  and (_18996_, _18967_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_18997_, _18996_, _18994_);
  nor (_18999_, _18997_, _18964_);
  nand (_19000_, _18967_, _18915_);
  nor (_19002_, _18967_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_19003_, _19002_, _18973_);
  and (_19005_, _19003_, _19000_);
  nor (_19006_, _19005_, _18999_);
  nor (_19008_, _19006_, _18668_);
  nor (_19009_, _18967_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not (_19011_, _19009_);
  nor (_19012_, _18973_, _18927_);
  and (_19014_, _19012_, _19011_);
  nor (_19015_, _18967_, _18931_);
  and (_19017_, _18967_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_19018_, _19017_, _19015_);
  nor (_19020_, _19018_, _18964_);
  nor (_19021_, _19020_, _19014_);
  nor (_19022_, _19021_, _18691_);
  nor (_19023_, _19022_, _19008_);
  and (_19024_, _19023_, _18993_);
  and (_19025_, _18844_, _18809_);
  and (_19026_, _18839_, _18815_);
  or (_19027_, _19026_, _19025_);
  or (_19028_, _19027_, _18964_);
  and (_19029_, _18856_, _18809_);
  and (_19030_, _18851_, _18815_);
  nor (_19031_, _19030_, _19029_);
  nand (_19032_, _19031_, _18964_);
  and (_19033_, _19032_, _19028_);
  and (_19034_, _19033_, _18967_);
  not (_19035_, _18967_);
  and (_19036_, _18818_, _18809_);
  and (_19037_, _18813_, _18815_);
  nor (_19038_, _19037_, _19036_);
  nor (_19039_, _19038_, _18964_);
  and (_19040_, _18830_, _18809_);
  and (_19041_, _18825_, _18815_);
  or (_19042_, _19041_, _19040_);
  and (_19043_, _19042_, _18964_);
  or (_19044_, _19043_, _19039_);
  and (_19045_, _19044_, _19035_);
  nor (_19046_, _19045_, _19034_);
  nor (_19047_, _19046_, _19024_);
  and (_19048_, _19024_, word_in[31]);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _19048_, _19047_);
  or (_19049_, _18647_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_25618_, _19049_, _27355_);
  and (_19050_, _19024_, _27355_);
  and (_19051_, _19050_, _18967_);
  and (_19052_, _19051_, _18964_);
  and (_19053_, _19052_, _18657_);
  not (_19054_, _19053_);
  and (_19055_, _18904_, _27355_);
  and (_19056_, _19055_, _18689_);
  nor (_19057_, _18939_, rst);
  nor (_19058_, _18874_, _18699_);
  and (_19059_, _19058_, _19057_);
  and (_19060_, _19059_, _19056_);
  not (_19061_, _19060_);
  and (_19062_, _18808_, _27355_);
  and (_19063_, _19062_, _18758_);
  and (_19064_, _19063_, _18775_);
  and (_19065_, _19064_, _18679_);
  and (_19066_, _18753_, _18639_);
  and (_19067_, _18694_, _27355_);
  and (_19068_, _19067_, word_in[7]);
  and (_19069_, _19068_, _19066_);
  nand (_19070_, _19067_, _19066_);
  and (_19071_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor (_19072_, _19071_, _19069_);
  nor (_19073_, _19072_, _19065_);
  and (_19074_, _19062_, word_in[15]);
  and (_19075_, _19074_, _19065_);
  or (_19076_, _19075_, _19073_);
  and (_19077_, _19076_, _19061_);
  and (_19078_, _19060_, word_in[23]);
  or (_19079_, _19078_, _19077_);
  and (_19080_, _19079_, _19054_);
  and (_19081_, _19050_, word_in[31]);
  and (_19082_, _19081_, _19053_);
  or (_25622_, _19082_, _19080_);
  and (_19083_, _18657_, _18642_);
  or (_19084_, _18965_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_19085_, _19084_, _19083_);
  and (_25625_, _19085_, _27355_);
  or (_19086_, _19066_, _18870_);
  and (_19087_, _18679_, _18647_);
  or (_19088_, _19087_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_19089_, _19088_, _19086_);
  and (_25629_, _19089_, _27355_);
  and (_19090_, _18679_, _18642_);
  or (_19091_, _19090_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_19092_, _19091_, _19086_);
  and (_25634_, _19092_, _27355_);
  or (_19093_, _18642_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_25640_, _19093_, _27355_);
  and (_19094_, _18667_, _18642_);
  and (_19095_, _18668_, _18642_);
  and (_19096_, _19095_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_19097_, _19096_, _19094_);
  not (_19098_, _18642_);
  and (_19099_, _18657_, _18640_);
  nand (_19100_, _18966_, _18668_);
  and (_19101_, _19100_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_19102_, _19101_, _19099_);
  and (_19103_, _19102_, _19098_);
  nor (_19104_, _19103_, _19097_);
  nor (_19105_, _19104_, _18760_);
  or (_19106_, _19102_, _19096_);
  and (_19107_, _19106_, _19066_);
  and (_19108_, _18815_, _18642_);
  and (_19109_, _18870_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_19110_, _19109_, _19108_);
  or (_19111_, _19110_, _19107_);
  or (_19112_, _19111_, _19105_);
  and (_25647_, _19112_, _27355_);
  and (_19113_, _18690_, _18640_);
  or (_19114_, _19113_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_19115_, _18966_, _19066_);
  and (_19116_, _19115_, _19114_);
  or (_19117_, _19116_, _19099_);
  and (_19118_, _18690_, _18642_);
  and (_19119_, _19118_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_19120_, _19119_, _19090_);
  and (_19121_, _19083_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_19122_, _19114_, _19066_);
  or (_19123_, _19122_, _19121_);
  or (_19124_, _19123_, _19120_);
  or (_19125_, _19124_, _19094_);
  or (_19126_, _19125_, _19117_);
  and (_25655_, _19126_, _27355_);
  or (_19127_, _19094_, _19099_);
  or (_19128_, _19127_, _19113_);
  and (_19129_, _19095_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_19130_, _18700_, _18639_);
  and (_19131_, _18679_, _18640_);
  or (_19132_, _18653_, _18639_);
  nor (_19133_, _18642_, _18798_);
  and (_19134_, _19133_, _19132_);
  or (_19135_, _19134_, _19131_);
  and (_19136_, _19135_, _19130_);
  or (_19137_, _19136_, _19129_);
  or (_19138_, _19137_, _19128_);
  and (_25663_, _19138_, _27355_);
  or (_19139_, _18874_, _18639_);
  not (_19140_, _19139_);
  nor (_19141_, _19140_, _19086_);
  and (_19142_, _18664_, _18689_);
  nand (_19143_, _18680_, _18640_);
  and (_19144_, _19143_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_19145_, _19144_, _19142_);
  or (_19146_, _19145_, _18755_);
  and (_19147_, _19146_, _18775_);
  and (_19148_, _19094_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_19149_, _19148_, _19131_);
  or (_19150_, _19149_, _19142_);
  or (_19151_, _19150_, _19147_);
  and (_19152_, _19151_, _19141_);
  and (_19153_, _19145_, _19066_);
  or (_19154_, _19148_, _19099_);
  and (_19155_, _18870_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_19156_, _19090_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_19157_, _19156_, _19155_);
  or (_19158_, _19157_, _19154_);
  or (_19159_, _19158_, _19153_);
  or (_19160_, _19159_, _19113_);
  or (_19161_, _19160_, _19152_);
  and (_25673_, _19161_, _27355_);
  and (_19162_, _18815_, _18640_);
  and (_19163_, _18963_, _18639_);
  or (_19164_, _19163_, _18755_);
  or (_19165_, _19164_, _19162_);
  or (_19166_, _19165_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_25683_, _19166_, _27355_);
  not (_19167_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_19168_, _19130_, _19167_);
  and (_19169_, _18690_, _18645_);
  or (_19170_, _19169_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_19171_, _19170_, _19130_);
  or (_19172_, _19171_, _18963_);
  and (_19173_, _19172_, _18639_);
  or (_19174_, _19173_, _18755_);
  or (_19175_, _19174_, _19131_);
  or (_19176_, _19175_, _19168_);
  and (_28201_[9], _19176_, _27355_);
  or (_19177_, _19058_, _19087_);
  or (_19178_, _19177_, _19066_);
  and (_19179_, _19083_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_19180_, _18679_, _18645_);
  and (_19181_, _19108_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_19182_, _19181_, _19180_);
  or (_19183_, _19182_, _19179_);
  or (_19184_, _19127_, _19162_);
  and (_19185_, _19184_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_19186_, _19164_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_19187_, _18757_);
  and (_19188_, _19187_, _18639_);
  or (_19189_, _19188_, _19169_);
  and (_19190_, _19189_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_19191_, _19190_, _19186_);
  or (_19192_, _19191_, _19185_);
  or (_19193_, _19192_, _19183_);
  and (_19194_, _19193_, _19178_);
  not (_19195_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_19196_, _19139_, _19195_);
  and (_19197_, _19131_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_19198_, _18870_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_19199_, _19198_, _18755_);
  or (_19200_, _19199_, _19197_);
  or (_19201_, _19200_, _19196_);
  or (_19202_, _19201_, _19169_);
  or (_19203_, _19202_, _19163_);
  or (_19204_, _19203_, _19194_);
  and (_28201_[10], _19204_, _27355_);
  and (_19205_, _18667_, _18645_);
  or (_19206_, _19205_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_19207_, _19187_, _18754_);
  and (_19208_, _19207_, _19206_);
  and (_19209_, _18663_, _18689_);
  and (_19210_, _18755_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_19211_, _19210_, _19180_);
  or (_19212_, _19211_, _19209_);
  or (_19213_, _19099_, _19113_);
  and (_19214_, _19213_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_19215_, _19131_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_19216_, _19094_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_19217_, _19108_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_19218_, _19217_, _19216_);
  or (_19219_, _19218_, _19215_);
  or (_19220_, _19219_, _19214_);
  or (_19221_, _19220_, _19212_);
  or (_19222_, _19221_, _19208_);
  and (_19223_, _19222_, _19177_);
  and (_19224_, _19066_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_19225_, _19083_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_19226_, _19225_, _19163_);
  or (_19227_, _19226_, _19210_);
  or (_19228_, _19227_, _19220_);
  or (_19229_, _19228_, _19169_);
  or (_19230_, _19229_, _19224_);
  or (_19231_, _19230_, _19223_);
  and (_28201_[11], _19231_, _27355_);
  and (_19232_, _18965_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_19233_, _18690_, _18647_);
  not (_19234_, _19233_);
  and (_19235_, _19058_, _19234_);
  and (_19236_, _19108_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_19237_, _19162_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_19238_, _19237_, _19236_);
  or (_19239_, _19238_, _19235_);
  and (_19240_, _19099_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_19241_, _18963_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_19242_, _19241_, _19169_);
  or (_19243_, _19242_, _19240_);
  and (_19244_, _19094_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_19245_, _18755_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_19246_, _19245_, _19244_);
  or (_19247_, _19246_, _19243_);
  or (_19248_, _19247_, _19239_);
  or (_19249_, _19248_, _19232_);
  and (_28201_[12], _19249_, _27355_);
  or (_19250_, _19058_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_28201_[13], _19250_, _27355_);
  or (_19251_, _19207_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_28201_[14], _19251_, _27355_);
  and (_19252_, _19050_, word_in[24]);
  and (_19253_, _19050_, _18964_);
  nor (_19254_, _19051_, _19253_);
  and (_19255_, _19254_, _18690_);
  and (_19256_, _19255_, _19252_);
  and (_19257_, _19057_, _18689_);
  nor (_19258_, _19257_, _19055_);
  and (_19259_, _19258_, _19057_);
  and (_19260_, _19259_, _18872_);
  not (_19261_, _19260_);
  or (_19262_, _19261_, word_in[16]);
  and (_19263_, _19255_, _19050_);
  not (_19264_, _19263_);
  and (_19265_, _19062_, _19066_);
  and (_19266_, _19067_, word_in[0]);
  and (_19267_, _19266_, _19083_);
  not (_19268_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_19269_, _19067_, _19083_);
  nor (_19270_, _19269_, _19268_);
  or (_19271_, _19270_, _19267_);
  or (_19272_, _19271_, _19265_);
  not (_19273_, _19265_);
  or (_19274_, _19273_, word_in[8]);
  and (_19275_, _19274_, _19272_);
  or (_19276_, _19275_, _19260_);
  and (_19277_, _19276_, _19264_);
  and (_19278_, _19277_, _19262_);
  or (_28202_[0], _19278_, _19256_);
  and (_19279_, _19050_, word_in[25]);
  and (_19280_, _19279_, _19255_);
  or (_19281_, _19261_, word_in[17]);
  and (_19282_, _19062_, word_in[9]);
  and (_19283_, _19282_, _19066_);
  not (_19284_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or (_19285_, _19269_, _19284_);
  and (_19286_, _19067_, word_in[1]);
  nand (_19287_, _19286_, _19269_);
  and (_19288_, _19287_, _19285_);
  nor (_19289_, _19288_, _19265_);
  or (_19290_, _19289_, _19283_);
  or (_19291_, _19290_, _19260_);
  and (_19292_, _19291_, _19264_);
  and (_19293_, _19292_, _19281_);
  or (_28202_[1], _19293_, _19280_);
  and (_19294_, _19050_, word_in[26]);
  and (_19295_, _19294_, _19255_);
  or (_19296_, _19261_, word_in[18]);
  not (_19297_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_19298_, _19269_, _19297_);
  and (_19299_, _19067_, word_in[2]);
  and (_19300_, _19299_, _19269_);
  or (_19301_, _19300_, _19298_);
  or (_19302_, _19301_, _19265_);
  or (_19303_, _19273_, word_in[10]);
  and (_19304_, _19303_, _19302_);
  or (_19305_, _19304_, _19260_);
  and (_19306_, _19305_, _19264_);
  and (_19307_, _19306_, _19296_);
  or (_28202_[2], _19307_, _19295_);
  and (_19308_, _19050_, word_in[27]);
  and (_19309_, _19308_, _19255_);
  or (_19310_, _19261_, word_in[19]);
  not (_19311_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_19312_, _19269_, _19311_);
  and (_19313_, _19067_, word_in[3]);
  and (_19314_, _19313_, _19269_);
  or (_19315_, _19314_, _19312_);
  or (_19316_, _19315_, _19265_);
  or (_19317_, _19273_, word_in[11]);
  and (_19318_, _19317_, _19316_);
  or (_19319_, _19318_, _19260_);
  and (_19320_, _19319_, _19264_);
  and (_19321_, _19320_, _19310_);
  or (_28202_[3], _19321_, _19309_);
  and (_19322_, _19050_, word_in[28]);
  and (_19323_, _19322_, _19255_);
  or (_19324_, _19261_, word_in[20]);
  not (_19325_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_19326_, _19269_, _19325_);
  and (_19327_, _19067_, word_in[4]);
  and (_19328_, _19327_, _19083_);
  or (_19329_, _19328_, _19326_);
  or (_19330_, _19329_, _19265_);
  or (_19331_, _19273_, word_in[12]);
  and (_19332_, _19331_, _19330_);
  or (_19333_, _19332_, _19260_);
  and (_19334_, _19333_, _19264_);
  and (_19335_, _19334_, _19324_);
  or (_28202_[4], _19335_, _19323_);
  or (_19336_, _19261_, word_in[21]);
  not (_19337_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_19338_, _19269_, _19337_);
  and (_19339_, _19067_, word_in[5]);
  and (_19340_, _19339_, _19269_);
  or (_19341_, _19340_, _19338_);
  or (_19342_, _19341_, _19265_);
  or (_19343_, _19273_, word_in[13]);
  and (_19344_, _19343_, _19342_);
  or (_19345_, _19344_, _19260_);
  and (_19346_, _19345_, _19264_);
  and (_19347_, _19346_, _19336_);
  and (_19348_, _19050_, word_in[29]);
  and (_19349_, _19348_, _19263_);
  or (_28202_[5], _19349_, _19347_);
  and (_19350_, _19050_, word_in[30]);
  and (_19351_, _19350_, _19255_);
  or (_19352_, _19261_, word_in[22]);
  not (_19353_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_19354_, _19269_, _19353_);
  and (_19355_, _19067_, word_in[6]);
  and (_19356_, _19355_, _19269_);
  or (_19357_, _19356_, _19354_);
  or (_19358_, _19357_, _19265_);
  or (_19359_, _19273_, word_in[14]);
  and (_19360_, _19359_, _19358_);
  or (_19361_, _19360_, _19260_);
  and (_19362_, _19361_, _19264_);
  and (_19363_, _19362_, _19352_);
  or (_28202_[6], _19363_, _19351_);
  and (_19364_, _19255_, _19081_);
  or (_19365_, _19261_, word_in[23]);
  nor (_19366_, _19269_, _18810_);
  and (_19367_, _19269_, _19068_);
  or (_19368_, _19367_, _19366_);
  or (_19369_, _19368_, _19265_);
  or (_19370_, _19273_, word_in[15]);
  and (_19371_, _19370_, _19369_);
  or (_19372_, _19371_, _19260_);
  and (_19373_, _19372_, _19264_);
  and (_19374_, _19373_, _19365_);
  or (_28202_[7], _19374_, _19364_);
  and (_19375_, _19050_, _18679_);
  and (_19376_, _19375_, _19254_);
  and (_19377_, _19376_, _19252_);
  and (_19378_, _19057_, _18871_);
  and (_19379_, _19055_, _18656_);
  not (_19380_, _19379_);
  nor (_19381_, _19380_, _19378_);
  and (_19382_, _19062_, _19083_);
  and (_19383_, _19266_, _19118_);
  nand (_19384_, _19067_, _19118_);
  and (_19385_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or (_19386_, _19385_, _19383_);
  or (_19387_, _19386_, _19382_);
  not (_19388_, _19382_);
  or (_19389_, _19388_, word_in[8]);
  and (_19390_, _19389_, _19387_);
  or (_19391_, _19390_, _19381_);
  not (_19392_, _19376_);
  and (_19393_, _19057_, word_in[16]);
  not (_19394_, _19381_);
  or (_19395_, _19394_, _19393_);
  and (_19396_, _19395_, _19392_);
  and (_19397_, _19396_, _19391_);
  or (_28209_[0], _19397_, _19377_);
  and (_19398_, _19286_, _19118_);
  and (_19399_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_19400_, _19399_, _19398_);
  nor (_19401_, _19400_, _19382_);
  and (_19402_, _19382_, word_in[9]);
  nor (_19403_, _19402_, _19401_);
  nor (_19404_, _19403_, _19381_);
  and (_19405_, _19057_, word_in[17]);
  and (_19406_, _19381_, _19405_);
  or (_19407_, _19406_, _19376_);
  or (_19408_, _19407_, _19404_);
  or (_19409_, _19392_, _19279_);
  and (_28209_[1], _19409_, _19408_);
  and (_19410_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_19411_, _19299_, _19118_);
  nor (_19412_, _19411_, _19410_);
  nor (_19413_, _19412_, _19382_);
  and (_19414_, _19382_, word_in[10]);
  nor (_19415_, _19414_, _19413_);
  nor (_19416_, _19415_, _19381_);
  and (_19417_, _19057_, word_in[18]);
  and (_19418_, _19381_, _19417_);
  or (_19419_, _19418_, _19376_);
  or (_19420_, _19419_, _19416_);
  or (_19421_, _19392_, _19294_);
  and (_28209_[2], _19421_, _19420_);
  and (_19422_, _19313_, _19118_);
  and (_19423_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_19424_, _19423_, _19422_);
  nor (_19425_, _19424_, _19382_);
  and (_19426_, _19382_, word_in[11]);
  nor (_19427_, _19426_, _19425_);
  nor (_19428_, _19427_, _19381_);
  and (_19429_, _19057_, word_in[19]);
  and (_19430_, _19381_, _19429_);
  or (_19431_, _19430_, _19376_);
  or (_19432_, _19431_, _19428_);
  or (_19433_, _19392_, _19308_);
  and (_28209_[3], _19433_, _19432_);
  and (_19434_, _19327_, _19118_);
  and (_19435_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or (_19436_, _19435_, _19434_);
  or (_19437_, _19436_, _19382_);
  or (_19438_, _19388_, word_in[12]);
  nand (_19439_, _19438_, _19437_);
  nor (_19440_, _19439_, _19381_);
  and (_19441_, _19057_, word_in[20]);
  and (_19442_, _19381_, _19441_);
  or (_19443_, _19442_, _19376_);
  or (_19444_, _19443_, _19440_);
  or (_19445_, _19392_, word_in[28]);
  and (_28209_[4], _19445_, _19444_);
  and (_19446_, _19339_, _19118_);
  and (_19447_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or (_19448_, _19447_, _19446_);
  or (_19449_, _19448_, _19382_);
  or (_19450_, _19388_, word_in[13]);
  nand (_19451_, _19450_, _19449_);
  nor (_19452_, _19451_, _19381_);
  and (_19453_, _19057_, word_in[21]);
  and (_19454_, _19381_, _19453_);
  or (_19455_, _19454_, _19376_);
  or (_19456_, _19455_, _19452_);
  or (_19457_, _19392_, word_in[29]);
  and (_28209_[5], _19457_, _19456_);
  and (_19458_, _19355_, _19118_);
  and (_19459_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_19460_, _19459_, _19458_);
  nor (_19461_, _19460_, _19382_);
  and (_19462_, _19382_, word_in[14]);
  nor (_19463_, _19462_, _19461_);
  nor (_19464_, _19463_, _19381_);
  and (_19465_, _19057_, word_in[22]);
  and (_19466_, _19381_, _19465_);
  or (_19467_, _19466_, _19376_);
  or (_19468_, _19467_, _19464_);
  or (_19469_, _19392_, _19350_);
  and (_28209_[6], _19469_, _19468_);
  and (_19470_, _19068_, _19118_);
  and (_19471_, _19384_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_19472_, _19471_, _19470_);
  nor (_19473_, _19472_, _19382_);
  and (_19474_, _19382_, word_in[15]);
  nor (_19475_, _19474_, _19473_);
  nor (_19476_, _19475_, _19381_);
  and (_19477_, _19057_, word_in[23]);
  and (_19478_, _19381_, _19477_);
  or (_19479_, _19478_, _19376_);
  or (_19480_, _19479_, _19476_);
  or (_19481_, _19392_, _19081_);
  and (_28209_[7], _19481_, _19480_);
  and (_19482_, _19050_, _18667_);
  and (_19483_, _19482_, _19254_);
  not (_19484_, _19483_);
  not (_19485_, _19055_);
  and (_19486_, _19257_, _19485_);
  and (_19487_, _19486_, _18872_);
  and (_19488_, _19062_, _19118_);
  nand (_19489_, _19067_, _19090_);
  and (_19490_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_19491_, _19266_, _19090_);
  nor (_19492_, _19491_, _19490_);
  nor (_19493_, _19492_, _19488_);
  and (_19494_, _19488_, word_in[8]);
  nor (_19495_, _19494_, _19493_);
  nor (_19496_, _19495_, _19487_);
  and (_19497_, _19487_, _19393_);
  or (_19499_, _19497_, _19496_);
  and (_19500_, _19499_, _19484_);
  and (_19501_, _19483_, word_in[24]);
  or (_28210_[0], _19501_, _19500_);
  and (_19502_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_19503_, _19286_, _19090_);
  or (_19504_, _19503_, _19502_);
  or (_19505_, _19504_, _19488_);
  not (_19506_, _19488_);
  or (_19507_, _19506_, word_in[9]);
  nand (_19509_, _19507_, _19505_);
  nor (_19510_, _19509_, _19487_);
  and (_19511_, _19487_, _19405_);
  or (_19512_, _19511_, _19483_);
  or (_19513_, _19512_, _19510_);
  or (_19514_, _19484_, word_in[25]);
  and (_28210_[1], _19514_, _19513_);
  and (_19515_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_19516_, _19299_, _19090_);
  nor (_19517_, _19516_, _19515_);
  nor (_19519_, _19517_, _19488_);
  and (_19520_, _19488_, word_in[10]);
  nor (_19521_, _19520_, _19519_);
  nor (_19522_, _19521_, _19487_);
  and (_19523_, _19487_, _19417_);
  or (_19524_, _19523_, _19522_);
  and (_19525_, _19524_, _19484_);
  and (_19526_, _19483_, word_in[26]);
  or (_28210_[2], _19526_, _19525_);
  and (_19527_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_19529_, _19313_, _19090_);
  nor (_19530_, _19529_, _19527_);
  nor (_19531_, _19530_, _19488_);
  and (_19532_, _19488_, word_in[11]);
  nor (_19533_, _19532_, _19531_);
  nor (_19534_, _19533_, _19487_);
  and (_19535_, _19487_, _19429_);
  or (_19536_, _19535_, _19534_);
  and (_19537_, _19536_, _19484_);
  and (_19538_, _19483_, word_in[27]);
  or (_28210_[3], _19538_, _19537_);
  and (_19540_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_19541_, _19327_, _19090_);
  nor (_19542_, _19541_, _19540_);
  nor (_19543_, _19542_, _19488_);
  and (_19544_, _19488_, word_in[12]);
  nor (_19545_, _19544_, _19543_);
  nor (_19546_, _19545_, _19487_);
  and (_19547_, _19487_, _19441_);
  or (_19548_, _19547_, _19546_);
  and (_19550_, _19548_, _19484_);
  and (_19551_, _19483_, word_in[28]);
  or (_28210_[4], _19551_, _19550_);
  and (_19552_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_19553_, _19339_, _19090_);
  or (_19554_, _19553_, _19552_);
  or (_19555_, _19554_, _19488_);
  or (_19556_, _19506_, word_in[13]);
  nand (_19557_, _19556_, _19555_);
  nor (_19558_, _19557_, _19487_);
  and (_19560_, _19487_, _19453_);
  or (_19561_, _19560_, _19483_);
  or (_19562_, _19561_, _19558_);
  or (_19563_, _19484_, word_in[29]);
  and (_28210_[5], _19563_, _19562_);
  and (_19564_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_19565_, _19355_, _19090_);
  nor (_19566_, _19565_, _19564_);
  nor (_19567_, _19566_, _19488_);
  and (_19568_, _19488_, word_in[14]);
  nor (_19569_, _19568_, _19567_);
  nor (_19570_, _19569_, _19487_);
  and (_19571_, _19487_, _19465_);
  or (_19572_, _19571_, _19570_);
  and (_19573_, _19572_, _19484_);
  and (_19574_, _19483_, word_in[30]);
  or (_28210_[6], _19574_, _19573_);
  and (_19575_, _19489_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_19576_, _19068_, _19090_);
  nor (_19577_, _19576_, _19575_);
  nor (_19578_, _19577_, _19488_);
  and (_19579_, _19488_, word_in[15]);
  nor (_19580_, _19579_, _19578_);
  nor (_19581_, _19580_, _19487_);
  and (_19582_, _19487_, _19477_);
  or (_19583_, _19582_, _19581_);
  and (_19584_, _19583_, _19484_);
  and (_19585_, _19483_, word_in[31]);
  or (_28210_[7], _19585_, _19584_);
  not (_19586_, _19056_);
  nor (_19587_, _19378_, _19586_);
  and (_19588_, _19062_, _19090_);
  nand (_19589_, _19067_, _19094_);
  and (_19590_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_19591_, _19266_, _19094_);
  or (_19592_, _19591_, _19590_);
  or (_19593_, _19592_, _19588_);
  not (_19594_, _19588_);
  or (_19595_, _19594_, word_in[8]);
  and (_19596_, _19595_, _19593_);
  or (_19597_, _19596_, _19587_);
  and (_19598_, _19050_, _19083_);
  not (_19599_, _19598_);
  not (_19600_, _19587_);
  or (_19601_, _19600_, _19393_);
  and (_19602_, _19601_, _19599_);
  and (_19603_, _19602_, _19597_);
  and (_19604_, _19598_, word_in[24]);
  or (_28211_[0], _19604_, _19603_);
  and (_19605_, _19587_, _19405_);
  and (_19606_, _19286_, _19094_);
  and (_19607_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_19608_, _19607_, _19606_);
  nor (_19609_, _19608_, _19588_);
  and (_19610_, _19588_, word_in[9]);
  nor (_19611_, _19610_, _19609_);
  nor (_19612_, _19611_, _19587_);
  or (_19613_, _19612_, _19605_);
  and (_19614_, _19613_, _19599_);
  and (_19615_, _19598_, word_in[25]);
  or (_28211_[1], _19615_, _19614_);
  and (_19616_, _19587_, _19417_);
  and (_19617_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_19618_, _19299_, _19094_);
  nor (_19619_, _19618_, _19617_);
  nor (_19620_, _19619_, _19588_);
  and (_19621_, _19588_, word_in[10]);
  nor (_19622_, _19621_, _19620_);
  nor (_19623_, _19622_, _19587_);
  or (_19624_, _19623_, _19616_);
  and (_19625_, _19624_, _19599_);
  and (_19626_, _19598_, word_in[26]);
  or (_28211_[2], _19626_, _19625_);
  and (_19627_, _19598_, _19308_);
  and (_19628_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_19629_, _19313_, _19094_);
  or (_19630_, _19629_, _19628_);
  or (_19631_, _19630_, _19588_);
  or (_19632_, _19594_, word_in[11]);
  and (_19633_, _19632_, _19631_);
  or (_19634_, _19633_, _19587_);
  or (_19635_, _19600_, _19429_);
  and (_19636_, _19635_, _19599_);
  and (_19637_, _19636_, _19634_);
  or (_28211_[3], _19637_, _19627_);
  and (_19638_, _19587_, _19441_);
  and (_19639_, _19327_, _19094_);
  and (_19640_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_19641_, _19640_, _19639_);
  nor (_19642_, _19641_, _19588_);
  and (_19643_, _19588_, word_in[12]);
  nor (_19644_, _19643_, _19642_);
  nor (_19645_, _19644_, _19587_);
  or (_19646_, _19645_, _19638_);
  and (_19647_, _19646_, _19599_);
  and (_19648_, _19598_, word_in[28]);
  or (_28211_[4], _19648_, _19647_);
  and (_19649_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_19650_, _19339_, _19094_);
  or (_19651_, _19650_, _19649_);
  or (_19652_, _19651_, _19588_);
  or (_19653_, _19594_, word_in[13]);
  and (_19654_, _19653_, _19652_);
  or (_19655_, _19654_, _19587_);
  or (_19656_, _19600_, _19453_);
  and (_19657_, _19656_, _19599_);
  and (_19658_, _19657_, _19655_);
  and (_19659_, _19598_, word_in[29]);
  or (_28211_[5], _19659_, _19658_);
  and (_19660_, _19587_, _19465_);
  and (_19661_, _19355_, _19094_);
  and (_19662_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_19663_, _19662_, _19661_);
  nor (_19664_, _19663_, _19588_);
  and (_19665_, _19588_, word_in[14]);
  nor (_19666_, _19665_, _19664_);
  nor (_19667_, _19666_, _19587_);
  or (_19668_, _19667_, _19660_);
  and (_19669_, _19668_, _19599_);
  and (_19670_, _19598_, word_in[30]);
  or (_28211_[6], _19670_, _19669_);
  and (_19671_, _19587_, _19477_);
  and (_19672_, _19589_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_19673_, _19068_, _19094_);
  nor (_19674_, _19673_, _19672_);
  nor (_19675_, _19674_, _19588_);
  and (_19676_, _19588_, word_in[15]);
  nor (_19677_, _19676_, _19675_);
  nor (_19678_, _19677_, _19587_);
  or (_19679_, _19678_, _19671_);
  and (_19680_, _19679_, _19599_);
  and (_19681_, _19598_, word_in[31]);
  or (_28211_[7], _19681_, _19680_);
  and (_19682_, _19253_, _18699_);
  and (_19683_, _19682_, _18690_);
  not (_19684_, _19683_);
  and (_19685_, _19140_, _19057_);
  and (_19686_, _19685_, _19258_);
  and (_19687_, _19062_, _19094_);
  not (_19688_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_19689_, _19067_, _19099_);
  nor (_19690_, _19689_, _19688_);
  and (_19691_, _19266_, _19099_);
  nor (_19692_, _19691_, _19690_);
  nor (_19693_, _19692_, _19687_);
  and (_19694_, _19687_, word_in[8]);
  nor (_19695_, _19694_, _19693_);
  nor (_19696_, _19695_, _19686_);
  and (_19697_, _19686_, _19393_);
  or (_19698_, _19697_, _19696_);
  and (_19699_, _19698_, _19684_);
  and (_19700_, _19683_, _19252_);
  or (_28212_[0], _19700_, _19699_);
  not (_19701_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_19702_, _19689_, _19701_);
  and (_19703_, _19286_, _19099_);
  or (_19704_, _19703_, _19702_);
  or (_19705_, _19704_, _19687_);
  not (_19706_, _19687_);
  or (_19707_, _19706_, word_in[9]);
  and (_19708_, _19707_, _19705_);
  or (_19709_, _19708_, _19686_);
  not (_19710_, _19686_);
  or (_19711_, _19710_, _19405_);
  and (_19712_, _19711_, _19709_);
  or (_19713_, _19712_, _19683_);
  or (_19714_, _19684_, _19279_);
  and (_28212_[1], _19714_, _19713_);
  not (_19715_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_19716_, _19689_, _19715_);
  and (_19717_, _19299_, _19099_);
  nor (_19718_, _19717_, _19716_);
  nor (_19719_, _19718_, _19687_);
  and (_19720_, _19687_, word_in[10]);
  nor (_19721_, _19720_, _19719_);
  nor (_19722_, _19721_, _19686_);
  and (_19723_, _19686_, _19417_);
  or (_19724_, _19723_, _19722_);
  and (_19725_, _19724_, _19684_);
  and (_19726_, _19683_, _19294_);
  or (_28212_[2], _19726_, _19725_);
  not (_19727_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_19728_, _19689_, _19727_);
  and (_19729_, _19313_, _19099_);
  nor (_19730_, _19729_, _19728_);
  nor (_19731_, _19730_, _19687_);
  and (_19732_, _19687_, word_in[11]);
  nor (_19733_, _19732_, _19731_);
  nor (_19734_, _19733_, _19686_);
  and (_19735_, _19686_, _19429_);
  or (_19736_, _19735_, _19734_);
  and (_19737_, _19736_, _19684_);
  and (_19738_, _19683_, _19308_);
  or (_28212_[3], _19738_, _19737_);
  not (_19739_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_19740_, _19689_, _19739_);
  and (_19741_, _19327_, _19099_);
  nor (_19742_, _19741_, _19740_);
  nor (_19743_, _19742_, _19687_);
  and (_19744_, _19687_, word_in[12]);
  nor (_19745_, _19744_, _19743_);
  nor (_19746_, _19745_, _19686_);
  and (_19747_, _19686_, _19441_);
  or (_19748_, _19747_, _19746_);
  and (_19749_, _19748_, _19684_);
  and (_19750_, _19683_, _19322_);
  or (_28212_[4], _19750_, _19749_);
  not (_19751_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_19752_, _19689_, _19751_);
  and (_19753_, _19339_, _19099_);
  or (_19754_, _19753_, _19752_);
  or (_19755_, _19754_, _19687_);
  or (_19756_, _19706_, word_in[13]);
  and (_19757_, _19756_, _19755_);
  or (_19758_, _19757_, _19686_);
  or (_19759_, _19710_, _19453_);
  and (_19760_, _19759_, _19758_);
  or (_19761_, _19760_, _19683_);
  or (_19762_, _19684_, _19348_);
  and (_28212_[5], _19762_, _19761_);
  not (_19763_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_19764_, _19689_, _19763_);
  and (_19765_, _19355_, _19099_);
  or (_19766_, _19765_, _19764_);
  or (_19767_, _19766_, _19687_);
  or (_19768_, _19706_, word_in[14]);
  and (_19769_, _19768_, _19767_);
  or (_19770_, _19769_, _19686_);
  or (_19771_, _19710_, _19465_);
  and (_19772_, _19771_, _19770_);
  or (_19773_, _19772_, _19683_);
  or (_19774_, _19684_, _19350_);
  and (_28212_[6], _19774_, _19773_);
  nor (_19775_, _19689_, _18822_);
  and (_19776_, _19689_, _19068_);
  or (_19777_, _19776_, _19775_);
  or (_19778_, _19777_, _19687_);
  or (_19779_, _19706_, word_in[15]);
  and (_19780_, _19779_, _19778_);
  or (_19781_, _19780_, _19686_);
  or (_19782_, _19710_, _19477_);
  and (_19783_, _19782_, _19781_);
  or (_19784_, _19783_, _19683_);
  or (_19785_, _19684_, _19081_);
  and (_28212_[7], _19785_, _19784_);
  and (_19786_, _19685_, _19379_);
  not (_19787_, _19786_);
  and (_19788_, _19063_, _18756_);
  and (_19789_, _19788_, _18657_);
  not (_19790_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_19791_, _19067_, _19113_);
  nor (_19792_, _19791_, _19790_);
  and (_19793_, _19266_, _19113_);
  nor (_19794_, _19793_, _19792_);
  nor (_19795_, _19794_, _19789_);
  and (_19796_, _19062_, word_in[8]);
  and (_19797_, _19789_, _19796_);
  or (_19798_, _19797_, _19795_);
  and (_19799_, _19798_, _19787_);
  and (_19800_, _19682_, _18679_);
  and (_19801_, _19786_, _19393_);
  or (_19802_, _19801_, _19800_);
  or (_19803_, _19802_, _19799_);
  not (_19804_, _19800_);
  or (_19805_, _19804_, _19252_);
  and (_28213_[0], _19805_, _19803_);
  not (_19806_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_19807_, _19791_, _19806_);
  and (_19808_, _19286_, _19113_);
  nor (_19809_, _19808_, _19807_);
  nor (_19810_, _19809_, _19789_);
  and (_19811_, _19789_, _19282_);
  or (_19812_, _19811_, _19810_);
  or (_19813_, _19812_, _19786_);
  or (_19814_, _19787_, _19405_);
  and (_19815_, _19814_, _19804_);
  and (_19816_, _19815_, _19813_);
  and (_19817_, _19800_, _19279_);
  or (_28213_[1], _19817_, _19816_);
  not (_19818_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_19819_, _19791_, _19818_);
  and (_19820_, _19299_, _19113_);
  nor (_19821_, _19820_, _19819_);
  nor (_19822_, _19821_, _19789_);
  and (_19823_, _19062_, word_in[10]);
  and (_19824_, _19789_, _19823_);
  or (_19825_, _19824_, _19822_);
  and (_19826_, _19825_, _19787_);
  and (_19827_, _19786_, _19417_);
  or (_19828_, _19827_, _19800_);
  or (_19829_, _19828_, _19826_);
  or (_19830_, _19804_, _19294_);
  and (_28213_[2], _19830_, _19829_);
  not (_19831_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_19832_, _19791_, _19831_);
  and (_19833_, _19313_, _19113_);
  nor (_19834_, _19833_, _19832_);
  nor (_19835_, _19834_, _19789_);
  and (_19836_, _19062_, word_in[11]);
  and (_19837_, _19789_, _19836_);
  or (_19838_, _19837_, _19835_);
  and (_19839_, _19838_, _19787_);
  and (_19840_, _19786_, _19429_);
  or (_19841_, _19840_, _19800_);
  or (_19842_, _19841_, _19839_);
  or (_19843_, _19804_, _19308_);
  and (_28213_[3], _19843_, _19842_);
  not (_19844_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_19845_, _19791_, _19844_);
  and (_19846_, _19327_, _19113_);
  or (_19847_, _19846_, _19845_);
  or (_19848_, _19847_, _19789_);
  and (_19849_, _19062_, word_in[12]);
  not (_19850_, _19789_);
  or (_19851_, _19850_, _19849_);
  and (_19852_, _19851_, _19848_);
  or (_19853_, _19852_, _19786_);
  or (_19854_, _19787_, _19441_);
  and (_19855_, _19854_, _19804_);
  and (_19856_, _19855_, _19853_);
  and (_19857_, _19800_, _19322_);
  or (_28213_[4], _19857_, _19856_);
  and (_19858_, _19786_, _19453_);
  not (_19859_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_19860_, _19791_, _19859_);
  and (_19861_, _19339_, _19113_);
  nor (_19862_, _19861_, _19860_);
  nor (_19863_, _19862_, _19789_);
  and (_19864_, _19062_, word_in[13]);
  and (_19865_, _19789_, _19864_);
  or (_19866_, _19865_, _19863_);
  and (_19867_, _19866_, _19787_);
  or (_19868_, _19867_, _19858_);
  and (_19869_, _19868_, _19804_);
  and (_19870_, _19800_, _19348_);
  or (_28213_[5], _19870_, _19869_);
  not (_19871_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_19872_, _19791_, _19871_);
  and (_19873_, _19355_, _19113_);
  nor (_19874_, _19873_, _19872_);
  nor (_19875_, _19874_, _19789_);
  and (_19876_, _19062_, word_in[14]);
  and (_19877_, _19789_, _19876_);
  or (_19878_, _19877_, _19875_);
  and (_19879_, _19878_, _19787_);
  and (_19880_, _19786_, _19465_);
  or (_19881_, _19880_, _19800_);
  or (_19882_, _19881_, _19879_);
  or (_19883_, _19804_, _19350_);
  and (_28213_[6], _19883_, _19882_);
  and (_19884_, _19791_, word_in[7]);
  nor (_19885_, _19791_, _18716_);
  nor (_19886_, _19885_, _19884_);
  nor (_19887_, _19886_, _19789_);
  and (_19888_, _19789_, _19074_);
  or (_19889_, _19888_, _19887_);
  and (_19890_, _19889_, _19787_);
  and (_19891_, _19786_, _19477_);
  or (_19892_, _19891_, _19800_);
  or (_19893_, _19892_, _19890_);
  or (_19894_, _19804_, _19081_);
  and (_28213_[7], _19894_, _19893_);
  and (_19895_, _19685_, _19486_);
  and (_19896_, _19788_, _18690_);
  and (_19897_, _19067_, _19131_);
  and (_19898_, _19897_, word_in[0]);
  not (_19899_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_19900_, _19897_, _19899_);
  nor (_19901_, _19900_, _19898_);
  nor (_19902_, _19901_, _19896_);
  and (_19903_, _19896_, _19796_);
  or (_19904_, _19903_, _19902_);
  or (_19905_, _19904_, _19895_);
  and (_19906_, _19682_, _18667_);
  not (_19907_, _19906_);
  not (_19908_, _19895_);
  or (_19909_, _19908_, _19393_);
  and (_19910_, _19909_, _19907_);
  and (_19911_, _19910_, _19905_);
  and (_19912_, _19906_, _19252_);
  or (_28214_[0], _19912_, _19911_);
  not (_19913_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_19914_, _19897_, _19913_);
  and (_19915_, _19897_, _19286_);
  or (_19916_, _19915_, _19914_);
  or (_19917_, _19916_, _19896_);
  not (_19918_, _19896_);
  or (_19919_, _19918_, _19282_);
  and (_19920_, _19919_, _19917_);
  or (_19921_, _19920_, _19895_);
  or (_19922_, _19908_, _19405_);
  and (_19923_, _19922_, _19907_);
  and (_19924_, _19923_, _19921_);
  and (_19925_, _19906_, _19279_);
  or (_28214_[1], _19925_, _19924_);
  not (_19926_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_19927_, _19897_, _19926_);
  and (_19928_, _19897_, _19299_);
  or (_19929_, _19928_, _19927_);
  or (_19930_, _19929_, _19896_);
  or (_19931_, _19918_, _19823_);
  and (_19932_, _19931_, _19930_);
  or (_19933_, _19932_, _19895_);
  or (_19934_, _19908_, _19417_);
  and (_19935_, _19934_, _19933_);
  or (_19936_, _19935_, _19906_);
  or (_19937_, _19907_, _19294_);
  and (_28214_[2], _19937_, _19936_);
  or (_19938_, _19908_, _19429_);
  not (_19939_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_19940_, _19897_, _19939_);
  and (_19941_, _19897_, _19313_);
  or (_19942_, _19941_, _19940_);
  or (_19943_, _19942_, _19896_);
  or (_19944_, _19918_, _19836_);
  and (_19945_, _19944_, _19943_);
  or (_19946_, _19945_, _19895_);
  and (_19947_, _19946_, _19938_);
  or (_19948_, _19947_, _19906_);
  or (_19949_, _19907_, _19308_);
  and (_28214_[3], _19949_, _19948_);
  not (_19950_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_19951_, _19897_, _19950_);
  and (_19952_, _19897_, _19327_);
  or (_19953_, _19952_, _19951_);
  or (_19954_, _19953_, _19896_);
  or (_19955_, _19918_, _19849_);
  and (_19956_, _19955_, _19954_);
  or (_19957_, _19956_, _19895_);
  or (_19958_, _19908_, _19441_);
  and (_19959_, _19958_, _19907_);
  and (_19960_, _19959_, _19957_);
  and (_19961_, _19906_, _19322_);
  or (_28214_[4], _19961_, _19960_);
  not (_19962_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_19963_, _19897_, _19962_);
  and (_19964_, _19897_, _19339_);
  or (_19965_, _19964_, _19963_);
  or (_19966_, _19965_, _19896_);
  or (_19967_, _19918_, _19864_);
  and (_19968_, _19967_, _19966_);
  or (_19969_, _19968_, _19895_);
  or (_19970_, _19908_, _19453_);
  and (_19971_, _19970_, _19907_);
  and (_19972_, _19971_, _19969_);
  and (_19973_, _19906_, _19348_);
  or (_28214_[5], _19973_, _19972_);
  or (_19974_, _19908_, _19465_);
  not (_19975_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_19976_, _19897_, _19975_);
  and (_19977_, _19897_, _19355_);
  or (_19978_, _19977_, _19976_);
  or (_19979_, _19978_, _19896_);
  or (_19980_, _19918_, _19876_);
  and (_19981_, _19980_, _19979_);
  or (_19982_, _19981_, _19895_);
  and (_19983_, _19982_, _19974_);
  or (_19984_, _19983_, _19906_);
  or (_19985_, _19907_, _19350_);
  and (_28214_[6], _19985_, _19984_);
  nor (_19986_, _19897_, _18827_);
  and (_19987_, _19897_, _19068_);
  or (_19988_, _19987_, _19986_);
  or (_19989_, _19988_, _19896_);
  or (_19990_, _19918_, _19074_);
  and (_19991_, _19990_, _19989_);
  or (_19992_, _19991_, _19895_);
  or (_19993_, _19908_, _19477_);
  and (_19994_, _19993_, _19907_);
  and (_19995_, _19994_, _19992_);
  and (_19996_, _19906_, _19081_);
  or (_28214_[7], _19996_, _19995_);
  and (_19997_, _19252_, _19099_);
  and (_19998_, _19685_, _19056_);
  and (_19999_, _19788_, _18679_);
  and (_20000_, _19067_, _18755_);
  and (_20001_, _20000_, word_in[0]);
  not (_20002_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_20003_, _20000_, _20002_);
  nor (_20004_, _20003_, _20001_);
  nor (_20005_, _20004_, _19999_);
  and (_20006_, _19999_, _19796_);
  or (_20007_, _20006_, _20005_);
  or (_20008_, _20007_, _19998_);
  and (_20009_, _19050_, _19099_);
  not (_20010_, _20009_);
  not (_20011_, _19998_);
  or (_20012_, _20011_, _19393_);
  and (_20013_, _20012_, _20010_);
  and (_20014_, _20013_, _20008_);
  or (_28215_[0], _20014_, _19997_);
  and (_20015_, _19279_, _19099_);
  not (_20016_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_20017_, _20000_, _20016_);
  and (_20018_, _20000_, _19286_);
  or (_20019_, _20018_, _20017_);
  or (_20020_, _20019_, _19999_);
  not (_20021_, _19999_);
  or (_20022_, _20021_, _19282_);
  and (_20023_, _20022_, _20020_);
  or (_20024_, _20023_, _19998_);
  or (_20025_, _20011_, _19405_);
  and (_20026_, _20025_, _20010_);
  and (_20027_, _20026_, _20024_);
  or (_28215_[1], _20027_, _20015_);
  and (_20028_, _19294_, _19099_);
  and (_20029_, _20000_, word_in[2]);
  not (_20030_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_20031_, _20000_, _20030_);
  nor (_20032_, _20031_, _20029_);
  nor (_20033_, _20032_, _19999_);
  and (_20034_, _19999_, _19823_);
  or (_20035_, _20034_, _20033_);
  or (_20036_, _20035_, _19998_);
  or (_20037_, _20011_, _19417_);
  and (_20038_, _20037_, _20010_);
  and (_20039_, _20038_, _20036_);
  or (_28215_[2], _20039_, _20028_);
  and (_20040_, _19308_, _19099_);
  and (_20041_, _20000_, word_in[3]);
  not (_20042_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_20043_, _20000_, _20042_);
  nor (_20044_, _20043_, _20041_);
  nor (_20045_, _20044_, _19999_);
  and (_20046_, _19999_, _19836_);
  or (_20047_, _20046_, _20045_);
  or (_20048_, _20047_, _19998_);
  or (_20049_, _20011_, _19429_);
  and (_20050_, _20049_, _20010_);
  and (_20051_, _20050_, _20048_);
  or (_28215_[3], _20051_, _20040_);
  and (_20052_, _20000_, word_in[4]);
  not (_20053_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_20054_, _20000_, _20053_);
  nor (_20055_, _20054_, _20052_);
  nor (_20056_, _20055_, _19999_);
  and (_20057_, _19999_, _19849_);
  or (_20058_, _20057_, _20056_);
  and (_20059_, _20058_, _20011_);
  and (_20060_, _19998_, _19441_);
  or (_20061_, _20060_, _20059_);
  and (_20062_, _20061_, _20010_);
  and (_20063_, _20009_, word_in[28]);
  or (_28215_[4], _20063_, _20062_);
  and (_20064_, _20009_, word_in[29]);
  and (_20065_, _20000_, word_in[5]);
  not (_20066_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_20067_, _20000_, _20066_);
  nor (_20068_, _20067_, _20065_);
  nor (_20069_, _20068_, _19999_);
  and (_20070_, _19999_, _19864_);
  or (_20071_, _20070_, _20069_);
  or (_20072_, _20071_, _19998_);
  or (_20073_, _20011_, _19453_);
  and (_20074_, _20073_, _20010_);
  and (_20075_, _20074_, _20072_);
  or (_28215_[5], _20075_, _20064_);
  not (_20076_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_20077_, _20000_, _20076_);
  and (_20078_, _20000_, _19355_);
  or (_20079_, _20078_, _20077_);
  or (_20080_, _20079_, _19999_);
  or (_20081_, _20021_, _19876_);
  and (_20082_, _20081_, _20080_);
  or (_20083_, _20082_, _19998_);
  or (_20084_, _20011_, _19465_);
  and (_20085_, _20084_, _20083_);
  or (_20086_, _20085_, _20009_);
  or (_20087_, _20010_, word_in[30]);
  and (_28215_[6], _20087_, _20086_);
  and (_20088_, _20009_, word_in[31]);
  and (_20089_, _20000_, word_in[7]);
  nor (_20090_, _20000_, _18695_);
  nor (_20091_, _20090_, _20089_);
  nor (_20092_, _20091_, _19999_);
  and (_20093_, _19999_, _19074_);
  or (_20094_, _20093_, _20092_);
  or (_20095_, _20094_, _19998_);
  or (_20096_, _20011_, _19477_);
  and (_20097_, _20096_, _20010_);
  and (_20098_, _20097_, _20095_);
  or (_28215_[7], _20098_, _20088_);
  and (_20099_, _19051_, _18973_);
  and (_20100_, _20099_, _18690_);
  not (_20101_, _20100_);
  and (_20102_, _18689_, _18645_);
  or (_20103_, _20102_, _18701_);
  and (_20104_, _20103_, _19057_);
  and (_20105_, _20104_, _19258_);
  and (_20106_, _19062_, _18755_);
  and (_20107_, _19067_, _19163_);
  and (_20108_, _20107_, word_in[0]);
  not (_20109_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_20110_, _20107_, _20109_);
  nor (_20111_, _20110_, _20108_);
  nor (_20112_, _20111_, _20106_);
  and (_20113_, _20106_, word_in[8]);
  nor (_20114_, _20113_, _20112_);
  nor (_20115_, _20114_, _20105_);
  and (_20116_, _20105_, word_in[16]);
  or (_20117_, _20116_, _20115_);
  and (_20118_, _20117_, _20101_);
  and (_20119_, _20100_, _19252_);
  or (_28216_[0], _20119_, _20118_);
  not (_20120_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_20121_, _20107_, _20120_);
  and (_20122_, _20107_, _19286_);
  or (_20123_, _20122_, _20121_);
  or (_20124_, _20123_, _20106_);
  not (_20125_, _20106_);
  or (_20126_, _20125_, word_in[9]);
  and (_20127_, _20126_, _20124_);
  or (_20128_, _20127_, _20105_);
  not (_20129_, _20105_);
  or (_20130_, _20129_, word_in[17]);
  and (_20131_, _20130_, _20128_);
  or (_20132_, _20131_, _20100_);
  or (_20133_, _20101_, _19279_);
  and (_28216_[1], _20133_, _20132_);
  and (_20134_, _20107_, word_in[2]);
  not (_20135_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_20136_, _20107_, _20135_);
  nor (_20137_, _20136_, _20134_);
  nor (_20138_, _20137_, _20106_);
  and (_20139_, _20106_, word_in[10]);
  nor (_20140_, _20139_, _20138_);
  nor (_20141_, _20140_, _20105_);
  and (_20142_, _20105_, word_in[18]);
  or (_20143_, _20142_, _20141_);
  and (_20144_, _20143_, _20101_);
  and (_20145_, _20100_, _19294_);
  or (_28216_[2], _20145_, _20144_);
  and (_20146_, _20107_, word_in[3]);
  not (_20147_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_20148_, _20107_, _20147_);
  nor (_20149_, _20148_, _20146_);
  nor (_20150_, _20149_, _20106_);
  and (_20151_, _20106_, word_in[11]);
  nor (_20152_, _20151_, _20150_);
  nor (_20153_, _20152_, _20105_);
  and (_20154_, _20105_, word_in[19]);
  or (_20155_, _20154_, _20153_);
  and (_20156_, _20155_, _20101_);
  and (_20157_, _20100_, _19308_);
  or (_28216_[3], _20157_, _20156_);
  not (_20158_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_20159_, _20107_, _20158_);
  and (_20160_, _20107_, _19327_);
  or (_20161_, _20160_, _20159_);
  or (_20162_, _20161_, _20106_);
  or (_20163_, _20125_, word_in[12]);
  and (_20164_, _20163_, _20162_);
  or (_20165_, _20164_, _20105_);
  or (_20166_, _20129_, word_in[20]);
  and (_20167_, _20166_, _20165_);
  or (_20168_, _20167_, _20100_);
  or (_20169_, _20101_, _19322_);
  and (_28216_[4], _20169_, _20168_);
  not (_20170_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_20171_, _20107_, _20170_);
  and (_20172_, _20107_, _19339_);
  or (_20173_, _20172_, _20171_);
  or (_20174_, _20173_, _20106_);
  or (_20175_, _20125_, word_in[13]);
  and (_20176_, _20175_, _20174_);
  or (_20177_, _20176_, _20105_);
  or (_20178_, _20129_, word_in[21]);
  and (_20179_, _20178_, _20177_);
  or (_20180_, _20179_, _20100_);
  or (_20181_, _20101_, _19348_);
  and (_28216_[5], _20181_, _20180_);
  not (_20182_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_20183_, _20107_, _20182_);
  and (_20184_, _20107_, _19355_);
  or (_20185_, _20184_, _20183_);
  or (_20186_, _20185_, _20106_);
  or (_20187_, _20125_, word_in[14]);
  and (_20188_, _20187_, _20186_);
  or (_20189_, _20188_, _20105_);
  or (_20190_, _20129_, word_in[22]);
  and (_20191_, _20190_, _20189_);
  or (_20192_, _20191_, _20100_);
  or (_20193_, _20101_, _19350_);
  and (_28216_[6], _20193_, _20192_);
  and (_20194_, _20107_, word_in[7]);
  nor (_20195_, _20107_, _18836_);
  nor (_20196_, _20195_, _20194_);
  nor (_20197_, _20196_, _20106_);
  and (_20198_, _20106_, word_in[15]);
  nor (_20199_, _20198_, _20197_);
  nor (_20200_, _20199_, _20105_);
  and (_20201_, _20105_, word_in[23]);
  or (_20202_, _20201_, _20200_);
  and (_20203_, _20202_, _20101_);
  and (_20204_, _20100_, _19081_);
  or (_28216_[7], _20204_, _20203_);
  and (_20205_, _20104_, _19379_);
  and (_20206_, _19062_, _18768_);
  and (_20207_, _20206_, _18657_);
  and (_20208_, _19266_, _19169_);
  not (_20209_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_20210_, _19067_, _19169_);
  nor (_20211_, _20210_, _20209_);
  nor (_20212_, _20211_, _20208_);
  nor (_20213_, _20212_, _20207_);
  and (_20214_, _20207_, word_in[8]);
  nor (_20215_, _20214_, _20213_);
  nor (_20216_, _20215_, _20205_);
  and (_20217_, _20099_, _18679_);
  and (_20218_, _20205_, _19393_);
  or (_20219_, _20218_, _20217_);
  or (_20220_, _20219_, _20216_);
  not (_20221_, _20217_);
  or (_20222_, _20221_, _19252_);
  and (_28217_[0], _20222_, _20220_);
  not (_20223_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_20224_, _20210_, _20223_);
  and (_20225_, _19286_, _19169_);
  or (_20226_, _20225_, _20224_);
  or (_20227_, _20226_, _20207_);
  not (_20228_, _20207_);
  or (_20229_, _20228_, word_in[9]);
  and (_20230_, _20229_, _20227_);
  or (_20231_, _20230_, _20205_);
  not (_20232_, _20205_);
  or (_20233_, _20232_, _19405_);
  and (_20234_, _20233_, _20231_);
  or (_20235_, _20234_, _20217_);
  or (_20236_, _20221_, _19279_);
  and (_28217_[1], _20236_, _20235_);
  not (_20237_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_20238_, _20210_, _20237_);
  and (_20239_, _19299_, _19169_);
  or (_20240_, _20239_, _20238_);
  or (_20241_, _20240_, _20207_);
  or (_20242_, _20228_, word_in[10]);
  and (_20243_, _20242_, _20241_);
  or (_20244_, _20243_, _20205_);
  or (_20245_, _20232_, _19417_);
  and (_20246_, _20245_, _20244_);
  or (_20247_, _20246_, _20217_);
  or (_20248_, _20221_, _19294_);
  and (_28217_[2], _20248_, _20247_);
  not (_20249_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_20250_, _20210_, _20249_);
  and (_20251_, _19313_, _19169_);
  nor (_20252_, _20251_, _20250_);
  nor (_20253_, _20252_, _20207_);
  and (_20254_, _20207_, word_in[11]);
  nor (_20255_, _20254_, _20253_);
  nor (_20256_, _20255_, _20205_);
  and (_20257_, _20205_, _19429_);
  or (_20258_, _20257_, _20256_);
  and (_20259_, _20258_, _20221_);
  and (_20260_, _20217_, _19308_);
  or (_28217_[3], _20260_, _20259_);
  not (_20261_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_20262_, _20210_, _20261_);
  and (_20263_, _19327_, _19169_);
  or (_20264_, _20263_, _20262_);
  or (_20265_, _20264_, _20207_);
  or (_20266_, _20228_, word_in[12]);
  and (_20267_, _20266_, _20265_);
  or (_20268_, _20267_, _20205_);
  or (_20269_, _20232_, _19441_);
  and (_20270_, _20269_, _20268_);
  or (_20271_, _20270_, _20217_);
  or (_20272_, _20221_, _19322_);
  and (_28217_[4], _20272_, _20271_);
  not (_20273_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_20274_, _20210_, _20273_);
  and (_20275_, _20210_, _19339_);
  or (_20276_, _20275_, _20274_);
  or (_20277_, _20276_, _20207_);
  or (_20278_, _20228_, word_in[13]);
  and (_20279_, _20278_, _20277_);
  or (_20280_, _20279_, _20205_);
  or (_20281_, _20232_, _19453_);
  and (_20282_, _20281_, _20221_);
  and (_20283_, _20282_, _20280_);
  and (_20284_, _20217_, _19348_);
  or (_28217_[5], _20284_, _20283_);
  and (_20285_, _20210_, word_in[6]);
  not (_20286_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_20287_, _20210_, _20286_);
  nor (_20288_, _20287_, _20285_);
  nor (_20289_, _20288_, _20207_);
  and (_20290_, _20207_, word_in[14]);
  or (_20291_, _20290_, _20289_);
  or (_20292_, _20291_, _20205_);
  or (_20293_, _20232_, _19465_);
  and (_20294_, _20293_, _20221_);
  and (_20295_, _20294_, _20292_);
  and (_20296_, _20217_, _19350_);
  or (_28217_[6], _20296_, _20295_);
  and (_20297_, _20210_, word_in[7]);
  nor (_20298_, _20210_, _18728_);
  nor (_20299_, _20298_, _20297_);
  nor (_20300_, _20299_, _20207_);
  and (_20301_, _20207_, word_in[15]);
  nor (_20302_, _20301_, _20300_);
  nor (_20303_, _20302_, _20205_);
  and (_20304_, _20205_, _19477_);
  or (_20305_, _20304_, _20303_);
  and (_20306_, _20305_, _20221_);
  and (_20307_, _20217_, _19081_);
  or (_28217_[7], _20307_, _20306_);
  and (_20308_, _19051_, _18753_);
  not (_20309_, _20308_);
  and (_20310_, _20104_, _19486_);
  and (_20311_, _20206_, _18690_);
  not (_20312_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_20313_, _19067_, _19180_);
  nor (_20314_, _20313_, _20312_);
  and (_20315_, _20313_, _19266_);
  nor (_20316_, _20315_, _20314_);
  nor (_20317_, _20316_, _20311_);
  and (_20318_, _20311_, word_in[8]);
  nor (_20319_, _20318_, _20317_);
  nor (_20320_, _20319_, _20310_);
  and (_20321_, _20310_, _19393_);
  or (_20322_, _20321_, _20320_);
  and (_20323_, _20322_, _20309_);
  and (_20324_, _20308_, _19252_);
  or (_28203_[0], _20324_, _20323_);
  not (_20325_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_20326_, _20313_, _20325_);
  and (_20327_, _20313_, _19286_);
  or (_20328_, _20327_, _20326_);
  or (_20329_, _20328_, _20311_);
  not (_20330_, _20311_);
  or (_20331_, _20330_, word_in[9]);
  and (_20332_, _20331_, _20329_);
  or (_20333_, _20332_, _20310_);
  not (_20334_, _20310_);
  or (_20335_, _20334_, _19405_);
  and (_20336_, _20335_, _20309_);
  and (_20337_, _20336_, _20333_);
  and (_20338_, _20308_, _19279_);
  or (_28203_[1], _20338_, _20337_);
  not (_20339_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_20340_, _20313_, _20339_);
  and (_20341_, _20313_, _19299_);
  or (_20342_, _20341_, _20340_);
  or (_20343_, _20342_, _20311_);
  or (_20344_, _20330_, word_in[10]);
  and (_20345_, _20344_, _20343_);
  or (_20346_, _20345_, _20310_);
  or (_20347_, _20334_, _19417_);
  and (_20348_, _20347_, _20309_);
  and (_20349_, _20348_, _20346_);
  and (_20350_, _20308_, _19294_);
  or (_28203_[2], _20350_, _20349_);
  and (_20351_, _20310_, _19429_);
  and (_20352_, _20313_, word_in[3]);
  not (_20353_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_20354_, _20313_, _20353_);
  nor (_20355_, _20354_, _20352_);
  nor (_20356_, _20355_, _20311_);
  and (_20357_, _20311_, word_in[11]);
  nor (_20358_, _20357_, _20356_);
  nor (_20359_, _20358_, _20310_);
  or (_20360_, _20359_, _20351_);
  and (_20361_, _20360_, _20309_);
  and (_20362_, _20308_, _19308_);
  or (_28203_[3], _20362_, _20361_);
  not (_20363_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_20364_, _20313_, _20363_);
  and (_20365_, _20313_, _19327_);
  or (_20366_, _20365_, _20364_);
  or (_20367_, _20366_, _20311_);
  or (_20368_, _20330_, word_in[12]);
  nand (_20369_, _20368_, _20367_);
  nor (_20370_, _20369_, _20310_);
  and (_20371_, _20310_, _19441_);
  or (_20372_, _20371_, _20308_);
  or (_20373_, _20372_, _20370_);
  or (_20374_, _20309_, _19322_);
  and (_28203_[4], _20374_, _20373_);
  not (_20375_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_20376_, _20313_, _20375_);
  and (_20377_, _20313_, _19339_);
  or (_20378_, _20377_, _20376_);
  or (_20379_, _20378_, _20311_);
  or (_20380_, _20330_, word_in[13]);
  and (_20381_, _20380_, _20379_);
  or (_20382_, _20381_, _20310_);
  or (_20383_, _20334_, _19453_);
  and (_20384_, _20383_, _20309_);
  and (_20385_, _20384_, _20382_);
  and (_20386_, _20308_, _19348_);
  or (_28203_[5], _20386_, _20385_);
  and (_20387_, _20313_, word_in[6]);
  not (_20388_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_20389_, _20313_, _20388_);
  nor (_20390_, _20389_, _20387_);
  nor (_20391_, _20390_, _20311_);
  and (_20392_, _20311_, word_in[14]);
  or (_20393_, _20392_, _20391_);
  or (_20394_, _20393_, _20310_);
  or (_20395_, _20334_, _19465_);
  and (_20396_, _20395_, _20309_);
  and (_20397_, _20396_, _20394_);
  and (_20398_, _20308_, _19350_);
  or (_28203_[6], _20398_, _20397_);
  nor (_20399_, _20313_, _18841_);
  and (_20400_, _20313_, _19068_);
  or (_20401_, _20400_, _20399_);
  or (_20402_, _20401_, _20311_);
  or (_20403_, _20330_, word_in[15]);
  and (_20404_, _20403_, _20402_);
  or (_20405_, _20404_, _20310_);
  or (_20406_, _20334_, _19477_);
  and (_20407_, _20406_, _20309_);
  and (_20408_, _20407_, _20405_);
  and (_20409_, _20308_, _19081_);
  or (_28203_[7], _20409_, _20408_);
  and (_20410_, _20104_, _19056_);
  and (_20411_, _20206_, _18679_);
  not (_20412_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_20413_, _19067_, _19205_);
  nor (_20414_, _20413_, _20412_);
  and (_20415_, _20413_, _19266_);
  or (_20416_, _20415_, _20414_);
  or (_20417_, _20416_, _20411_);
  not (_20418_, _20411_);
  or (_20419_, _20418_, word_in[8]);
  and (_20420_, _20419_, _20417_);
  or (_20421_, _20420_, _20410_);
  and (_20422_, _19050_, _19163_);
  not (_20423_, _20422_);
  not (_20424_, _20410_);
  or (_20425_, _20424_, word_in[16]);
  and (_20426_, _20425_, _20423_);
  and (_20427_, _20426_, _20421_);
  and (_20428_, _20422_, word_in[24]);
  or (_28204_[0], _20428_, _20427_);
  not (_20429_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_20430_, _20413_, _20429_);
  and (_20431_, _20413_, _19286_);
  or (_20432_, _20431_, _20430_);
  or (_20433_, _20432_, _20411_);
  or (_20434_, _20418_, word_in[9]);
  and (_20435_, _20434_, _20433_);
  or (_20436_, _20435_, _20410_);
  or (_20437_, _20424_, word_in[17]);
  and (_20438_, _20437_, _20423_);
  and (_20439_, _20438_, _20436_);
  and (_20440_, _20422_, word_in[25]);
  or (_28204_[1], _20440_, _20439_);
  and (_20441_, _20413_, word_in[2]);
  not (_20442_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_20443_, _20413_, _20442_);
  nor (_20444_, _20443_, _20441_);
  nor (_20445_, _20444_, _20411_);
  and (_20446_, _20411_, word_in[10]);
  nor (_20447_, _20446_, _20445_);
  nor (_20448_, _20447_, _20410_);
  and (_20449_, _20410_, word_in[18]);
  or (_20450_, _20449_, _20448_);
  and (_20451_, _20450_, _20423_);
  and (_20452_, _20422_, word_in[26]);
  or (_28204_[2], _20452_, _20451_);
  not (_20453_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_20454_, _20413_, _20453_);
  and (_20455_, _20413_, _19313_);
  or (_20456_, _20455_, _20454_);
  or (_20457_, _20456_, _20411_);
  or (_20458_, _20418_, word_in[11]);
  and (_20459_, _20458_, _20457_);
  or (_20460_, _20459_, _20410_);
  or (_20461_, _20424_, word_in[19]);
  and (_20462_, _20461_, _20423_);
  and (_20463_, _20462_, _20460_);
  and (_20464_, _20422_, word_in[27]);
  or (_28204_[3], _20464_, _20463_);
  not (_20465_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_20466_, _20413_, _20465_);
  and (_20467_, _20413_, _19327_);
  or (_20468_, _20467_, _20466_);
  or (_20469_, _20468_, _20411_);
  or (_20470_, _20418_, word_in[12]);
  and (_20471_, _20470_, _20469_);
  or (_20472_, _20471_, _20410_);
  or (_20473_, _20424_, word_in[20]);
  and (_20474_, _20473_, _20423_);
  and (_20475_, _20474_, _20472_);
  and (_20476_, _20422_, word_in[28]);
  or (_28204_[4], _20476_, _20475_);
  not (_20477_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_20478_, _20413_, _20477_);
  and (_20479_, _20413_, _19339_);
  or (_20480_, _20479_, _20478_);
  or (_20481_, _20480_, _20411_);
  or (_20482_, _20418_, word_in[13]);
  and (_20483_, _20482_, _20481_);
  or (_20484_, _20483_, _20410_);
  or (_20485_, _20424_, _19453_);
  and (_20486_, _20485_, _20423_);
  and (_20487_, _20486_, _20484_);
  and (_20488_, _20422_, word_in[29]);
  or (_28204_[5], _20488_, _20487_);
  and (_20489_, _20413_, word_in[6]);
  not (_20490_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_20491_, _20413_, _20490_);
  nor (_20492_, _20491_, _20489_);
  nor (_20493_, _20492_, _20411_);
  and (_20494_, _20411_, word_in[14]);
  nor (_20495_, _20494_, _20493_);
  nor (_20496_, _20495_, _20410_);
  and (_20497_, _20410_, word_in[22]);
  or (_20498_, _20497_, _20496_);
  and (_20499_, _20498_, _20423_);
  and (_20500_, _20422_, word_in[30]);
  or (_28204_[6], _20500_, _20499_);
  nor (_20501_, _20413_, _18723_);
  and (_20502_, _20413_, _19068_);
  or (_20503_, _20502_, _20501_);
  or (_20504_, _20503_, _20411_);
  or (_20505_, _20418_, word_in[15]);
  and (_20506_, _20505_, _20504_);
  or (_20507_, _20506_, _20410_);
  or (_20508_, _20424_, word_in[23]);
  and (_20509_, _20508_, _20423_);
  and (_20510_, _20509_, _20507_);
  and (_20511_, _20422_, word_in[31]);
  or (_28204_[7], _20511_, _20510_);
  and (_20512_, _19052_, _18690_);
  and (_20513_, _19258_, _19059_);
  and (_20514_, _19062_, _19205_);
  and (_20515_, _18657_, _18647_);
  and (_20516_, _19067_, _20515_);
  and (_20517_, _20516_, _19266_);
  not (_20518_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_20519_, _20516_, _20518_);
  or (_20520_, _20519_, _20517_);
  or (_20521_, _20520_, _20514_);
  not (_20522_, _20514_);
  or (_20523_, _20522_, word_in[8]);
  and (_20524_, _20523_, _20521_);
  or (_20525_, _20524_, _20513_);
  not (_20526_, _20513_);
  or (_20527_, _20526_, word_in[16]);
  and (_20528_, _20527_, _20525_);
  or (_20529_, _20528_, _20512_);
  not (_20530_, _20512_);
  or (_20531_, _20530_, _19252_);
  and (_28205_[0], _20531_, _20529_);
  not (_20532_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_20533_, _20516_, _20532_);
  and (_20534_, _20516_, _19286_);
  nor (_20535_, _20534_, _20533_);
  nor (_20536_, _20535_, _20514_);
  and (_20537_, _20514_, word_in[9]);
  nor (_20538_, _20537_, _20536_);
  nor (_20539_, _20538_, _20513_);
  and (_20540_, _20513_, word_in[17]);
  or (_20541_, _20540_, _20539_);
  and (_20542_, _20541_, _20530_);
  and (_20543_, _20512_, _19279_);
  or (_28205_[1], _20543_, _20542_);
  not (_20544_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_20545_, _20516_, _20544_);
  and (_20546_, _20516_, _19299_);
  or (_20547_, _20546_, _20545_);
  or (_20548_, _20547_, _20514_);
  or (_20549_, _20522_, word_in[10]);
  and (_20550_, _20549_, _20548_);
  or (_20551_, _20550_, _20513_);
  or (_20552_, _20526_, word_in[18]);
  and (_20553_, _20552_, _20551_);
  or (_20554_, _20553_, _20512_);
  or (_20555_, _20530_, _19294_);
  and (_28205_[2], _20555_, _20554_);
  and (_20556_, _20516_, word_in[3]);
  not (_20557_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_20558_, _20516_, _20557_);
  nor (_20559_, _20558_, _20556_);
  nor (_20560_, _20559_, _20514_);
  and (_20561_, _20514_, word_in[11]);
  nor (_20562_, _20561_, _20560_);
  nor (_20563_, _20562_, _20513_);
  and (_20564_, _20513_, word_in[19]);
  or (_20565_, _20564_, _20563_);
  and (_20566_, _20565_, _20530_);
  and (_20567_, _20512_, _19308_);
  or (_28205_[3], _20567_, _20566_);
  not (_20568_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_20569_, _20516_, _20568_);
  and (_20570_, _20516_, _19327_);
  or (_20571_, _20570_, _20569_);
  or (_20572_, _20571_, _20514_);
  or (_20573_, _20522_, word_in[12]);
  and (_20574_, _20573_, _20572_);
  or (_20575_, _20574_, _20513_);
  or (_20576_, _20526_, word_in[20]);
  and (_20577_, _20576_, _20575_);
  or (_20578_, _20577_, _20512_);
  or (_20579_, _20530_, _19322_);
  and (_28205_[4], _20579_, _20578_);
  not (_20580_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_20581_, _20516_, _20580_);
  and (_20582_, _20516_, word_in[5]);
  nor (_20583_, _20582_, _20581_);
  nor (_20584_, _20583_, _20514_);
  and (_20585_, _20514_, word_in[13]);
  nor (_20586_, _20585_, _20584_);
  nor (_20587_, _20586_, _20513_);
  and (_20588_, _20513_, word_in[21]);
  or (_20589_, _20588_, _20587_);
  and (_20590_, _20589_, _20530_);
  and (_20591_, _20512_, _19348_);
  or (_28205_[5], _20591_, _20590_);
  and (_20592_, _20516_, word_in[6]);
  not (_20593_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_20594_, _20516_, _20593_);
  nor (_20595_, _20594_, _20592_);
  nor (_20596_, _20595_, _20514_);
  and (_20597_, _20514_, word_in[14]);
  nor (_20598_, _20597_, _20596_);
  nor (_20599_, _20598_, _20513_);
  and (_20600_, _20513_, word_in[22]);
  or (_20601_, _20600_, _20599_);
  and (_20602_, _20601_, _20530_);
  and (_20603_, _20512_, _19350_);
  or (_28205_[6], _20603_, _20602_);
  nor (_20604_, _20516_, _18848_);
  and (_20605_, _20516_, _19068_);
  or (_20606_, _20605_, _20604_);
  or (_20607_, _20606_, _20514_);
  or (_20608_, _20522_, word_in[15]);
  and (_20609_, _20608_, _20607_);
  or (_20610_, _20609_, _20513_);
  or (_20611_, _20526_, word_in[23]);
  and (_20612_, _20611_, _20610_);
  or (_20613_, _20612_, _20512_);
  or (_20614_, _20530_, _19081_);
  and (_28205_[7], _20614_, _20613_);
  and (_20615_, _19052_, _18679_);
  not (_20616_, _20615_);
  and (_20617_, _19379_, _19059_);
  not (_20618_, _20617_);
  and (_20619_, _19064_, _18657_);
  not (_20620_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_20621_, _19067_, _19233_);
  nor (_20622_, _20621_, _20620_);
  and (_20623_, _19266_, _19233_);
  nor (_20624_, _20623_, _20622_);
  nor (_20625_, _20624_, _20619_);
  and (_20626_, _20619_, _19796_);
  or (_20627_, _20626_, _20625_);
  and (_20628_, _20627_, _20618_);
  and (_20629_, _20617_, _19393_);
  or (_20630_, _20629_, _20628_);
  and (_20631_, _20630_, _20616_);
  and (_20632_, _20615_, _19252_);
  or (_28206_[0], _20632_, _20631_);
  not (_20633_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_20634_, _20621_, _20633_);
  and (_20635_, _19286_, _19233_);
  nor (_20636_, _20635_, _20634_);
  nor (_20637_, _20636_, _20619_);
  and (_20638_, _20619_, _19282_);
  or (_20639_, _20638_, _20637_);
  or (_20640_, _20639_, _20617_);
  or (_20641_, _20618_, _19405_);
  and (_20642_, _20641_, _20616_);
  and (_20643_, _20642_, _20640_);
  and (_20644_, _20615_, _19279_);
  or (_28206_[1], _20644_, _20643_);
  not (_20645_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_20646_, _20621_, _20645_);
  and (_20647_, _20621_, _19299_);
  or (_20648_, _20647_, _20646_);
  or (_20649_, _20648_, _20619_);
  not (_20650_, _20619_);
  or (_20651_, _20650_, _19823_);
  and (_20652_, _20651_, _20649_);
  or (_20653_, _20652_, _20617_);
  or (_20654_, _20618_, _19417_);
  and (_20655_, _20654_, _20616_);
  and (_20656_, _20655_, _20653_);
  and (_20657_, _20615_, _19294_);
  or (_28206_[2], _20657_, _20656_);
  and (_20658_, _20621_, word_in[3]);
  not (_20659_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_20660_, _20621_, _20659_);
  nor (_20661_, _20660_, _20658_);
  nor (_20662_, _20661_, _20619_);
  and (_20663_, _20619_, _19836_);
  or (_20664_, _20663_, _20662_);
  and (_20665_, _20664_, _20618_);
  and (_20666_, _20617_, _19429_);
  or (_20667_, _20666_, _20615_);
  or (_20668_, _20667_, _20665_);
  or (_20669_, _20616_, _19308_);
  and (_28206_[3], _20669_, _20668_);
  not (_20670_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_20671_, _20621_, _20670_);
  and (_20672_, _19327_, _19233_);
  nor (_20673_, _20672_, _20671_);
  nor (_20674_, _20673_, _20619_);
  and (_20675_, _20619_, _19849_);
  or (_20676_, _20675_, _20674_);
  and (_20677_, _20676_, _20618_);
  and (_20678_, _20617_, _19441_);
  or (_20679_, _20678_, _20677_);
  and (_20680_, _20679_, _20616_);
  and (_20681_, _20615_, _19322_);
  or (_28206_[4], _20681_, _20680_);
  not (_20682_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_20683_, _20621_, _20682_);
  and (_20684_, _20621_, _19339_);
  or (_20685_, _20684_, _20683_);
  or (_20686_, _20685_, _20619_);
  or (_20687_, _20650_, _19864_);
  and (_20688_, _20687_, _20686_);
  or (_20689_, _20688_, _20617_);
  or (_20690_, _20618_, _19453_);
  and (_20691_, _20690_, _20616_);
  and (_20692_, _20691_, _20689_);
  and (_20693_, _20615_, _19348_);
  or (_28206_[5], _20693_, _20692_);
  not (_20694_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_20695_, _20621_, _20694_);
  and (_20696_, _20621_, _19355_);
  or (_20697_, _20696_, _20695_);
  or (_20698_, _20697_, _20619_);
  or (_20699_, _20650_, _19876_);
  and (_20700_, _20699_, _20698_);
  or (_20701_, _20700_, _20617_);
  or (_20702_, _20618_, _19465_);
  and (_20703_, _20702_, _20701_);
  or (_20704_, _20703_, _20615_);
  or (_20705_, _20616_, _19350_);
  and (_28206_[6], _20705_, _20704_);
  nor (_20706_, _20621_, _18711_);
  and (_20707_, _20621_, _19068_);
  or (_20708_, _20707_, _20706_);
  or (_20709_, _20708_, _20619_);
  or (_20710_, _20650_, _19074_);
  and (_20711_, _20710_, _20709_);
  or (_20712_, _20711_, _20617_);
  or (_20713_, _20618_, _19477_);
  and (_20714_, _20713_, _20616_);
  and (_20715_, _20714_, _20712_);
  and (_20716_, _20615_, _19081_);
  or (_28206_[7], _20716_, _20715_);
  and (_20717_, _19486_, _19058_);
  and (_20718_, _19064_, _18690_);
  not (_20719_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_20720_, _19067_, _19087_);
  nor (_20721_, _20720_, _20719_);
  and (_20722_, _20720_, _19266_);
  nor (_20723_, _20722_, _20721_);
  nor (_20724_, _20723_, _20718_);
  and (_20725_, _20718_, _19796_);
  nor (_20726_, _20725_, _20724_);
  nor (_20727_, _20726_, _20717_);
  and (_20728_, _19052_, _18667_);
  and (_20729_, _20717_, _19393_);
  or (_20730_, _20729_, _20728_);
  or (_20731_, _20730_, _20727_);
  not (_20732_, _20728_);
  or (_20733_, _20732_, _19252_);
  and (_28207_[0], _20733_, _20731_);
  not (_20734_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_20735_, _20720_, _20734_);
  and (_20736_, _20720_, _19286_);
  or (_20737_, _20736_, _20735_);
  or (_20738_, _20737_, _20718_);
  not (_20739_, _20718_);
  or (_20740_, _20739_, _19282_);
  and (_20741_, _20740_, _20738_);
  or (_20742_, _20741_, _20717_);
  not (_20743_, _20717_);
  or (_20744_, _20743_, _19405_);
  and (_20745_, _20744_, _20732_);
  and (_20746_, _20745_, _20742_);
  and (_20747_, _20728_, _19279_);
  or (_28207_[1], _20747_, _20746_);
  not (_20748_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_20749_, _20720_, _20748_);
  and (_20750_, _20720_, _19299_);
  or (_20751_, _20750_, _20749_);
  or (_20752_, _20751_, _20718_);
  or (_20753_, _20739_, _19823_);
  and (_20754_, _20753_, _20752_);
  or (_20755_, _20754_, _20717_);
  or (_20756_, _20743_, _19417_);
  and (_20757_, _20756_, _20755_);
  or (_20758_, _20757_, _20728_);
  or (_20759_, _20732_, _19294_);
  and (_28207_[2], _20759_, _20758_);
  not (_20760_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_20761_, _20720_, _20760_);
  and (_20762_, _20720_, _19313_);
  or (_20763_, _20762_, _20761_);
  or (_20764_, _20763_, _20718_);
  or (_20765_, _20739_, _19836_);
  and (_20766_, _20765_, _20764_);
  or (_20767_, _20766_, _20717_);
  or (_20768_, _20743_, _19429_);
  and (_20769_, _20768_, _20767_);
  or (_20770_, _20769_, _20728_);
  or (_20771_, _20732_, _19308_);
  and (_28207_[3], _20771_, _20770_);
  not (_20772_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_20773_, _20720_, _20772_);
  and (_20774_, _20720_, _19327_);
  or (_20775_, _20774_, _20773_);
  or (_20776_, _20775_, _20718_);
  or (_20777_, _20739_, _19849_);
  and (_20778_, _20777_, _20776_);
  or (_20779_, _20778_, _20717_);
  or (_20780_, _20743_, _19441_);
  and (_20781_, _20780_, _20779_);
  or (_20782_, _20781_, _20728_);
  or (_20783_, _20732_, _19322_);
  and (_28207_[4], _20783_, _20782_);
  and (_20784_, _20720_, word_in[5]);
  not (_20785_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_20786_, _20720_, _20785_);
  nor (_20787_, _20786_, _20784_);
  nor (_20788_, _20787_, _20718_);
  and (_20789_, _20718_, _19864_);
  or (_20790_, _20789_, _20788_);
  or (_20791_, _20790_, _20717_);
  or (_20792_, _20743_, _19453_);
  and (_20793_, _20792_, _20732_);
  and (_20794_, _20793_, _20791_);
  and (_20795_, _20728_, _19348_);
  or (_28207_[5], _20795_, _20794_);
  not (_20796_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_20797_, _20720_, _20796_);
  and (_20798_, _20720_, _19355_);
  or (_20799_, _20798_, _20797_);
  or (_20800_, _20799_, _20718_);
  or (_20801_, _20739_, _19876_);
  and (_20802_, _20801_, _20800_);
  or (_20803_, _20802_, _20717_);
  or (_20804_, _20743_, _19465_);
  and (_20805_, _20804_, _20803_);
  or (_20806_, _20805_, _20728_);
  or (_20807_, _20732_, _19350_);
  and (_28207_[6], _20807_, _20806_);
  nor (_20808_, _20720_, _18853_);
  and (_20809_, _20720_, _19068_);
  or (_20810_, _20809_, _20808_);
  or (_20811_, _20810_, _20718_);
  or (_20812_, _20739_, _19074_);
  and (_20813_, _20812_, _20811_);
  or (_20814_, _20813_, _20717_);
  or (_20815_, _20743_, _19477_);
  and (_20816_, _20815_, _20732_);
  and (_20817_, _20816_, _20814_);
  and (_20818_, _20728_, _19081_);
  or (_28207_[7], _20818_, _20817_);
  and (_20819_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_20820_, _19266_, _19066_);
  nor (_20821_, _20820_, _20819_);
  nor (_20822_, _20821_, _19065_);
  and (_20823_, _19796_, _19065_);
  or (_20824_, _20823_, _20822_);
  and (_20825_, _20824_, _19061_);
  and (_20826_, _19060_, word_in[16]);
  or (_20827_, _20826_, _20825_);
  and (_20828_, _20827_, _19054_);
  and (_20829_, _19252_, _19053_);
  or (_28208_[0], _20829_, _20828_);
  and (_20830_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_20831_, _19286_, _19066_);
  nor (_20832_, _20831_, _20830_);
  nor (_20833_, _20832_, _19065_);
  and (_20834_, _19282_, _19065_);
  or (_20835_, _20834_, _20833_);
  and (_20836_, _20835_, _19061_);
  and (_20837_, _19060_, word_in[17]);
  or (_20838_, _20837_, _20836_);
  and (_20839_, _20838_, _19054_);
  and (_20840_, _19279_, _19053_);
  or (_28208_[1], _20840_, _20839_);
  and (_20841_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_20842_, _19299_, _19066_);
  nor (_20843_, _20842_, _20841_);
  nor (_20844_, _20843_, _19065_);
  and (_20845_, _19823_, _19065_);
  or (_20846_, _20845_, _20844_);
  and (_20847_, _20846_, _19061_);
  and (_20848_, _19060_, word_in[18]);
  or (_20849_, _20848_, _20847_);
  and (_20850_, _20849_, _19054_);
  and (_20851_, _19294_, _19053_);
  or (_28208_[2], _20851_, _20850_);
  and (_20852_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_20853_, _19313_, _19066_);
  nor (_20854_, _20853_, _20852_);
  nor (_20855_, _20854_, _19065_);
  and (_20856_, _19836_, _19065_);
  or (_20857_, _20856_, _20855_);
  and (_20858_, _20857_, _19061_);
  and (_20859_, _19060_, word_in[19]);
  or (_20860_, _20859_, _20858_);
  and (_20861_, _20860_, _19054_);
  and (_20862_, _19308_, _19053_);
  or (_28208_[3], _20862_, _20861_);
  and (_20863_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_20864_, _19327_, _19066_);
  nor (_20865_, _20864_, _20863_);
  nor (_20866_, _20865_, _19065_);
  and (_20867_, _19849_, _19065_);
  or (_20868_, _20867_, _20866_);
  and (_20869_, _20868_, _19061_);
  and (_20870_, _19060_, word_in[20]);
  or (_20871_, _20870_, _20869_);
  and (_20872_, _20871_, _19054_);
  and (_20873_, _19322_, _19053_);
  or (_28208_[4], _20873_, _20872_);
  and (_20874_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_20875_, _19339_, _19066_);
  nor (_20876_, _20875_, _20874_);
  nor (_20877_, _20876_, _19065_);
  and (_20878_, _19864_, _19065_);
  or (_20879_, _20878_, _20877_);
  and (_20880_, _20879_, _19061_);
  and (_20881_, _19060_, word_in[21]);
  or (_20882_, _20881_, _20880_);
  and (_20883_, _20882_, _19054_);
  and (_20884_, _19348_, _19053_);
  or (_28208_[5], _20884_, _20883_);
  and (_20885_, _19070_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_20886_, _19355_, _19066_);
  nor (_20887_, _20886_, _20885_);
  nor (_20888_, _20887_, _19065_);
  and (_20889_, _19876_, _19065_);
  or (_20890_, _20889_, _20888_);
  and (_20891_, _20890_, _19061_);
  and (_20892_, _19060_, word_in[22]);
  or (_20893_, _20892_, _20891_);
  and (_20894_, _20893_, _19054_);
  and (_20895_, _19350_, _19053_);
  or (_28208_[6], _20895_, _20894_);
  and (_20896_, _18694_, word_in[0]);
  nand (_20897_, _18653_, _20412_);
  or (_20898_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_20899_, _20898_, _20897_);
  and (_20900_, _20899_, _18873_);
  nand (_20901_, _18653_, _20620_);
  or (_20902_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_20903_, _20902_, _20901_);
  and (_20904_, _20903_, _18710_);
  nor (_20905_, _18656_, _18635_);
  nand (_20906_, _18653_, _20209_);
  or (_20907_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_20908_, _20907_, _20906_);
  and (_20909_, _20908_, _20905_);
  or (_20910_, _20909_, _20904_);
  or (_20911_, _20910_, _20900_);
  and (_20912_, _20911_, _18639_);
  nand (_20913_, _18653_, _19790_);
  or (_20914_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_20915_, _20914_, _20913_);
  and (_20916_, _20915_, _18710_);
  not (_20917_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand (_20918_, _18653_, _20917_);
  or (_20919_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_20920_, _20919_, _20918_);
  and (_20921_, _20920_, _20905_);
  or (_20922_, _20921_, _20916_);
  nand (_20923_, _18653_, _20002_);
  or (_20924_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_20925_, _20924_, _20923_);
  and (_20926_, _20925_, _18700_);
  not (_20927_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand (_20928_, _18653_, _20927_);
  or (_20929_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_20930_, _20929_, _20928_);
  and (_20931_, _20930_, _18873_);
  or (_20932_, _20931_, _20926_);
  or (_20933_, _20932_, _20922_);
  and (_20934_, _20933_, _18699_);
  not (_20935_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nand (_20936_, _18653_, _20935_);
  or (_20937_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_20938_, _20937_, _20936_);
  and (_20939_, _20938_, _18707_);
  or (_20940_, _20939_, _20934_);
  nor (_20941_, _20940_, _20912_);
  nor (_20942_, _20941_, _18694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _20942_, _20896_);
  and (_20943_, _18694_, word_in[1]);
  nand (_20944_, _18653_, _20223_);
  or (_20945_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_20946_, _20945_, _20944_);
  and (_20947_, _20946_, _20905_);
  nand (_20948_, _18653_, _20429_);
  or (_20949_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_20950_, _20949_, _20948_);
  and (_20951_, _20950_, _18873_);
  or (_20952_, _20951_, _20947_);
  nand (_20953_, _18653_, _20633_);
  or (_20954_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_20955_, _20954_, _20953_);
  and (_20956_, _20955_, _18710_);
  or (_20957_, _20956_, _20952_);
  and (_20958_, _20957_, _18639_);
  nand (_20959_, _18653_, _19806_);
  or (_20960_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_20961_, _20960_, _20959_);
  and (_20962_, _20961_, _18710_);
  not (_20963_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand (_20964_, _18653_, _20963_);
  or (_20965_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_20966_, _20965_, _20964_);
  and (_20967_, _20966_, _18873_);
  or (_20968_, _20967_, _20962_);
  nand (_20969_, _18653_, _20016_);
  or (_20970_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_20971_, _20970_, _20969_);
  and (_20972_, _20971_, _18700_);
  not (_20973_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nand (_20974_, _18653_, _20973_);
  or (_20975_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_20976_, _20975_, _20974_);
  and (_20977_, _20976_, _20905_);
  or (_20978_, _20977_, _20972_);
  or (_20979_, _20978_, _20968_);
  and (_20980_, _20979_, _18699_);
  not (_20981_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nand (_20982_, _18653_, _20981_);
  or (_20983_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_20984_, _20983_, _20982_);
  and (_20985_, _20984_, _18707_);
  or (_20986_, _20985_, _20980_);
  nor (_20987_, _20986_, _20958_);
  nor (_20988_, _20987_, _18694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _20988_, _20943_);
  and (_20989_, _18694_, word_in[2]);
  nand (_20990_, _18653_, _20442_);
  or (_20991_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_20992_, _20991_, _20990_);
  and (_20993_, _20992_, _18873_);
  nand (_20994_, _18653_, _20645_);
  or (_20995_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_20996_, _20995_, _20994_);
  and (_20997_, _20996_, _18710_);
  nand (_20998_, _18653_, _20237_);
  or (_20999_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_21000_, _20999_, _20998_);
  and (_21001_, _21000_, _20905_);
  or (_21002_, _21001_, _20997_);
  or (_21003_, _21002_, _20993_);
  and (_21004_, _21003_, _18639_);
  nand (_21005_, _18653_, _19818_);
  or (_21006_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_21007_, _21006_, _21005_);
  and (_21008_, _21007_, _18710_);
  not (_21009_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_21010_, _18653_, _21009_);
  or (_21011_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_21012_, _21011_, _21010_);
  and (_21013_, _21012_, _20905_);
  or (_21014_, _21013_, _21008_);
  nand (_21015_, _18653_, _20030_);
  or (_21016_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_21017_, _21016_, _21015_);
  and (_21018_, _21017_, _18700_);
  not (_21019_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand (_21020_, _18653_, _21019_);
  or (_21021_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_21022_, _21021_, _21020_);
  and (_21023_, _21022_, _18873_);
  or (_21024_, _21023_, _21018_);
  or (_21025_, _21024_, _21014_);
  and (_21026_, _21025_, _18699_);
  not (_21027_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nand (_21028_, _18653_, _21027_);
  or (_21029_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_21030_, _21029_, _21028_);
  and (_21031_, _21030_, _18707_);
  or (_21032_, _21031_, _21026_);
  nor (_21033_, _21032_, _21004_);
  nor (_21034_, _21033_, _18694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _21034_, _20989_);
  and (_21035_, _18694_, word_in[3]);
  nand (_21036_, _18653_, _19831_);
  or (_21037_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_21038_, _21037_, _21036_);
  and (_21039_, _21038_, _18710_);
  not (_21040_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nand (_21041_, _18653_, _21040_);
  or (_21042_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_21043_, _21042_, _21041_);
  and (_21044_, _21043_, _18873_);
  or (_21045_, _21044_, _21039_);
  nand (_21046_, _18653_, _20042_);
  or (_21047_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_21048_, _21047_, _21046_);
  and (_21049_, _21048_, _18700_);
  not (_21050_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nand (_21051_, _18653_, _21050_);
  or (_21052_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_21053_, _21052_, _21051_);
  and (_21054_, _21053_, _20905_);
  or (_21055_, _21054_, _21049_);
  or (_21056_, _21055_, _21045_);
  and (_21057_, _21056_, _18699_);
  nand (_21058_, _18653_, _20249_);
  or (_21059_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_21060_, _21059_, _21058_);
  and (_21061_, _21060_, _20905_);
  nand (_21062_, _18653_, _20453_);
  or (_21063_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_21064_, _21063_, _21062_);
  and (_21065_, _21064_, _18873_);
  or (_21066_, _21065_, _21061_);
  nand (_21067_, _18653_, _20659_);
  or (_21068_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_21069_, _21068_, _21067_);
  and (_21070_, _21069_, _18710_);
  or (_21071_, _21070_, _21066_);
  and (_21072_, _21071_, _18639_);
  not (_21073_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nand (_21074_, _18653_, _21073_);
  or (_21075_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_21076_, _21075_, _21074_);
  and (_21077_, _21076_, _18707_);
  or (_21078_, _21077_, _21072_);
  nor (_21079_, _21078_, _21057_);
  nor (_21080_, _21079_, _18694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _21080_, _21035_);
  and (_21081_, _18694_, word_in[4]);
  nand (_21082_, _18653_, _19844_);
  or (_21083_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_21084_, _21083_, _21082_);
  and (_21085_, _21084_, _18710_);
  not (_21086_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand (_21087_, _18653_, _21086_);
  or (_21088_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_21089_, _21088_, _21087_);
  and (_21090_, _21089_, _20905_);
  or (_21091_, _21090_, _21085_);
  nand (_21092_, _18653_, _20053_);
  or (_21093_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_21094_, _21093_, _21092_);
  and (_21095_, _21094_, _18700_);
  not (_21096_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand (_21097_, _18653_, _21096_);
  or (_21098_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_21099_, _21098_, _21097_);
  and (_21100_, _21099_, _18873_);
  or (_21101_, _21100_, _21095_);
  or (_21102_, _21101_, _21091_);
  and (_21103_, _21102_, _18699_);
  nand (_21104_, _18653_, _20465_);
  or (_21105_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_21106_, _21105_, _21104_);
  and (_21107_, _21106_, _18873_);
  nand (_21108_, _18653_, _20670_);
  or (_21109_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_21110_, _21109_, _21108_);
  and (_21111_, _21110_, _18710_);
  nand (_21112_, _18653_, _20261_);
  or (_21113_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_21114_, _21113_, _21112_);
  and (_21115_, _21114_, _20905_);
  or (_21116_, _21115_, _21111_);
  or (_21117_, _21116_, _21107_);
  and (_21118_, _21117_, _18639_);
  not (_21119_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nand (_21120_, _18653_, _21119_);
  or (_21121_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_21122_, _21121_, _21120_);
  and (_21123_, _21122_, _18707_);
  or (_21124_, _21123_, _21118_);
  nor (_21125_, _21124_, _21103_);
  nor (_21126_, _21125_, _18694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _21126_, _21081_);
  and (_21127_, _18694_, word_in[5]);
  nand (_21128_, _18653_, _20477_);
  or (_21129_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_21130_, _21129_, _21128_);
  and (_21131_, _21130_, _18873_);
  nand (_21132_, _18653_, _20682_);
  or (_21133_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_21134_, _21133_, _21132_);
  and (_21135_, _21134_, _18710_);
  nand (_21136_, _18653_, _20273_);
  or (_21137_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_21138_, _21137_, _21136_);
  and (_21139_, _21138_, _20905_);
  or (_21140_, _21139_, _21135_);
  or (_21141_, _21140_, _21131_);
  and (_21142_, _21141_, _18639_);
  nand (_21143_, _18653_, _19859_);
  or (_21144_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_21145_, _21144_, _21143_);
  and (_21146_, _21145_, _18710_);
  not (_21147_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nand (_21148_, _18653_, _21147_);
  or (_21149_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_21150_, _21149_, _21148_);
  and (_21151_, _21150_, _20905_);
  or (_21152_, _21151_, _21146_);
  nand (_21153_, _18653_, _20066_);
  or (_21154_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_21155_, _21154_, _21153_);
  and (_21156_, _21155_, _18700_);
  not (_21157_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nand (_21158_, _18653_, _21157_);
  or (_21159_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_21160_, _21159_, _21158_);
  and (_21161_, _21160_, _18873_);
  or (_21162_, _21161_, _21156_);
  or (_21163_, _21162_, _21152_);
  and (_21164_, _21163_, _18699_);
  not (_21165_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nand (_21166_, _18653_, _21165_);
  or (_21167_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_21168_, _21167_, _21166_);
  and (_21169_, _21168_, _18707_);
  or (_21170_, _21169_, _21164_);
  nor (_21171_, _21170_, _21142_);
  nor (_21172_, _21171_, _18694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _21172_, _21127_);
  and (_21173_, _18694_, word_in[6]);
  nand (_21174_, _18653_, _20490_);
  or (_21175_, _18653_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_21176_, _21175_, _21174_);
  and (_21177_, _21176_, _18873_);
  nand (_21178_, _18653_, _20694_);
  or (_21179_, _18653_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_21180_, _21179_, _21178_);
  and (_21181_, _21180_, _18710_);
  nand (_21182_, _18653_, _20286_);
  or (_21183_, _18653_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_21184_, _21183_, _21182_);
  and (_21185_, _21184_, _20905_);
  or (_21186_, _21185_, _21181_);
  or (_21187_, _21186_, _21177_);
  and (_21188_, _21187_, _18639_);
  nand (_21189_, _18653_, _19871_);
  or (_21190_, _18653_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_21191_, _21190_, _21189_);
  and (_21192_, _21191_, _18710_);
  not (_21193_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nand (_21194_, _18653_, _21193_);
  or (_21195_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_21196_, _21195_, _21194_);
  and (_21197_, _21196_, _18873_);
  or (_21198_, _21197_, _21192_);
  nand (_21199_, _18653_, _20076_);
  or (_21200_, _18653_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_21201_, _21200_, _21199_);
  and (_21202_, _21201_, _18700_);
  not (_21203_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nand (_21204_, _18653_, _21203_);
  or (_21205_, _18653_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_21206_, _21205_, _21204_);
  and (_21207_, _21206_, _20905_);
  or (_21208_, _21207_, _21202_);
  or (_21209_, _21208_, _21198_);
  and (_21210_, _21209_, _18699_);
  not (_21211_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nand (_21212_, _18653_, _21211_);
  or (_21213_, _18653_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_21214_, _21213_, _21212_);
  and (_21215_, _21214_, _18707_);
  or (_21216_, _21215_, _21210_);
  nor (_21217_, _21216_, _21188_);
  nor (_21218_, _21217_, _18694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _21218_, _21173_);
  and (_21219_, _18808_, word_in[8]);
  nand (_21220_, _18653_, _19268_);
  or (_21221_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_21222_, _21221_, _21220_);
  and (_21223_, _21222_, _18809_);
  and (_21224_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_21225_, _18653_, _20927_);
  or (_21226_, _21225_, _21224_);
  and (_21227_, _21226_, _18815_);
  nor (_21228_, _21227_, _21223_);
  nor (_21229_, _21228_, _18758_);
  nand (_21230_, _18653_, _19688_);
  or (_21231_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_21232_, _21231_, _21230_);
  and (_21233_, _21232_, _18809_);
  nand (_21234_, _18653_, _19899_);
  or (_21235_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_21236_, _21235_, _21234_);
  and (_21237_, _21236_, _18815_);
  or (_21238_, _21237_, _21233_);
  and (_21239_, _21238_, _18758_);
  or (_21240_, _21239_, _21229_);
  and (_21241_, _21240_, _18756_);
  nand (_21242_, _18653_, _20109_);
  or (_21243_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_21244_, _21243_, _21242_);
  and (_21245_, _21244_, _18809_);
  nand (_21246_, _18653_, _20312_);
  or (_21247_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_21248_, _21247_, _21246_);
  and (_21249_, _21248_, _18815_);
  nor (_21250_, _21249_, _21245_);
  nor (_21251_, _21250_, _18758_);
  nand (_21252_, _18653_, _20518_);
  or (_21253_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_21254_, _21253_, _21252_);
  and (_21255_, _21254_, _18809_);
  nand (_21256_, _18653_, _20719_);
  or (_21257_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_21258_, _21257_, _21256_);
  and (_21259_, _21258_, _18815_);
  or (_21260_, _21259_, _21255_);
  and (_21261_, _21260_, _18758_);
  nor (_21262_, _21261_, _21251_);
  nor (_21263_, _21262_, _18756_);
  nor (_21264_, _21263_, _21241_);
  nor (_21265_, _21264_, _18808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _21265_, _21219_);
  and (_21266_, _18808_, word_in[9]);
  nand (_21267_, _18653_, _19284_);
  or (_21268_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_21269_, _21268_, _21267_);
  and (_21270_, _21269_, _18809_);
  and (_21271_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_21272_, _18653_, _20963_);
  or (_21273_, _21272_, _21271_);
  and (_21274_, _21273_, _18815_);
  nor (_21275_, _21274_, _21270_);
  nor (_21276_, _21275_, _18758_);
  nand (_21277_, _18653_, _19701_);
  or (_21278_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_21279_, _21278_, _21277_);
  and (_21280_, _21279_, _18809_);
  nand (_21281_, _18653_, _19913_);
  or (_21282_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_21283_, _21282_, _21281_);
  and (_21284_, _21283_, _18815_);
  or (_21285_, _21284_, _21280_);
  and (_21286_, _21285_, _18758_);
  or (_21287_, _21286_, _21276_);
  and (_21288_, _21287_, _18756_);
  nand (_21289_, _18653_, _20120_);
  or (_21290_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_21291_, _21290_, _21289_);
  and (_21292_, _21291_, _18809_);
  nand (_21293_, _18653_, _20325_);
  or (_21294_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_21295_, _21294_, _21293_);
  and (_21296_, _21295_, _18815_);
  nor (_21297_, _21296_, _21292_);
  nor (_21298_, _21297_, _18758_);
  nand (_21299_, _18653_, _20532_);
  or (_21300_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_21301_, _21300_, _21299_);
  and (_21302_, _21301_, _18809_);
  nand (_21303_, _18653_, _20734_);
  or (_21304_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_21305_, _21304_, _21303_);
  and (_21306_, _21305_, _18815_);
  or (_21307_, _21306_, _21302_);
  and (_21308_, _21307_, _18758_);
  nor (_21309_, _21308_, _21298_);
  nor (_21310_, _21309_, _18756_);
  nor (_21311_, _21310_, _21288_);
  nor (_21312_, _21311_, _18808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _21312_, _21266_);
  and (_21313_, _18808_, word_in[10]);
  nand (_21314_, _18653_, _19297_);
  or (_21315_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_21316_, _21315_, _21314_);
  and (_21317_, _21316_, _18809_);
  and (_21318_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_21319_, _18653_, _21019_);
  or (_21320_, _21319_, _21318_);
  and (_21321_, _21320_, _18815_);
  nor (_21322_, _21321_, _21317_);
  nor (_21323_, _21322_, _18758_);
  nand (_21324_, _18653_, _19715_);
  or (_21325_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_21326_, _21325_, _21324_);
  and (_21327_, _21326_, _18809_);
  nand (_21328_, _18653_, _19926_);
  or (_21329_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_21330_, _21329_, _21328_);
  and (_21331_, _21330_, _18815_);
  or (_21332_, _21331_, _21327_);
  and (_21333_, _21332_, _18758_);
  or (_21334_, _21333_, _21323_);
  and (_21335_, _21334_, _18756_);
  nand (_21336_, _18653_, _20135_);
  or (_21337_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_21338_, _21337_, _21336_);
  and (_21339_, _21338_, _18809_);
  nand (_21340_, _18653_, _20339_);
  or (_21341_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_21342_, _21341_, _21340_);
  and (_21343_, _21342_, _18815_);
  nor (_21344_, _21343_, _21339_);
  nor (_21345_, _21344_, _18758_);
  nand (_21346_, _18653_, _20544_);
  or (_21347_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_21348_, _21347_, _21346_);
  and (_21349_, _21348_, _18809_);
  nand (_21350_, _18653_, _20748_);
  or (_21351_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_21352_, _21351_, _21350_);
  and (_21353_, _21352_, _18815_);
  or (_21354_, _21353_, _21349_);
  and (_21355_, _21354_, _18758_);
  nor (_21356_, _21355_, _21345_);
  nor (_21357_, _21356_, _18756_);
  nor (_21358_, _21357_, _21335_);
  nor (_21359_, _21358_, _18808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _21359_, _21313_);
  and (_21360_, _18808_, word_in[11]);
  nand (_21361_, _18653_, _19311_);
  or (_21362_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_21363_, _21362_, _21361_);
  and (_21364_, _21363_, _18809_);
  and (_21365_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_21366_, _18653_, _21040_);
  or (_21367_, _21366_, _21365_);
  and (_21368_, _21367_, _18815_);
  nor (_21369_, _21368_, _21364_);
  nor (_21370_, _21369_, _18758_);
  nand (_21371_, _18653_, _19727_);
  or (_21372_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_21373_, _21372_, _21371_);
  and (_21374_, _21373_, _18809_);
  nand (_21375_, _18653_, _19939_);
  or (_21376_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_21377_, _21376_, _21375_);
  and (_21378_, _21377_, _18815_);
  or (_21379_, _21378_, _21374_);
  and (_21380_, _21379_, _18758_);
  or (_21381_, _21380_, _21370_);
  and (_21382_, _21381_, _18756_);
  nand (_21383_, _18653_, _20147_);
  or (_21384_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_21385_, _21384_, _21383_);
  and (_21386_, _21385_, _18809_);
  nand (_21387_, _18653_, _20353_);
  or (_21388_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_21389_, _21388_, _21387_);
  and (_21390_, _21389_, _18815_);
  nor (_21391_, _21390_, _21386_);
  nor (_21392_, _21391_, _18758_);
  nand (_21393_, _18653_, _20557_);
  or (_21394_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_21395_, _21394_, _21393_);
  and (_21396_, _21395_, _18809_);
  nand (_21397_, _18653_, _20760_);
  or (_21398_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_21399_, _21398_, _21397_);
  and (_21400_, _21399_, _18815_);
  or (_21401_, _21400_, _21396_);
  and (_21402_, _21401_, _18758_);
  nor (_21403_, _21402_, _21392_);
  nor (_21404_, _21403_, _18756_);
  nor (_21405_, _21404_, _21382_);
  nor (_21406_, _21405_, _18808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _21406_, _21360_);
  and (_21407_, _18808_, word_in[12]);
  nand (_21408_, _18653_, _19325_);
  or (_21409_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_21410_, _21409_, _21408_);
  and (_21411_, _21410_, _18809_);
  and (_21412_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_21413_, _18653_, _21096_);
  or (_21414_, _21413_, _21412_);
  and (_21415_, _21414_, _18815_);
  nor (_21416_, _21415_, _21411_);
  nor (_21417_, _21416_, _18758_);
  nand (_21418_, _18653_, _19739_);
  or (_21419_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_21420_, _21419_, _21418_);
  and (_21421_, _21420_, _18809_);
  nand (_21422_, _18653_, _19950_);
  or (_21423_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_21424_, _21423_, _21422_);
  and (_21425_, _21424_, _18815_);
  or (_21426_, _21425_, _21421_);
  and (_21427_, _21426_, _18758_);
  or (_21428_, _21427_, _21417_);
  and (_21429_, _21428_, _18756_);
  nand (_21430_, _18653_, _20158_);
  or (_21431_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_21432_, _21431_, _21430_);
  and (_21433_, _21432_, _18809_);
  nand (_21434_, _18653_, _20363_);
  or (_21435_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_21436_, _21435_, _21434_);
  and (_21437_, _21436_, _18815_);
  nor (_21438_, _21437_, _21433_);
  nor (_21439_, _21438_, _18758_);
  nand (_21440_, _18653_, _20568_);
  or (_21441_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_21442_, _21441_, _21440_);
  and (_21443_, _21442_, _18809_);
  nand (_21444_, _18653_, _20772_);
  or (_21445_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_21446_, _21445_, _21444_);
  and (_21447_, _21446_, _18815_);
  or (_21448_, _21447_, _21443_);
  and (_21449_, _21448_, _18758_);
  nor (_21450_, _21449_, _21439_);
  nor (_21451_, _21450_, _18756_);
  nor (_21452_, _21451_, _21429_);
  nor (_21453_, _21452_, _18808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _21453_, _21407_);
  and (_21454_, _18808_, word_in[13]);
  nand (_21455_, _18653_, _19337_);
  or (_21456_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_21457_, _21456_, _21455_);
  and (_21458_, _21457_, _18809_);
  and (_21459_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_21460_, _18653_, _21157_);
  or (_21461_, _21460_, _21459_);
  and (_21462_, _21461_, _18815_);
  nor (_21463_, _21462_, _21458_);
  nor (_21464_, _21463_, _18758_);
  nand (_21465_, _18653_, _19751_);
  or (_21466_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_21467_, _21466_, _21465_);
  and (_21468_, _21467_, _18809_);
  nand (_21469_, _18653_, _19962_);
  or (_21470_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_21471_, _21470_, _21469_);
  and (_21472_, _21471_, _18815_);
  or (_21473_, _21472_, _21468_);
  and (_21474_, _21473_, _18758_);
  or (_21475_, _21474_, _21464_);
  and (_21476_, _21475_, _18756_);
  nand (_21477_, _18653_, _20170_);
  or (_21478_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_21479_, _21478_, _21477_);
  and (_21480_, _21479_, _18809_);
  nand (_21481_, _18653_, _20375_);
  or (_21482_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_21483_, _21482_, _21481_);
  and (_21484_, _21483_, _18815_);
  nor (_21485_, _21484_, _21480_);
  nor (_21486_, _21485_, _18758_);
  nand (_21487_, _18653_, _20580_);
  or (_21488_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_21489_, _21488_, _21487_);
  and (_21490_, _21489_, _18809_);
  nand (_21491_, _18653_, _20785_);
  or (_21492_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_21493_, _21492_, _21491_);
  and (_21494_, _21493_, _18815_);
  or (_21495_, _21494_, _21490_);
  and (_21496_, _21495_, _18758_);
  nor (_21497_, _21496_, _21486_);
  nor (_21498_, _21497_, _18756_);
  nor (_21499_, _21498_, _21476_);
  nor (_21500_, _21499_, _18808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _21500_, _21454_);
  and (_21501_, _18808_, word_in[14]);
  nand (_21502_, _18653_, _19353_);
  or (_21503_, _18653_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_21504_, _21503_, _21502_);
  and (_21505_, _21504_, _18809_);
  and (_21506_, _18653_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_21507_, _18653_, _21193_);
  or (_21508_, _21507_, _21506_);
  and (_21509_, _21508_, _18815_);
  nor (_21510_, _21509_, _21505_);
  nor (_21511_, _21510_, _18758_);
  nand (_21512_, _18653_, _19763_);
  or (_21513_, _18653_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_21514_, _21513_, _21512_);
  and (_21515_, _21514_, _18809_);
  nand (_21516_, _18653_, _19975_);
  or (_21517_, _18653_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_21518_, _21517_, _21516_);
  and (_21519_, _21518_, _18815_);
  or (_21520_, _21519_, _21515_);
  and (_21521_, _21520_, _18758_);
  or (_21522_, _21521_, _21511_);
  and (_21523_, _21522_, _18756_);
  nand (_21524_, _18653_, _20182_);
  or (_21525_, _18653_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_21526_, _21525_, _21524_);
  and (_21527_, _21526_, _18809_);
  nand (_21528_, _18653_, _20388_);
  or (_21529_, _18653_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_21530_, _21529_, _21528_);
  and (_21531_, _21530_, _18815_);
  nor (_21532_, _21531_, _21527_);
  nor (_21533_, _21532_, _18758_);
  nand (_21534_, _18653_, _20593_);
  or (_21535_, _18653_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_21536_, _21535_, _21534_);
  and (_21537_, _21536_, _18809_);
  nand (_21538_, _18653_, _20796_);
  or (_21539_, _18653_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_21540_, _21539_, _21538_);
  and (_21541_, _21540_, _18815_);
  or (_21542_, _21541_, _21537_);
  and (_21543_, _21542_, _18758_);
  nor (_21544_, _21543_, _21533_);
  nor (_21545_, _21544_, _18756_);
  nor (_21546_, _21545_, _21523_);
  nor (_21547_, _21546_, _18808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _21547_, _21501_);
  and (_21548_, _18960_, word_in[16]);
  and (_21549_, _20903_, _18873_);
  and (_21550_, _20899_, _20905_);
  or (_21551_, _21550_, _21549_);
  and (_21552_, _20938_, _18710_);
  and (_21553_, _20908_, _18700_);
  or (_21554_, _21553_, _21552_);
  or (_21555_, _21554_, _21551_);
  or (_21556_, _21555_, _18868_);
  and (_21557_, _20925_, _18710_);
  and (_21558_, _20930_, _20905_);
  or (_21559_, _21558_, _21557_);
  and (_21560_, _20915_, _18873_);
  and (_21561_, _20920_, _18700_);
  or (_21562_, _21561_, _21560_);
  nor (_21563_, _21562_, _21559_);
  nand (_21564_, _21563_, _18868_);
  and (_21565_, _21564_, _21556_);
  and (_21566_, _21565_, _18939_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _21566_, _21548_);
  and (_21567_, _18960_, word_in[17]);
  and (_21568_, _20946_, _18700_);
  and (_21569_, _20950_, _20905_);
  or (_21570_, _21569_, _21568_);
  and (_21571_, _20984_, _18710_);
  and (_21572_, _20955_, _18873_);
  or (_21573_, _21572_, _21571_);
  or (_21574_, _21573_, _21570_);
  or (_21575_, _21574_, _18868_);
  and (_21576_, _20961_, _18873_);
  and (_21577_, _20966_, _20905_);
  or (_21578_, _21577_, _21576_);
  and (_21579_, _20971_, _18710_);
  and (_21580_, _20976_, _18700_);
  or (_21581_, _21580_, _21579_);
  nor (_21582_, _21581_, _21578_);
  nand (_21583_, _21582_, _18868_);
  and (_21584_, _21583_, _21575_);
  and (_21585_, _21584_, _18939_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _21585_, _21567_);
  and (_21586_, _18960_, word_in[18]);
  and (_21587_, _21030_, _18710_);
  and (_21588_, _20996_, _18873_);
  or (_21589_, _21588_, _21587_);
  and (_21590_, _21000_, _18700_);
  and (_21591_, _20992_, _20905_);
  or (_21592_, _21591_, _21590_);
  or (_21593_, _21592_, _21589_);
  or (_21594_, _21593_, _18868_);
  and (_21595_, _21007_, _18873_);
  and (_21596_, _21022_, _20905_);
  or (_21597_, _21596_, _21595_);
  and (_21598_, _21017_, _18710_);
  and (_21599_, _21012_, _18700_);
  or (_21600_, _21599_, _21598_);
  nor (_21601_, _21600_, _21597_);
  nand (_21602_, _21601_, _18868_);
  and (_21603_, _21602_, _21594_);
  and (_21604_, _21603_, _18939_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _21604_, _21586_);
  and (_21605_, _18960_, word_in[19]);
  and (_21606_, _21076_, _18710_);
  and (_21607_, _21069_, _18873_);
  or (_21608_, _21607_, _21606_);
  and (_21609_, _21060_, _18700_);
  and (_21610_, _21064_, _20905_);
  or (_21611_, _21610_, _21609_);
  or (_21612_, _21611_, _21608_);
  or (_21613_, _21612_, _18868_);
  and (_21614_, _21038_, _18873_);
  and (_21615_, _21043_, _20905_);
  or (_21616_, _21615_, _21614_);
  and (_21617_, _21048_, _18710_);
  and (_21618_, _21053_, _18700_);
  or (_21619_, _21618_, _21617_);
  nor (_21620_, _21619_, _21616_);
  nand (_21621_, _21620_, _18868_);
  and (_21622_, _21621_, _21613_);
  and (_21623_, _21622_, _18939_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _21623_, _21605_);
  and (_21624_, _18960_, word_in[20]);
  and (_21625_, _21094_, _18710_);
  and (_21626_, _21084_, _18873_);
  or (_21627_, _21626_, _21625_);
  and (_21628_, _21089_, _18700_);
  and (_21629_, _21099_, _20905_);
  or (_21630_, _21629_, _21628_);
  nor (_21631_, _21630_, _21627_);
  nand (_21632_, _21631_, _18868_);
  and (_21633_, _21110_, _18873_);
  and (_21634_, _21106_, _20905_);
  or (_21635_, _21634_, _21633_);
  and (_21636_, _21122_, _18710_);
  and (_21637_, _21114_, _18700_);
  or (_21638_, _21637_, _21636_);
  or (_21639_, _21638_, _21635_);
  or (_21640_, _21639_, _18868_);
  and (_21641_, _21640_, _21632_);
  and (_21642_, _21641_, _18939_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _21642_, _21624_);
  and (_21643_, _18960_, word_in[21]);
  and (_21644_, _21168_, _18710_);
  and (_21645_, _21134_, _18873_);
  or (_21646_, _21645_, _21644_);
  and (_21647_, _21138_, _18700_);
  and (_21648_, _21130_, _20905_);
  or (_21649_, _21648_, _21647_);
  or (_21650_, _21649_, _21646_);
  or (_21651_, _21650_, _18868_);
  and (_21652_, _21155_, _18710_);
  and (_21653_, _21145_, _18873_);
  or (_21654_, _21653_, _21652_);
  and (_21655_, _21150_, _18700_);
  and (_21656_, _21160_, _20905_);
  or (_21657_, _21656_, _21655_);
  nor (_21658_, _21657_, _21654_);
  nand (_21659_, _21658_, _18868_);
  and (_21660_, _21659_, _21651_);
  and (_21661_, _21660_, _18939_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _21661_, _21643_);
  and (_21662_, _18960_, word_in[22]);
  and (_21663_, _21180_, _18873_);
  and (_21664_, _21176_, _20905_);
  or (_21665_, _21664_, _21663_);
  and (_21666_, _21214_, _18710_);
  and (_21667_, _21184_, _18700_);
  or (_21668_, _21667_, _21666_);
  or (_21669_, _21668_, _21665_);
  or (_21670_, _21669_, _18868_);
  and (_21671_, _21191_, _18873_);
  and (_21672_, _21196_, _20905_);
  or (_21673_, _21672_, _21671_);
  and (_21674_, _21201_, _18710_);
  and (_21675_, _21206_, _18700_);
  or (_21676_, _21675_, _21674_);
  nor (_21677_, _21676_, _21673_);
  nand (_21678_, _21677_, _18868_);
  and (_21679_, _21678_, _21670_);
  and (_21680_, _21679_, _18939_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _21680_, _21662_);
  and (_21681_, _19024_, word_in[24]);
  and (_21682_, _21226_, _18809_);
  and (_21683_, _21222_, _18815_);
  or (_21684_, _21683_, _21682_);
  or (_21685_, _21684_, _18964_);
  and (_21686_, _21236_, _18809_);
  and (_21687_, _21232_, _18815_);
  nor (_21688_, _21687_, _21686_);
  and (_21689_, _21688_, _18964_);
  nor (_21690_, _21689_, _18967_);
  and (_21691_, _21690_, _21685_);
  and (_21692_, _21248_, _18809_);
  and (_21693_, _21244_, _18815_);
  or (_21694_, _21693_, _21692_);
  or (_21695_, _21694_, _18964_);
  and (_21696_, _21258_, _18809_);
  and (_21697_, _21254_, _18815_);
  nor (_21698_, _21697_, _21696_);
  nand (_21699_, _21698_, _18964_);
  and (_21700_, _21699_, _18967_);
  and (_21701_, _21700_, _21695_);
  nor (_21702_, _21701_, _21691_);
  nor (_21703_, _21702_, _19024_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _21703_, _21681_);
  and (_21704_, _19024_, word_in[25]);
  or (_21705_, _21269_, _18809_);
  or (_21706_, _21273_, _18815_);
  and (_21707_, _21706_, _21705_);
  or (_21708_, _21707_, _18964_);
  or (_21709_, _21279_, _18809_);
  or (_21710_, _21283_, _18815_);
  nand (_21711_, _21710_, _21709_);
  nand (_21712_, _21711_, _18964_);
  and (_21713_, _21712_, _21708_);
  and (_21714_, _21713_, _19035_);
  and (_21715_, _21291_, _18815_);
  and (_21716_, _21295_, _18809_);
  or (_21717_, _21716_, _21715_);
  or (_21718_, _21717_, _18964_);
  and (_21719_, _21305_, _18809_);
  and (_21720_, _21301_, _18815_);
  nor (_21721_, _21720_, _21719_);
  nand (_21722_, _21721_, _18964_);
  and (_21723_, _21722_, _21718_);
  and (_21724_, _21723_, _18967_);
  nor (_21725_, _21724_, _21714_);
  nor (_21726_, _21725_, _19024_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _21726_, _21704_);
  and (_21727_, _19024_, word_in[26]);
  or (_21728_, _21326_, _18809_);
  or (_21729_, _21330_, _18815_);
  nand (_21730_, _21729_, _21728_);
  nand (_21731_, _21730_, _18964_);
  or (_21732_, _21316_, _18809_);
  or (_21733_, _21320_, _18815_);
  and (_21734_, _21733_, _21732_);
  or (_21735_, _21734_, _18964_);
  and (_21736_, _21735_, _21731_);
  and (_21737_, _21736_, _19035_);
  and (_21738_, _21338_, _18815_);
  and (_21739_, _21342_, _18809_);
  or (_21740_, _21739_, _21738_);
  or (_21741_, _21740_, _18964_);
  and (_21742_, _21352_, _18809_);
  and (_21743_, _21348_, _18815_);
  nor (_21744_, _21743_, _21742_);
  nand (_21745_, _21744_, _18964_);
  and (_21746_, _21745_, _21741_);
  and (_21747_, _21746_, _18967_);
  nor (_21748_, _21747_, _21737_);
  nor (_21749_, _21748_, _19024_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _21749_, _21727_);
  and (_21750_, _19024_, word_in[27]);
  and (_21751_, _21367_, _18809_);
  and (_21752_, _21363_, _18815_);
  or (_21753_, _21752_, _21751_);
  or (_21754_, _21753_, _18964_);
  and (_21755_, _21377_, _18809_);
  and (_21756_, _21373_, _18815_);
  nor (_21757_, _21756_, _21755_);
  and (_21758_, _21757_, _18964_);
  nor (_21759_, _21758_, _18967_);
  and (_21760_, _21759_, _21754_);
  and (_21761_, _21389_, _18809_);
  and (_21762_, _21385_, _18815_);
  or (_21763_, _21762_, _21761_);
  or (_21764_, _21763_, _18964_);
  and (_21765_, _21399_, _18809_);
  and (_21766_, _21395_, _18815_);
  nor (_21767_, _21766_, _21765_);
  nand (_21768_, _21767_, _18964_);
  and (_21769_, _21768_, _18967_);
  and (_21770_, _21769_, _21764_);
  nor (_21771_, _21770_, _21760_);
  nor (_21772_, _21771_, _19024_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _21772_, _21750_);
  and (_21773_, _19024_, word_in[28]);
  or (_21774_, _21410_, _18809_);
  or (_21775_, _21414_, _18815_);
  and (_21776_, _21775_, _21774_);
  or (_21777_, _21776_, _18964_);
  or (_21778_, _21420_, _18809_);
  or (_21779_, _21424_, _18815_);
  nand (_21780_, _21779_, _21778_);
  nand (_21781_, _21780_, _18964_);
  and (_21782_, _21781_, _21777_);
  and (_21783_, _21782_, _19035_);
  and (_21784_, _21432_, _18815_);
  and (_21785_, _21436_, _18809_);
  or (_21786_, _21785_, _21784_);
  or (_21787_, _21786_, _18964_);
  and (_21788_, _21446_, _18809_);
  and (_21789_, _21442_, _18815_);
  nor (_21790_, _21789_, _21788_);
  nand (_21791_, _21790_, _18964_);
  and (_21792_, _21791_, _21787_);
  and (_21793_, _21792_, _18967_);
  nor (_21794_, _21793_, _21783_);
  nor (_21795_, _21794_, _19024_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _21795_, _21773_);
  and (_21796_, _19024_, word_in[29]);
  and (_21797_, _21461_, _18809_);
  and (_21798_, _21457_, _18815_);
  or (_21799_, _21798_, _21797_);
  or (_21800_, _21799_, _18964_);
  and (_21801_, _21471_, _18809_);
  and (_21802_, _21467_, _18815_);
  nor (_21803_, _21802_, _21801_);
  and (_21804_, _21803_, _18964_);
  nor (_21805_, _21804_, _18967_);
  and (_21806_, _21805_, _21800_);
  and (_21807_, _21483_, _18809_);
  and (_21808_, _21479_, _18815_);
  or (_21809_, _21808_, _21807_);
  or (_21810_, _21809_, _18964_);
  and (_21811_, _21493_, _18809_);
  and (_21812_, _21489_, _18815_);
  nor (_21813_, _21812_, _21811_);
  nand (_21814_, _21813_, _18964_);
  and (_21815_, _21814_, _18967_);
  and (_21816_, _21815_, _21810_);
  nor (_21817_, _21816_, _21806_);
  nor (_21818_, _21817_, _19024_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _21818_, _21796_);
  and (_21819_, _19024_, word_in[30]);
  or (_21820_, _21504_, _18809_);
  or (_21821_, _21508_, _18815_);
  and (_21822_, _21821_, _21820_);
  or (_21823_, _21822_, _18964_);
  or (_21824_, _21514_, _18809_);
  or (_21825_, _21518_, _18815_);
  nand (_21826_, _21825_, _21824_);
  nand (_21827_, _21826_, _18964_);
  and (_21828_, _21827_, _21823_);
  and (_21829_, _21828_, _19035_);
  and (_21830_, _21526_, _18815_);
  and (_21831_, _21530_, _18809_);
  or (_21832_, _21831_, _21830_);
  or (_21833_, _21832_, _18964_);
  and (_21834_, _21540_, _18809_);
  and (_21835_, _21536_, _18815_);
  nor (_21836_, _21835_, _21834_);
  nand (_21837_, _21836_, _18964_);
  and (_21838_, _21837_, _21833_);
  and (_21839_, _21838_, _18967_);
  nor (_21840_, _21839_, _21829_);
  nor (_21841_, _21840_, _19024_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _21841_, _21819_);
  not (_21842_, first_instr);
  nor (_21843_, pc_log_change, _21842_);
  or (_00001_, _21843_, rst);
  or (_21844_, pc_log_change_r, cy_reg);
  nand (_21845_, pc_log_change_r, _26928_);
  and (_00000_, _21845_, _21844_);
  and (_21846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21847_, _21846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_21848_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_21849_, _21848_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_21850_, _21849_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_21851_, _21850_, _21847_);
  and (_21852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_21853_, _21852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_21854_, _21853_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_21855_, _21854_, _21851_);
  and (_21856_, _21855_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_21857_, _21856_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_21858_, _21857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21859_, _21858_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_21860_, _21858_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_21861_, _21860_, _21859_);
  and (_21862_, _21861_, cy_reg);
  nor (_21863_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_21864_, _21863_);
  and (_21865_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _16515_);
  and (_21866_, _21846_, _16527_);
  nor (_21867_, _21846_, _16527_);
  nor (_21868_, _21867_, _21866_);
  nor (_21869_, _21868_, _16515_);
  nor (_21870_, _21869_, _21865_);
  not (_21871_, _21870_);
  and (_21872_, _16523_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21873_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _16519_);
  nor (_21874_, _21873_, _21872_);
  and (_21875_, _21874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21876_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21877_, _21876_, _21875_);
  nor (_21878_, _21877_, _18894_);
  and (_21879_, _21877_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_21880_, _21879_, _21878_);
  nor (_21881_, _21880_, _21871_);
  nor (_21882_, _21877_, _19167_);
  and (_21883_, _21877_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_21884_, _21883_, _21882_);
  nor (_21885_, _21884_, _21870_);
  nor (_21886_, _21885_, _21881_);
  nor (_21887_, _21886_, _21864_);
  and (_21888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _16515_);
  not (_21889_, _21888_);
  nor (_21890_, _21877_, _18865_);
  and (_21891_, _21877_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_21892_, _21891_, _21890_);
  nor (_21893_, _21892_, _21871_);
  not (_21894_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_21895_, _21877_, _21894_);
  and (_21896_, _21877_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_21897_, _21896_, _21895_);
  nor (_21898_, _21897_, _21870_);
  nor (_21899_, _21898_, _21893_);
  nor (_21900_, _21899_, _21889_);
  nor (_21901_, _21900_, _21887_);
  and (_21902_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_21903_, _21902_);
  nor (_21904_, _21877_, _18931_);
  and (_21905_, _21877_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_21906_, _21905_, _21904_);
  nor (_21907_, _21906_, _21871_);
  not (_21908_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_21909_, _21877_, _21908_);
  and (_21910_, _21877_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_21911_, _21910_, _21909_);
  nor (_21912_, _21911_, _21870_);
  nor (_21913_, _21912_, _21907_);
  nor (_21914_, _21913_, _21903_);
  and (_21915_, _16519_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_21916_, _21915_);
  nor (_21917_, _21877_, _18906_);
  and (_21918_, _21877_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_21919_, _21918_, _21917_);
  nor (_21920_, _21919_, _21871_);
  nor (_21921_, _21877_, _19195_);
  and (_21922_, _21877_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_21923_, _21922_, _21921_);
  nor (_21924_, _21923_, _21870_);
  nor (_21925_, _21924_, _21920_);
  nor (_21926_, _21925_, _21916_);
  nor (_21927_, _21926_, _21914_);
  and (_21928_, _21927_, _21901_);
  not (_21929_, _21877_);
  and (_21930_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_21931_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_21932_, _21931_, _21930_);
  and (_21933_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_21934_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_21935_, _21934_, _21933_);
  and (_21936_, _21935_, _21932_);
  and (_21937_, _21936_, _21929_);
  and (_21938_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_21939_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_21940_, _21939_, _21938_);
  and (_21941_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_21942_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_21943_, _21942_, _21941_);
  and (_21944_, _21943_, _21940_);
  and (_21945_, _21944_, _21877_);
  or (_21946_, _21945_, _21871_);
  nor (_21947_, _21946_, _21937_);
  and (_21948_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_21949_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_21950_, _21949_, _21948_);
  and (_21951_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_21952_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_21953_, _21952_, _21951_);
  and (_21954_, _21953_, _21950_);
  nor (_21955_, _21954_, _21877_);
  and (_21956_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_21957_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_21958_, _21957_, _21956_);
  and (_21959_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_21960_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_21961_, _21960_, _21959_);
  and (_21962_, _21961_, _21958_);
  nor (_21963_, _21962_, _21929_);
  or (_21964_, _21963_, _21955_);
  and (_21965_, _21964_, _21871_);
  nor (_21966_, _21965_, _21947_);
  nor (_21967_, _21966_, _21928_);
  nor (_21968_, _21857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21969_, _21968_, _21858_);
  and (_21970_, _21969_, _21967_);
  nor (_21971_, _21969_, _21967_);
  nor (_21972_, _21971_, _21970_);
  not (_21973_, _21972_);
  nor (_21974_, _21856_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_21975_, _21974_, _21857_);
  nor (_21976_, _21975_, _21967_);
  and (_21977_, _21975_, _21967_);
  not (_21978_, _21977_);
  nor (_21979_, _21855_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_21980_, _21979_, _21856_);
  and (_21981_, _21980_, _21967_);
  and (_21982_, _21853_, _21851_);
  nor (_21983_, _21982_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_21984_, _21982_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_21985_, _21984_, _21983_);
  and (_21986_, _21985_, _21967_);
  nor (_21987_, _21985_, _21967_);
  and (_21988_, _21851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_21989_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_21990_, _21989_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_21991_, _21990_, _21982_);
  and (_21992_, _21991_, _21967_);
  nor (_21993_, _21991_, _21967_);
  nor (_21994_, _21993_, _21992_);
  not (_21995_, _21994_);
  nor (_21996_, _21988_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_21997_, _21996_, _21989_);
  and (_21998_, _21997_, _21967_);
  nor (_21999_, _21851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22000_, _21999_, _21988_);
  and (_22001_, _22000_, _21967_);
  nor (_22002_, _21997_, _21967_);
  nor (_22003_, _22002_, _21998_);
  and (_22004_, _21849_, _21847_);
  nor (_22005_, _22004_, _16540_);
  and (_22006_, _22004_, _16540_);
  nor (_22007_, _22006_, _22005_);
  not (_22008_, _22007_);
  and (_22009_, _22008_, _21967_);
  nor (_22010_, _22008_, _21967_);
  and (_22011_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_22012_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_22013_, _22012_, _22011_);
  and (_22014_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_22015_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_22016_, _22015_, _22014_);
  and (_22017_, _22016_, _22013_);
  and (_22018_, _22017_, _21929_);
  and (_22019_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_22020_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_22021_, _22020_, _22019_);
  and (_22022_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_22023_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_22024_, _22023_, _22022_);
  and (_22025_, _22024_, _22021_);
  and (_22026_, _22025_, _21877_);
  or (_22027_, _22026_, _21871_);
  nor (_22028_, _22027_, _22018_);
  and (_22029_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_22030_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_22031_, _22030_, _22029_);
  and (_22032_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_22033_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_22034_, _22033_, _22032_);
  and (_22035_, _22034_, _22031_);
  nor (_22036_, _22035_, _21877_);
  and (_22037_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_22038_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_22039_, _22038_, _22037_);
  and (_22040_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_22041_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_22042_, _22041_, _22040_);
  and (_22043_, _22042_, _22039_);
  nor (_22044_, _22043_, _21929_);
  or (_22045_, _22044_, _22036_);
  and (_22046_, _22045_, _21871_);
  nor (_22047_, _22046_, _22028_);
  nor (_22048_, _22047_, _21928_);
  and (_22049_, _21848_, _21847_);
  nor (_22050_, _22049_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_22051_, _22050_, _22004_);
  and (_22052_, _22051_, _22048_);
  nor (_22053_, _22051_, _22048_);
  nor (_22054_, _22053_, _22052_);
  not (_22055_, _22054_);
  and (_22056_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_22057_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_22058_, _22057_, _22056_);
  and (_22059_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_22060_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_22061_, _22060_, _22059_);
  and (_22062_, _22061_, _22058_);
  and (_22063_, _22062_, _21929_);
  and (_22064_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_22065_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_22066_, _22065_, _22064_);
  and (_22067_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_22068_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_22069_, _22068_, _22067_);
  and (_22070_, _22069_, _22066_);
  and (_22071_, _22070_, _21877_);
  or (_22072_, _22071_, _21871_);
  nor (_22073_, _22072_, _22063_);
  and (_22074_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_22075_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_22076_, _22075_, _22074_);
  and (_22077_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_22078_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_22079_, _22078_, _22077_);
  and (_22080_, _22079_, _22076_);
  nor (_22081_, _22080_, _21877_);
  and (_22082_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_22083_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_22084_, _22083_, _22082_);
  and (_22085_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_22086_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_22087_, _22086_, _22085_);
  and (_22088_, _22087_, _22084_);
  nor (_22089_, _22088_, _21929_);
  or (_22090_, _22089_, _22081_);
  and (_22091_, _22090_, _21871_);
  nor (_22092_, _22091_, _22073_);
  nor (_22093_, _22092_, _21928_);
  and (_22094_, _21847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_22095_, _22094_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_22096_, _22095_, _22049_);
  and (_22097_, _22096_, _22093_);
  nor (_22098_, _22096_, _22093_);
  nor (_22099_, _22098_, _22097_);
  not (_22100_, _22099_);
  and (_22101_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_22102_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_22103_, _22102_, _22101_);
  and (_22104_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_22105_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_22106_, _22105_, _22104_);
  and (_22107_, _22106_, _22103_);
  and (_22108_, _22107_, _21929_);
  and (_22109_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_22110_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_22111_, _22110_, _22109_);
  and (_22112_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_22113_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_22114_, _22113_, _22112_);
  and (_22115_, _22114_, _22111_);
  and (_22116_, _22115_, _21877_);
  or (_22117_, _22116_, _21871_);
  nor (_22118_, _22117_, _22108_);
  and (_22119_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_22120_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_22121_, _22120_, _22119_);
  and (_22122_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_22123_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_22124_, _22123_, _22122_);
  and (_22125_, _22124_, _22121_);
  nor (_22126_, _22125_, _21877_);
  and (_22127_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_22128_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_22129_, _22128_, _22127_);
  and (_22130_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_22131_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_22132_, _22131_, _22130_);
  and (_22133_, _22132_, _22129_);
  nor (_22134_, _22133_, _21929_);
  or (_22135_, _22134_, _22126_);
  and (_22136_, _22135_, _21871_);
  nor (_22137_, _22136_, _22118_);
  nor (_22138_, _22137_, _21928_);
  nor (_22139_, _21847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_22140_, _22139_, _22094_);
  and (_22141_, _22140_, _22138_);
  not (_22142_, _21868_);
  and (_22143_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_22144_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_22145_, _22144_, _22143_);
  and (_22146_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_22147_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_22148_, _22147_, _22146_);
  and (_22149_, _22148_, _22145_);
  and (_22150_, _22149_, _21929_);
  and (_22151_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_22152_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_22153_, _22152_, _22151_);
  and (_22154_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_22155_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_22156_, _22155_, _22154_);
  and (_22157_, _22156_, _22153_);
  and (_22158_, _22157_, _21877_);
  or (_22159_, _22158_, _21871_);
  nor (_22160_, _22159_, _22150_);
  and (_22161_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_22162_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_22163_, _22162_, _22161_);
  and (_22164_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_22165_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_22166_, _22165_, _22164_);
  and (_22167_, _22166_, _22163_);
  nor (_22168_, _22167_, _21877_);
  and (_22169_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_22170_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_22171_, _22170_, _22169_);
  and (_22172_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_22173_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_22174_, _22173_, _22172_);
  and (_22175_, _22174_, _22171_);
  nor (_22176_, _22175_, _21929_);
  or (_22177_, _22176_, _22168_);
  and (_22178_, _22177_, _21871_);
  nor (_22179_, _22178_, _22160_);
  nor (_22180_, _22179_, _21928_);
  and (_22181_, _22180_, _22142_);
  nor (_22182_, _22180_, _22142_);
  nor (_22183_, _22182_, _22181_);
  not (_22184_, _22183_);
  not (_22185_, _21874_);
  and (_22186_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_22187_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_22188_, _22187_, _22186_);
  and (_22189_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_22190_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_22191_, _22190_, _22189_);
  and (_22192_, _22191_, _22188_);
  and (_22193_, _22192_, _21929_);
  and (_22194_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_22195_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_22196_, _22195_, _22194_);
  and (_22197_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_22198_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_22199_, _22198_, _22197_);
  and (_22200_, _22199_, _22196_);
  and (_22201_, _22200_, _21877_);
  or (_22202_, _22201_, _21871_);
  nor (_22203_, _22202_, _22193_);
  and (_22204_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_22205_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_22206_, _22205_, _22204_);
  and (_22207_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_22208_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_22209_, _22208_, _22207_);
  and (_22210_, _22209_, _22206_);
  nor (_22211_, _22210_, _21877_);
  and (_22212_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_22213_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_22214_, _22213_, _22212_);
  and (_22215_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_22216_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_22217_, _22216_, _22215_);
  and (_22218_, _22217_, _22214_);
  nor (_22219_, _22218_, _21929_);
  or (_22220_, _22219_, _22211_);
  and (_22221_, _22220_, _21871_);
  nor (_22222_, _22221_, _22203_);
  nor (_22223_, _22222_, _21928_);
  and (_22224_, _22223_, _22185_);
  and (_22225_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_22226_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_22227_, _22226_, _22225_);
  and (_22228_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_22229_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_22230_, _22229_, _22228_);
  and (_22231_, _22230_, _22227_);
  and (_22232_, _22231_, _21929_);
  and (_22233_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_22234_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_22235_, _22234_, _22233_);
  and (_22236_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_22237_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_22238_, _22237_, _22236_);
  and (_22239_, _22238_, _22235_);
  and (_22240_, _22239_, _21877_);
  or (_22241_, _22240_, _21871_);
  nor (_22242_, _22241_, _22232_);
  and (_22243_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_22244_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_22245_, _22244_, _22243_);
  and (_22246_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_22247_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_22248_, _22247_, _22246_);
  and (_22249_, _22248_, _22245_);
  nor (_22250_, _22249_, _21877_);
  and (_22251_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_22252_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_22253_, _22252_, _22251_);
  and (_22254_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_22255_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_22256_, _22255_, _22254_);
  and (_22257_, _22256_, _22253_);
  nor (_22258_, _22257_, _21929_);
  or (_22259_, _22258_, _22250_);
  and (_22260_, _22259_, _21871_);
  nor (_22261_, _22260_, _22242_);
  nor (_22262_, _22261_, _21928_);
  and (_22263_, _22262_, _16519_);
  and (_22264_, _21888_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_22265_, _21902_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_22266_, _22265_, _22264_);
  and (_22267_, _21915_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_22268_, _21863_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_22269_, _22268_, _22267_);
  and (_22270_, _22269_, _22266_);
  and (_22271_, _22270_, _21929_);
  and (_22272_, _21888_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_22273_, _21863_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_22274_, _22273_, _22272_);
  and (_22275_, _21915_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_22276_, _21902_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_22277_, _22276_, _22275_);
  and (_22278_, _22277_, _22274_);
  and (_22279_, _22278_, _21877_);
  or (_22280_, _22279_, _21871_);
  nor (_22281_, _22280_, _22271_);
  and (_22282_, _21915_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_22283_, _21863_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_22284_, _22283_, _22282_);
  and (_22285_, _21888_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_22286_, _21902_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_22287_, _22286_, _22285_);
  and (_22288_, _22287_, _22284_);
  nor (_22289_, _22288_, _21877_);
  and (_22290_, _21915_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_22291_, _21902_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_22292_, _22291_, _22290_);
  and (_22293_, _21888_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_22294_, _21863_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_22295_, _22294_, _22293_);
  and (_22296_, _22295_, _22292_);
  nor (_22297_, _22296_, _21929_);
  or (_22298_, _22297_, _22289_);
  and (_22299_, _22298_, _21871_);
  nor (_22300_, _22299_, _22281_);
  nor (_22301_, _22300_, _21928_);
  and (_22302_, _22301_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22303_, _22262_, _16519_);
  nor (_22304_, _22303_, _22263_);
  and (_22305_, _22304_, _22302_);
  nor (_22306_, _22305_, _22263_);
  nor (_22307_, _22223_, _22185_);
  nor (_22308_, _22307_, _22224_);
  not (_22309_, _22308_);
  nor (_22310_, _22309_, _22306_);
  nor (_22311_, _22310_, _22224_);
  nor (_22312_, _22311_, _22184_);
  nor (_22313_, _22312_, _22181_);
  nor (_22314_, _22140_, _22138_);
  nor (_22315_, _22314_, _22141_);
  not (_22316_, _22315_);
  nor (_22317_, _22316_, _22313_);
  nor (_22318_, _22317_, _22141_);
  nor (_22319_, _22318_, _22100_);
  nor (_22320_, _22319_, _22097_);
  nor (_22321_, _22320_, _22055_);
  nor (_22322_, _22321_, _22052_);
  nor (_22323_, _22322_, _22010_);
  or (_22324_, _22323_, _22009_);
  nor (_22325_, _22000_, _21967_);
  nor (_22326_, _22325_, _22001_);
  and (_22327_, _22326_, _22324_);
  and (_22328_, _22327_, _22003_);
  or (_22329_, _22328_, _22001_);
  nor (_22330_, _22329_, _21998_);
  nor (_22331_, _22330_, _21995_);
  nor (_22332_, _22331_, _21992_);
  nor (_22333_, _22332_, _21987_);
  or (_22334_, _22333_, _21986_);
  nor (_22335_, _21980_, _21967_);
  nor (_22336_, _22335_, _21981_);
  and (_22337_, _22336_, _22334_);
  nor (_22338_, _22337_, _21981_);
  and (_22339_, _22338_, _21978_);
  or (_22340_, _22339_, _21976_);
  nor (_22341_, _22340_, _21973_);
  nor (_22342_, _22341_, _21970_);
  and (_22343_, _21967_, _21861_);
  nor (_22344_, _21967_, _21861_);
  or (_22345_, _22344_, _22343_);
  and (_22346_, _22345_, _22342_);
  nor (_22347_, _22345_, _22342_);
  or (_22348_, _22347_, _22346_);
  nor (_22349_, _22348_, cy_reg);
  nor (_22350_, _22349_, _21862_);
  nor (_22351_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_22352_, _22350_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_22353_, _21969_, cy_reg);
  not (_22354_, cy_reg);
  and (_22355_, _22340_, _21973_);
  nor (_22356_, _22355_, _22341_);
  and (_22357_, _22356_, _22354_);
  nor (_22358_, _22357_, _22353_);
  nor (_22359_, _22358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_22360_, _22358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_22361_, _21976_, _21977_);
  nor (_22362_, _22361_, _22338_);
  and (_22363_, _22361_, _22338_);
  nor (_22364_, _22363_, _22362_);
  nor (_22365_, _22364_, cy_reg);
  and (_22366_, _21975_, cy_reg);
  nor (_22367_, _22366_, _22365_);
  and (_22368_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_22369_, _22367_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_22370_, _22336_, _22334_);
  nor (_22371_, _22370_, _22337_);
  nor (_22372_, _22371_, cy_reg);
  nor (_22373_, _21980_, _22354_);
  nor (_22374_, _22373_, _22372_);
  nor (_22375_, _22374_, _16503_);
  and (_22376_, _22374_, _16503_);
  and (_22377_, _21985_, cy_reg);
  nor (_22378_, _21986_, _21987_);
  nor (_22379_, _22378_, _22332_);
  and (_22380_, _22378_, _22332_);
  nor (_22381_, _22380_, _22379_);
  nor (_22382_, _22381_, cy_reg);
  nor (_22383_, _22382_, _22377_);
  and (_22384_, _22383_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_22385_, _22383_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_22386_, _22327_, _22001_);
  and (_22387_, _22386_, _22003_);
  nor (_22388_, _22386_, _22003_);
  nor (_22389_, _22388_, _22387_);
  nor (_22390_, _22389_, cy_reg);
  and (_22391_, _21997_, cy_reg);
  nor (_22392_, _22391_, _22390_);
  nand (_22393_, _22392_, _16491_);
  or (_22394_, _22392_, _16491_);
  and (_22395_, _22394_, _22393_);
  nor (_22396_, _22000_, _16487_);
  and (_22397_, _22000_, _16487_);
  or (_22398_, _22397_, _22396_);
  or (_22399_, _22007_, _16483_);
  nand (_22400_, _22007_, _16483_);
  and (_22401_, _22400_, _22399_);
  or (_22402_, _22401_, _22354_);
  or (_22403_, _22402_, _22398_);
  nor (_22404_, _22326_, _22324_);
  nor (_22405_, _22404_, _22327_);
  or (_22406_, _22405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_22407_, _22405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_22408_, _22407_, _22406_);
  nor (_22409_, _22009_, _22010_);
  nor (_22410_, _22409_, _22322_);
  and (_22411_, _22409_, _22322_);
  nor (_22412_, _22411_, _22410_);
  nor (_22413_, _22412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_22414_, _22412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_22415_, _22414_, _22413_);
  or (_22416_, _22415_, cy_reg);
  or (_22417_, _22416_, _22408_);
  and (_22418_, _22417_, _22403_);
  and (_22419_, _22051_, cy_reg);
  and (_22420_, _22320_, _22055_);
  nor (_22421_, _22420_, _22321_);
  and (_22422_, _22421_, _22354_);
  nor (_22423_, _22422_, _22419_);
  nor (_22424_, _22423_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_22425_, _22423_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_22426_, _22318_, _22100_);
  nor (_22427_, _22426_, _22319_);
  and (_22428_, _22427_, _22354_);
  and (_22429_, _22096_, cy_reg);
  nor (_22430_, _22429_, _22428_);
  and (_22431_, _22430_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_22432_, _22430_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_22433_, _22140_, cy_reg);
  and (_22434_, _22316_, _22313_);
  nor (_22435_, _22434_, _22317_);
  and (_22436_, _22435_, _22354_);
  nor (_22437_, _22436_, _22433_);
  and (_22438_, _22437_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_22439_, _22437_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_22440_, _22311_, _22184_);
  nor (_22441_, _22440_, _22312_);
  and (_22442_, _22441_, _22354_);
  nor (_22443_, _21868_, _22354_);
  nor (_22444_, _22443_, _22442_);
  nor (_22445_, _22444_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22446_, _22444_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22447_, cy_reg, _16519_);
  nor (_22448_, _22304_, _22302_);
  nor (_22449_, _22448_, _22305_);
  and (_22450_, _22449_, _22354_);
  nor (_22451_, _22450_, _22447_);
  and (_22452_, _22451_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22453_, _22301_, _22354_);
  and (_22454_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_22455_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_22456_, _22455_, _22454_);
  nor (_22457_, _22456_, _22453_);
  and (_22458_, _22456_, _22301_);
  and (_22459_, _22458_, _22354_);
  or (_22460_, _22459_, _22457_);
  nor (_22461_, _22451_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_22462_, _22461_, _22460_);
  or (_22463_, _22462_, _22452_);
  and (_22464_, _22309_, _22306_);
  nor (_22465_, _22464_, _22310_);
  and (_22466_, _22465_, _22354_);
  nor (_22467_, _21874_, _22354_);
  nor (_22468_, _22467_, _22466_);
  nor (_22469_, _22468_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_22470_, _22468_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_22471_, _22470_, _22469_);
  or (_22472_, _22471_, _22463_);
  or (_22473_, _22472_, _22446_);
  or (_22474_, _22473_, _22445_);
  or (_22475_, _22474_, _22439_);
  or (_22476_, _22475_, _22438_);
  or (_22477_, _22476_, _22432_);
  or (_22478_, _22477_, _22431_);
  or (_22479_, _22478_, _22425_);
  or (_22480_, _22479_, _22424_);
  or (_22481_, _22480_, _22418_);
  or (_22482_, _22481_, _22395_);
  and (_22483_, _21991_, cy_reg);
  and (_22484_, _22330_, _21995_);
  nor (_22485_, _22484_, _22331_);
  and (_22486_, _22485_, _22354_);
  nor (_22487_, _22486_, _22483_);
  and (_22488_, _22487_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_22489_, _22487_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_22490_, _22489_, _22488_);
  or (_22491_, _22490_, _22482_);
  or (_22492_, _22491_, _22385_);
  or (_22493_, _22492_, _22384_);
  or (_22494_, _22493_, _22376_);
  or (_22495_, _22494_, _22375_);
  or (_22496_, _22495_, _22369_);
  or (_22497_, _22496_, _22368_);
  or (_22498_, _22497_, _22360_);
  or (_22499_, _22498_, _22359_);
  or (_22500_, _22499_, _22352_);
  or (_22501_, _22500_, _22351_);
  and (_22502_, _18925_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22503_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22504_, _22503_, _22502_);
  and (_22505_, _22504_, _21873_);
  nor (_22506_, _22505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22507_, _18915_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_22508_, _22507_);
  nor (_22509_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22510_, _22509_, _16523_);
  and (_22511_, _22510_, _22508_);
  and (_22512_, _19195_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22513_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22514_, _22513_, _22512_);
  and (_22515_, _22514_, _16523_);
  nor (_22516_, _22515_, _22511_);
  nor (_22517_, _22516_, _16519_);
  nor (_22518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_22519_, _21908_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22520_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22521_, _22520_, _22519_);
  and (_22522_, _22521_, _22518_);
  nor (_22523_, _22522_, _22517_);
  and (_22524_, _22523_, _22506_);
  nor (_22525_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_22526_, _22525_);
  and (_22527_, _18879_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22528_, _22527_, _16523_);
  and (_22529_, _22528_, _22526_);
  and (_22530_, _21894_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22531_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22532_, _22531_, _22530_);
  and (_22533_, _22532_, _16523_);
  nor (_22534_, _22533_, _22529_);
  nor (_22535_, _22534_, _16519_);
  nor (_22536_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_22537_, _19167_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22538_, _22537_, _22536_);
  and (_22539_, _22538_, _22518_);
  nor (_22540_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_22541_, _18887_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22542_, _22541_, _22540_);
  and (_22543_, _22542_, _21873_);
  or (_22544_, _22543_, _16515_);
  or (_22545_, _22544_, _22539_);
  nor (_22546_, _22545_, _22535_);
  nor (_22547_, _22546_, _22524_);
  nor (_22548_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22549_, _21040_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22550_, _22549_, _22548_);
  and (_22551_, _22550_, _21872_);
  nor (_22552_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22553_, _19831_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22554_, _22553_, _22552_);
  and (_22555_, _22554_, _21873_);
  nor (_22556_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22557_, _21050_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22558_, _22557_, _22556_);
  and (_22559_, _22558_, _22518_);
  nor (_22560_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22561_, _20042_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22562_, _22561_, _22560_);
  and (_22563_, _22562_, _21846_);
  or (_22564_, _22563_, _22559_);
  or (_22565_, _22564_, _22555_);
  or (_22566_, _22565_, _22551_);
  and (_22567_, _22566_, _16527_);
  nor (_22568_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22569_, _20453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22570_, _22569_, _22568_);
  and (_22571_, _22570_, _21872_);
  nor (_22572_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22573_, _20659_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22574_, _22573_, _22572_);
  and (_22575_, _22574_, _21873_);
  nor (_22576_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22577_, _20249_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22578_, _22577_, _22576_);
  and (_22579_, _22578_, _22518_);
  nor (_22580_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22581_, _21073_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22582_, _22581_, _22580_);
  and (_22583_, _22582_, _21846_);
  or (_22584_, _22583_, _22579_);
  or (_22585_, _22584_, _22575_);
  or (_22586_, _22585_, _22571_);
  and (_22587_, _22586_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_22588_, _22587_, _22567_);
  and (_22589_, _22588_, _22547_);
  nor (_22590_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22591_, _21019_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22592_, _22591_, _22590_);
  and (_22593_, _22592_, _21872_);
  nor (_22594_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22595_, _19818_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22596_, _22595_, _22594_);
  and (_22597_, _22596_, _21873_);
  nor (_22598_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22599_, _21009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22600_, _22599_, _22598_);
  and (_22601_, _22600_, _22518_);
  nor (_22602_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22603_, _20030_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22604_, _22603_, _22602_);
  and (_22605_, _22604_, _21846_);
  or (_22606_, _22605_, _22601_);
  or (_22607_, _22606_, _22597_);
  or (_22608_, _22607_, _22593_);
  and (_22609_, _22608_, _16527_);
  nor (_22610_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22611_, _20442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22612_, _22611_, _22610_);
  and (_22613_, _22612_, _21872_);
  nor (_22614_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22615_, _20645_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22616_, _22615_, _22614_);
  and (_22617_, _22616_, _21873_);
  nor (_22618_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22619_, _20237_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22620_, _22619_, _22618_);
  and (_22621_, _22620_, _22518_);
  nor (_22622_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22623_, _21027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22624_, _22623_, _22622_);
  and (_22625_, _22624_, _21846_);
  or (_22626_, _22625_, _22621_);
  or (_22627_, _22626_, _22617_);
  or (_22628_, _22627_, _22613_);
  and (_22629_, _22628_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_22630_, _22629_, _22609_);
  and (_22631_, _22630_, _22547_);
  nor (_22632_, _22631_, _22589_);
  nor (_22633_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22634_, _20963_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22635_, _22634_, _22633_);
  and (_22636_, _22635_, _21872_);
  nor (_22637_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22638_, _19806_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22639_, _22638_, _22637_);
  and (_22640_, _22639_, _21873_);
  nor (_22641_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22642_, _20973_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22643_, _22642_, _22641_);
  and (_22644_, _22643_, _22518_);
  nor (_22645_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22646_, _20016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22647_, _22646_, _22645_);
  and (_22648_, _22647_, _21846_);
  or (_22649_, _22648_, _22644_);
  or (_22650_, _22649_, _22640_);
  or (_22651_, _22650_, _22636_);
  and (_22652_, _22651_, _16527_);
  nor (_22653_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22654_, _20429_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22655_, _22654_, _22653_);
  and (_22656_, _22655_, _21872_);
  nor (_22657_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22658_, _20633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22659_, _22658_, _22657_);
  and (_22660_, _22659_, _21873_);
  nor (_22661_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22662_, _20223_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22663_, _22662_, _22661_);
  and (_22664_, _22663_, _22518_);
  nor (_22665_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22666_, _20981_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22667_, _22666_, _22665_);
  and (_22668_, _22667_, _21846_);
  or (_22669_, _22668_, _22664_);
  or (_22670_, _22669_, _22660_);
  or (_22671_, _22670_, _22656_);
  and (_22672_, _22671_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_22673_, _22672_, _22652_);
  and (_22674_, _22673_, _22547_);
  nor (_22675_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22676_, _20620_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22677_, _22676_, _22675_);
  and (_22678_, _22677_, _21873_);
  nor (_22679_, _22678_, _16527_);
  nor (_22680_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22681_, _20209_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22682_, _22681_, _22680_);
  and (_22683_, _22682_, _22518_);
  nor (_22684_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22685_, _20412_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22686_, _22685_, _22684_);
  and (_22687_, _22686_, _21872_);
  nor (_22688_, _22687_, _22683_);
  nor (_22689_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22690_, _20935_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22691_, _22690_, _22689_);
  and (_22692_, _22691_, _21846_);
  not (_22693_, _22692_);
  and (_22694_, _22693_, _22688_);
  and (_22695_, _22694_, _22679_);
  nor (_22696_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22697_, _19790_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22698_, _22697_, _22696_);
  and (_22699_, _22698_, _21873_);
  nor (_22700_, _22699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22701_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22702_, _20917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22703_, _22702_, _22701_);
  and (_22704_, _22703_, _22518_);
  nor (_22705_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22706_, _20927_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22707_, _22706_, _22705_);
  and (_22708_, _22707_, _21872_);
  nor (_22709_, _22708_, _22704_);
  nor (_22710_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22711_, _20002_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22712_, _22711_, _22710_);
  and (_22713_, _22712_, _21846_);
  not (_22714_, _22713_);
  and (_22715_, _22714_, _22709_);
  and (_22716_, _22715_, _22700_);
  nor (_22717_, _22716_, _22695_);
  and (_22718_, _22717_, _22547_);
  nor (_22719_, _22718_, _22674_);
  and (_22720_, _22719_, _22632_);
  nor (_22721_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22722_, _21096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22723_, _22722_, _22721_);
  and (_22724_, _22723_, _21872_);
  nor (_22725_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22726_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22727_, _22726_, _22725_);
  and (_22728_, _22727_, _21873_);
  nor (_22729_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22730_, _21086_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22731_, _22730_, _22729_);
  and (_22732_, _22731_, _22518_);
  nor (_22733_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22734_, _20053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22735_, _22734_, _22733_);
  and (_22736_, _22735_, _21846_);
  or (_22737_, _22736_, _22732_);
  or (_22738_, _22737_, _22728_);
  or (_22739_, _22738_, _22724_);
  and (_22740_, _22739_, _16527_);
  nor (_22741_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22742_, _20465_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22743_, _22742_, _22741_);
  and (_22744_, _22743_, _21872_);
  nor (_22745_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22746_, _20670_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22747_, _22746_, _22745_);
  and (_22748_, _22747_, _21873_);
  nor (_22749_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22750_, _20261_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22751_, _22750_, _22749_);
  and (_22752_, _22751_, _22518_);
  nor (_22753_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22754_, _21119_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22755_, _22754_, _22753_);
  and (_22756_, _22755_, _21846_);
  or (_22757_, _22756_, _22752_);
  or (_22758_, _22757_, _22748_);
  or (_22759_, _22758_, _22744_);
  and (_22760_, _22759_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_22761_, _22760_, _22740_);
  and (_22762_, _22761_, _22547_);
  nor (_22763_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22764_, _21157_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22765_, _22764_, _22763_);
  and (_22766_, _22765_, _21872_);
  nor (_22767_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22768_, _19859_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22769_, _22768_, _22767_);
  and (_22770_, _22769_, _21873_);
  nor (_22771_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22772_, _21147_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22773_, _22772_, _22771_);
  and (_22774_, _22773_, _22518_);
  nor (_22775_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22776_, _20066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22777_, _22776_, _22775_);
  and (_22778_, _22777_, _21846_);
  or (_22779_, _22778_, _22774_);
  or (_22780_, _22779_, _22770_);
  or (_22781_, _22780_, _22766_);
  and (_22782_, _22781_, _16527_);
  nor (_22783_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22784_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22785_, _22784_, _22783_);
  and (_22786_, _22785_, _21872_);
  nor (_22787_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22788_, _20682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22789_, _22788_, _22787_);
  and (_22790_, _22789_, _21873_);
  nor (_22791_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22792_, _20273_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22793_, _22792_, _22791_);
  and (_22794_, _22793_, _22518_);
  nor (_22795_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22796_, _21165_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22797_, _22796_, _22795_);
  and (_22798_, _22797_, _21846_);
  or (_22799_, _22798_, _22794_);
  or (_22800_, _22799_, _22790_);
  or (_22801_, _22800_, _22786_);
  and (_22802_, _22801_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_22803_, _22802_, _22782_);
  and (_22804_, _22803_, _22547_);
  not (_22805_, _22804_);
  and (_22806_, _22805_, _22762_);
  and (_22807_, _22806_, _22720_);
  or (_22808_, \oc8051_symbolic_cxrom1.regvalid [1], _16467_);
  and (_22809_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_22810_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22811_, _22810_, _22809_);
  and (_22812_, _22811_, _22808_);
  or (_22813_, \oc8051_symbolic_cxrom1.regvalid [13], _16467_);
  or (_22814_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22815_, _22814_, _22813_);
  and (_22816_, _16463_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22817_, _22816_, _22815_);
  or (_22818_, _22817_, _22812_);
  nor (_22819_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_22820_, _22819_, _16463_);
  nor (_22821_, _22820_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22822_, _22820_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_22823_, _22822_, _22821_);
  and (_22824_, _22823_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_22825_, _22819_, _16463_);
  nor (_22826_, _22825_, _22820_);
  nand (_22827_, \oc8051_symbolic_cxrom1.regvalid [7], _16467_);
  nand (_22828_, _22827_, _22826_);
  or (_22829_, _22828_, _22824_);
  and (_22830_, _22829_, _16459_);
  nand (_22831_, _22823_, _21894_);
  or (_22832_, _22823_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_22833_, _22832_, _22831_);
  or (_22834_, _22826_, _22833_);
  and (_22835_, _22834_, _22830_);
  or (_22836_, _22835_, _22818_);
  and (_22837_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22838_, \oc8051_symbolic_cxrom1.regvalid [0], _16467_);
  or (_22839_, _22838_, _22837_);
  and (_22840_, _22839_, _16463_);
  and (_22841_, \oc8051_symbolic_cxrom1.regvalid [4], _16467_);
  and (_22842_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22843_, _22842_, _22841_);
  and (_22844_, _22843_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_22845_, _22844_, _22840_);
  and (_22846_, _22845_, _16459_);
  and (_22847_, _22809_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_22848_, _22847_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22849_, _22847_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_22850_, _22849_, _22848_);
  or (_22851_, _22850_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_22852_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_22853_, _22852_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_22854_, _22853_, _22847_);
  and (_22855_, _22854_, _22813_);
  and (_22856_, _22855_, _22851_);
  or (_22857_, _22850_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_22858_, _22854_);
  nand (_22859_, _22850_, _19167_);
  and (_22860_, _22859_, _22858_);
  and (_22861_, _22860_, _22857_);
  or (_22862_, _22861_, _22856_);
  and (_22863_, _22862_, _22846_);
  or (_22864_, _22850_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_22865_, \oc8051_symbolic_cxrom1.regvalid [15], _16467_);
  and (_22866_, _22865_, _22854_);
  and (_22867_, _22866_, _22864_);
  or (_22868_, _22850_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_22869_, _22850_, _21894_);
  and (_22870_, _22869_, _22858_);
  and (_22871_, _22870_, _22868_);
  or (_22872_, _22871_, _22867_);
  and (_22873_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22874_, \oc8051_symbolic_cxrom1.regvalid [6], _16467_);
  or (_22875_, _22874_, _16463_);
  or (_22876_, _22875_, _22873_);
  or (_22877_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22878_, \oc8051_symbolic_cxrom1.regvalid [10], _16467_);
  and (_22879_, _22878_, _22877_);
  or (_22880_, _22879_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_22881_, _22880_, _22876_);
  and (_22882_, _22881_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22883_, _22843_, _22816_);
  or (_22884_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22885_, \oc8051_symbolic_cxrom1.regvalid [0], _16467_);
  and (_22886_, _22885_, _22809_);
  and (_22887_, _22886_, _22884_);
  or (_22888_, _22887_, _22883_);
  and (_22889_, _22888_, _22882_);
  and (_22890_, _22889_, _22872_);
  or (_22891_, _22890_, _22863_);
  or (_22892_, _22888_, _22881_);
  and (_22893_, _22892_, _16455_);
  and (_22894_, _22893_, _22891_);
  and (_22895_, _22894_, _22836_);
  or (_22896_, \oc8051_symbolic_cxrom1.regvalid [2], _16459_);
  or (_22897_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22898_, _22897_, _22896_);
  or (_22899_, _22898_, _22823_);
  or (_22900_, \oc8051_symbolic_cxrom1.regvalid [10], _16459_);
  or (_22901_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_22902_, _22901_, _22900_);
  and (_22903_, _22902_, _22823_);
  nor (_22904_, _22903_, _22826_);
  and (_22905_, _22904_, _22899_);
  and (_22906_, _22823_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_22907_, _22841_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_22908_, _22907_, _22906_);
  and (_22909_, _22823_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_22910_, _22874_, _16459_);
  or (_22911_, _22910_, _22909_);
  and (_22912_, _22911_, _22826_);
  and (_22913_, _22912_, _22908_);
  or (_22914_, _22913_, _22905_);
  or (_22915_, _22850_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_22916_, \oc8051_symbolic_cxrom1.regvalid [14], _16467_);
  and (_22917_, _22916_, _22915_);
  or (_22918_, _22917_, _22858_);
  nand (_22919_, _22850_, _19195_);
  or (_22920_, _22850_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_22921_, _22920_, _22919_);
  or (_22922_, _22921_, _22854_);
  and (_22923_, _22922_, _22918_);
  or (_22924_, _22923_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_22925_, _22850_, _18931_);
  and (_22926_, _22850_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_22927_, _22926_, _22925_);
  and (_22928_, _22927_, _22858_);
  or (_22929_, _22850_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_22930_, \oc8051_symbolic_cxrom1.regvalid [12], _16467_);
  and (_22931_, _22930_, _22854_);
  and (_22932_, _22931_, _22929_);
  or (_22933_, _22932_, _16459_);
  or (_22934_, _22933_, _22928_);
  or (_22935_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22936_, _22935_, _22865_);
  or (_22937_, _22936_, _16463_);
  or (_22938_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22939_, \oc8051_symbolic_cxrom1.regvalid [11], _16467_);
  and (_22940_, _22939_, _22938_);
  or (_22941_, _22940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_22942_, _22941_, _22937_);
  and (_22943_, _22942_, _22852_);
  and (_22944_, _16459_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_22945_, _22815_, _16463_);
  or (_22946_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22947_, \oc8051_symbolic_cxrom1.regvalid [9], _16467_);
  and (_22948_, _22947_, _22946_);
  or (_22949_, _22948_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_22950_, _22949_, _22945_);
  and (_22951_, _22950_, _22944_);
  or (_22952_, _22951_, _22943_);
  and (_22953_, _22942_, _16459_);
  or (_22954_, _22953_, _22818_);
  and (_22955_, _22954_, _22952_);
  and (_22956_, _22955_, _22934_);
  and (_22957_, _22956_, _22924_);
  and (_22958_, _22957_, _22914_);
  or (_22959_, _22958_, _22895_);
  nor (_22960_, _21863_, _16523_);
  and (_22961_, _22960_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22962_, _22960_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22963_, _22962_, _22961_);
  nand (_22964_, _22963_, _18879_);
  and (_22965_, _21876_, _16519_);
  nor (_22966_, _22965_, _22960_);
  and (_22967_, _22966_, _22526_);
  and (_22968_, _22967_, _22964_);
  not (_22969_, _22966_);
  and (_22970_, _22963_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_22971_, _22963_, _18865_);
  or (_22972_, _22971_, _22970_);
  and (_22973_, _22972_, _22969_);
  or (_22974_, _22973_, _22968_);
  and (_22975_, _22974_, _21863_);
  nand (_22976_, _22963_, _18887_);
  nor (_22977_, _22969_, _22540_);
  and (_22978_, _22977_, _22976_);
  and (_22979_, _22963_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_22980_, _22963_, _18894_);
  or (_22981_, _22980_, _22979_);
  and (_22982_, _22981_, _22969_);
  or (_22983_, _22982_, _22978_);
  and (_22984_, _22983_, _21888_);
  or (_22985_, _22984_, _22975_);
  or (_22986_, _22963_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_22987_, _22966_, _22508_);
  and (_22988_, _22987_, _22986_);
  and (_22989_, _22963_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_22990_, _22963_, _18906_);
  or (_22991_, _22990_, _22989_);
  and (_22992_, _22991_, _22969_);
  or (_22993_, _22992_, _22988_);
  and (_22994_, _22993_, _21902_);
  or (_22995_, _22963_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_22996_, _22969_, _22502_);
  and (_22997_, _22996_, _22995_);
  and (_22998_, _22963_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_22999_, _22963_, _18931_);
  or (_23000_, _22999_, _22998_);
  and (_23001_, _23000_, _22969_);
  or (_23002_, _23001_, _22997_);
  and (_23003_, _23002_, _21915_);
  or (_23004_, _23003_, _22994_);
  or (_23005_, _23004_, _22985_);
  nor (_23006_, _22516_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_23007_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_23008_, \oc8051_symbolic_cxrom1.regvalid [0], _16527_);
  and (_23009_, _23008_, _21846_);
  and (_23010_, _23009_, _23007_);
  and (_23011_, _22504_, _21872_);
  or (_23012_, _23011_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_23013_, _23012_, _23010_);
  or (_23014_, _23013_, _23006_);
  nor (_23015_, _22534_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_23016_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_23017_, \oc8051_symbolic_cxrom1.regvalid [1], _16527_);
  and (_23018_, _23017_, _21846_);
  and (_23019_, _23018_, _23016_);
  and (_23020_, _22542_, _21872_);
  or (_23021_, _23020_, _16515_);
  or (_23022_, _23021_, _23019_);
  or (_23023_, _23022_, _23015_);
  and (_23024_, _23023_, _23014_);
  and (_23025_, pc_log_change, _21842_);
  and (_23026_, _23025_, _22547_);
  nand (_23027_, _23026_, _23024_);
  nor (_23028_, _23027_, _21928_);
  and (_23029_, _23028_, _23005_);
  and (_23030_, _23029_, _22959_);
  nor (_23031_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23032_, _21193_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23033_, _23032_, _23031_);
  and (_23034_, _23033_, _21872_);
  nor (_23035_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23036_, _19871_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23037_, _23036_, _23035_);
  and (_23038_, _23037_, _21873_);
  nor (_23039_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23040_, _21203_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23041_, _23040_, _23039_);
  and (_23042_, _23041_, _22518_);
  nor (_23043_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23044_, _20076_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23045_, _23044_, _23043_);
  and (_23046_, _23045_, _21846_);
  or (_23047_, _23046_, _23042_);
  or (_23048_, _23047_, _23038_);
  or (_23049_, _23048_, _23034_);
  and (_23050_, _23049_, _16527_);
  nor (_23051_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23052_, _20490_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23053_, _23052_, _23051_);
  and (_23054_, _23053_, _21872_);
  nor (_23055_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23056_, _20694_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23057_, _23056_, _23055_);
  and (_23058_, _23057_, _21873_);
  nor (_23059_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23060_, _20286_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23061_, _23060_, _23059_);
  and (_23062_, _23061_, _22518_);
  nor (_23063_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23064_, _21211_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23065_, _23064_, _23063_);
  and (_23066_, _23065_, _21846_);
  or (_23067_, _23066_, _23062_);
  or (_23068_, _23067_, _23058_);
  or (_23069_, _23068_, _23054_);
  and (_23070_, _23069_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_23071_, _23070_, _23050_);
  and (_23072_, _23071_, _22547_);
  nor (_23073_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23074_, _18740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23075_, _23074_, _23073_);
  and (_23076_, _23075_, _22518_);
  nor (_23077_, _23076_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_23078_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23079_, _18716_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23080_, _23079_, _23078_);
  and (_23081_, _23080_, _21873_);
  not (_23082_, _23081_);
  nor (_23083_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23084_, _18735_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23085_, _23084_, _23083_);
  and (_23086_, _23085_, _21872_);
  nor (_23087_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23088_, _18695_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23089_, _23088_, _23087_);
  and (_23090_, _23089_, _21846_);
  nor (_23091_, _23090_, _23086_);
  and (_23092_, _23091_, _23082_);
  and (_23093_, _23092_, _23077_);
  nor (_23094_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23095_, _18728_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23096_, _23095_, _23094_);
  and (_23097_, _23096_, _22518_);
  nor (_23098_, _23097_, _16527_);
  nor (_23099_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23100_, _18711_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23101_, _23100_, _23099_);
  and (_23102_, _23101_, _21873_);
  not (_23103_, _23102_);
  nor (_23104_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23105_, _18723_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23106_, _23105_, _23104_);
  and (_23107_, _23106_, _21872_);
  nor (_23108_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23109_, _18703_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23110_, _23109_, _23108_);
  and (_23111_, _23110_, _21846_);
  nor (_23112_, _23111_, _23107_);
  and (_23113_, _23112_, _23103_);
  and (_23114_, _23113_, _23098_);
  nor (_23115_, _23114_, _23093_);
  not (_23116_, _23115_);
  and (_23117_, _23116_, _23072_);
  and (_23118_, _23117_, _23030_);
  and (_23119_, _23118_, _22807_);
  and (property_invalid_jnc, _23119_, _22501_);
  and (_23120_, _21861_, _22354_);
  nor (_23121_, _22348_, _22354_);
  nor (_23122_, _23121_, _23120_);
  nor (_23123_, _23122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_23124_, _23122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_23125_, _21969_, _22354_);
  and (_23126_, _22356_, cy_reg);
  nor (_23127_, _23126_, _23125_);
  nor (_23128_, _23127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_23129_, _23127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_23130_, _21975_, _22354_);
  nor (_23131_, _22364_, _22354_);
  nor (_23132_, _23131_, _23130_);
  and (_23133_, _23132_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_23134_, _23132_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_23135_, _21980_, cy_reg);
  nor (_23136_, _22371_, _22354_);
  nor (_23137_, _23136_, _23135_);
  nor (_23138_, _23137_, _16503_);
  and (_23139_, _23137_, _16503_);
  and (_23140_, _21985_, _22354_);
  nor (_23141_, _22381_, _22354_);
  nor (_23142_, _23141_, _23140_);
  and (_23143_, _23142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_23144_, _23142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_23145_, _21997_, _22354_);
  nor (_23146_, _22389_, _22354_);
  nor (_23147_, _23146_, _23145_);
  nor (_23148_, _23147_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_23149_, _23147_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_23150_, _22000_, _22354_);
  and (_23151_, _22405_, cy_reg);
  nor (_23152_, _23151_, _23150_);
  and (_23153_, _23152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_23154_, _23152_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_23155_, _22007_, cy_reg);
  nor (_23156_, _22412_, _22354_);
  nor (_23157_, _23156_, _23155_);
  nor (_23158_, _23157_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_23159_, _23157_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_23160_, _22051_, _22354_);
  and (_23161_, _22421_, cy_reg);
  nor (_23162_, _23161_, _23160_);
  nor (_23163_, _23162_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_23164_, _23162_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_23165_, _22096_, _22354_);
  and (_23166_, _22427_, cy_reg);
  nor (_23167_, _23166_, _23165_);
  nor (_23168_, _23167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_23169_, _23167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_23170_, _22140_, _22354_);
  and (_23171_, _22435_, cy_reg);
  nor (_23172_, _23171_, _23170_);
  nor (_23173_, _23172_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_23174_, _23172_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_23175_, _21868_, cy_reg);
  and (_23176_, _22441_, cy_reg);
  nor (_23177_, _23176_, _23175_);
  nor (_23178_, _23177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_23179_, _23177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_23180_, _22465_, cy_reg);
  nor (_23181_, _21874_, cy_reg);
  nor (_23182_, _23181_, _23180_);
  nor (_23183_, _23182_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_23184_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_23185_, _22449_, cy_reg);
  nor (_23186_, _23185_, _23184_);
  and (_23187_, _23186_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_23188_, _22456_, _22301_);
  or (_23189_, _23188_, _22458_);
  or (_23190_, _23189_, _22354_);
  nand (_23191_, _22456_, _22354_);
  and (_23192_, _23191_, _23190_);
  nor (_23193_, _23186_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_23194_, _23193_, _23192_);
  or (_23195_, _23194_, _23187_);
  and (_23196_, _23182_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_23197_, _23196_, _23195_);
  or (_23198_, _23197_, _23183_);
  or (_23199_, _23198_, _23179_);
  or (_23200_, _23199_, _23178_);
  or (_23201_, _23200_, _23174_);
  or (_23202_, _23201_, _23173_);
  or (_23203_, _23202_, _23169_);
  or (_23204_, _23203_, _23168_);
  or (_23205_, _23204_, _23164_);
  or (_23206_, _23205_, _23163_);
  or (_23207_, _23206_, _23159_);
  or (_23208_, _23207_, _23158_);
  or (_23209_, _23208_, _23154_);
  or (_23210_, _23209_, _23153_);
  or (_23211_, _23210_, _23149_);
  or (_23212_, _23211_, _23148_);
  and (_23213_, _21991_, _22354_);
  and (_23214_, _22485_, cy_reg);
  nor (_23215_, _23214_, _23213_);
  and (_23216_, _23215_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_23217_, _23215_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_23218_, _23217_, _23216_);
  or (_23219_, _23218_, _23212_);
  or (_23220_, _23219_, _23144_);
  or (_23221_, _23220_, _23143_);
  or (_23222_, _23221_, _23139_);
  or (_23223_, _23222_, _23138_);
  or (_23224_, _23223_, _23134_);
  or (_23225_, _23224_, _23133_);
  or (_23226_, _23225_, _23129_);
  or (_23227_, _23226_, _23128_);
  or (_23228_, _23227_, _23124_);
  or (_23229_, _23228_, _23123_);
  nor (_23230_, _22804_, _22762_);
  and (_23231_, _23230_, _22720_);
  and (_23232_, _23231_, _23118_);
  and (property_invalid_jc, _23232_, _23229_);
  or (_23233_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_23234_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_23235_, _23234_, _23233_);
  or (_23236_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_23237_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_23238_, _23237_, _23236_);
  or (_23239_, _23238_, _23235_);
  nor (_23240_, _22301_, _16455_);
  or (_23241_, _21861_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_23242_, _21861_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_23243_, _23242_, _23241_);
  nor (_23244_, _21975_, _16507_);
  and (_23245_, _21975_, _16507_);
  or (_23246_, _23245_, _23244_);
  or (_23247_, _21980_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_23248_, _21980_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_23249_, _23248_, _23247_);
  or (_23250_, _23249_, _23246_);
  or (_23251_, _21969_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_23252_, _21969_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_23253_, _23252_, _23251_);
  or (_23254_, _23253_, _23250_);
  or (_23255_, _23254_, _23243_);
  or (_23256_, _23255_, _23240_);
  and (_23257_, _22301_, _16455_);
  nor (_23258_, _22223_, _16463_);
  or (_23259_, _23258_, _23257_);
  or (_23260_, _23259_, _23256_);
  or (_23261_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_23262_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_23263_, _23262_, _23261_);
  and (_23264_, _22804_, _16487_);
  nor (_23265_, _22804_, _16487_);
  or (_23266_, _23265_, _23264_);
  and (_23267_, _23072_, _16491_);
  nor (_23268_, _23072_, _16491_);
  or (_23269_, _23268_, _23267_);
  or (_23270_, _23269_, _23266_);
  nor (_23271_, _21985_, _16499_);
  and (_23272_, _21985_, _16499_);
  or (_23273_, _23272_, _23271_);
  and (_23274_, _23115_, _22547_);
  nor (_23275_, _23274_, _16495_);
  and (_23276_, _23274_, _16495_);
  or (_23277_, _23276_, _23275_);
  or (_23278_, _23277_, _23273_);
  or (_23279_, _23278_, _23270_);
  or (_23280_, _23279_, _23263_);
  or (_23281_, _23280_, _23260_);
  and (_23282_, _22048_, _16479_);
  and (_23283_, _21967_, _16483_);
  nor (_23284_, _21967_, _16483_);
  or (_23285_, _23284_, _23283_);
  or (_23286_, _23285_, _23282_);
  and (_23287_, _22138_, _16471_);
  nor (_23288_, _22048_, _16479_);
  or (_23289_, _23288_, _23287_);
  and (_23290_, _22223_, _16463_);
  nor (_23291_, _22138_, _16471_);
  or (_23292_, _23291_, _23290_);
  or (_23293_, _23292_, _23289_);
  or (_23294_, _23293_, _23286_);
  or (_23295_, _23294_, _23281_);
  or (_23296_, _23295_, _23239_);
  not (_23297_, _22673_);
  and (_23298_, _22718_, _22632_);
  and (_23299_, _23298_, _23297_);
  and (_23300_, _23299_, _23030_);
  and (property_invalid_ajmp, _23300_, _23296_);
  and (_23301_, _22691_, _21873_);
  and (_23302_, _22677_, _21872_);
  or (_23303_, _23302_, _23301_);
  and (_23304_, _22686_, _22518_);
  and (_23305_, _22682_, _21846_);
  or (_23306_, _23305_, _23304_);
  or (_23307_, _23306_, _23303_);
  and (_23308_, _23307_, _22142_);
  and (_23309_, _22712_, _21873_);
  and (_23310_, _22698_, _21872_);
  or (_23311_, _23310_, _23309_);
  and (_23312_, _22707_, _22518_);
  and (_23313_, _22703_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_23314_, _23313_, _23312_);
  or (_23315_, _23314_, _23311_);
  and (_23316_, _23315_, _21868_);
  or (_23317_, _23316_, _23308_);
  and (_23318_, _23317_, _23024_);
  and (_23319_, _23318_, _16455_);
  nor (_23320_, _23318_, _16455_);
  or (_23321_, _23320_, _23319_);
  and (_23322_, _22647_, _21873_);
  or (_23323_, _23322_, _22142_);
  and (_23324_, _22643_, _21846_);
  and (_23325_, _22635_, _22518_);
  and (_23326_, _22639_, _21872_);
  or (_23327_, _23326_, _23325_);
  or (_23328_, _23327_, _23324_);
  or (_23329_, _23328_, _23323_);
  and (_23330_, _22663_, _21846_);
  or (_23331_, _23330_, _21868_);
  and (_23332_, _22659_, _21872_);
  and (_23333_, _22655_, _22518_);
  and (_23334_, _22667_, _21873_);
  or (_23335_, _23334_, _23333_);
  or (_23336_, _23335_, _23332_);
  or (_23337_, _23336_, _23331_);
  and (_23338_, _23337_, _23329_);
  and (_23339_, _23338_, _23024_);
  nor (_23340_, _23339_, _16459_);
  and (_23341_, _23339_, _16459_);
  or (_23342_, _23341_, _23340_);
  or (_23343_, _23342_, _23321_);
  and (_23344_, _22562_, _21873_);
  or (_23345_, _23344_, _22142_);
  and (_23346_, _22558_, _21846_);
  and (_23347_, _22550_, _22518_);
  and (_23348_, _22554_, _21872_);
  or (_23349_, _23348_, _23347_);
  or (_23350_, _23349_, _23346_);
  or (_23351_, _23350_, _23345_);
  and (_23352_, _22578_, _21846_);
  or (_23353_, _23352_, _21868_);
  and (_23354_, _22574_, _21872_);
  and (_23355_, _22570_, _22518_);
  and (_23356_, _22582_, _21873_);
  or (_23357_, _23356_, _23355_);
  or (_23358_, _23357_, _23354_);
  or (_23359_, _23358_, _23353_);
  and (_23360_, _23359_, _23351_);
  and (_23361_, _23360_, _23024_);
  nand (_23362_, _23361_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_23363_, _23361_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_23364_, _23363_, _23362_);
  and (_23365_, _22604_, _21873_);
  or (_23366_, _23365_, _22142_);
  and (_23367_, _22600_, _21846_);
  and (_23368_, _22592_, _22518_);
  and (_23369_, _22596_, _21872_);
  or (_23370_, _23369_, _23368_);
  or (_23371_, _23370_, _23367_);
  or (_23372_, _23371_, _23366_);
  and (_23373_, _22620_, _21846_);
  or (_23374_, _23373_, _21868_);
  and (_23375_, _22616_, _21872_);
  and (_23376_, _22612_, _22518_);
  and (_23377_, _22624_, _21873_);
  or (_23378_, _23377_, _23376_);
  or (_23379_, _23378_, _23375_);
  or (_23380_, _23379_, _23374_);
  and (_23381_, _23380_, _23372_);
  and (_23382_, _23381_, _23024_);
  nand (_23383_, _23382_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_23384_, _23382_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_23385_, _23384_, _23383_);
  or (_23386_, _23385_, _23364_);
  or (_23387_, _23386_, _23343_);
  and (_23388_, _22727_, _21872_);
  or (_23389_, _23388_, _22142_);
  and (_23390_, _22723_, _22518_);
  and (_23391_, _22731_, _21846_);
  or (_23392_, _23391_, _23390_);
  and (_23393_, _22735_, _21873_);
  or (_23394_, _23393_, _23392_);
  or (_23395_, _23394_, _23389_);
  and (_23396_, _22751_, _21846_);
  or (_23397_, _23396_, _21868_);
  and (_23398_, _22747_, _21872_);
  and (_23399_, _22743_, _22518_);
  and (_23400_, _22755_, _21873_);
  or (_23401_, _23400_, _23399_);
  or (_23402_, _23401_, _23398_);
  or (_23403_, _23402_, _23397_);
  and (_23404_, _23403_, _23395_);
  and (_23405_, _23404_, _23024_);
  or (_23406_, _23405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_23407_, _23405_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_23408_, _23407_, _23406_);
  and (_23409_, _22789_, _21872_);
  or (_23410_, _23409_, _21868_);
  and (_23411_, _22785_, _22518_);
  and (_23412_, _22793_, _21846_);
  or (_23413_, _23412_, _23411_);
  and (_23414_, _22797_, _21873_);
  or (_23415_, _23414_, _23413_);
  or (_23416_, _23415_, _23410_);
  and (_23417_, _22773_, _21846_);
  or (_23418_, _23417_, _22142_);
  and (_23419_, _22769_, _21872_);
  and (_23420_, _22765_, _22518_);
  and (_23421_, _22777_, _21873_);
  or (_23422_, _23421_, _23420_);
  or (_23423_, _23422_, _23419_);
  or (_23424_, _23423_, _23418_);
  and (_23425_, _23424_, _23416_);
  and (_23426_, _23425_, _23024_);
  nor (_23427_, _23426_, _16475_);
  and (_23428_, _23426_, _16475_);
  or (_23429_, _23428_, _23427_);
  or (_23430_, _23429_, _23408_);
  and (_23431_, _23080_, _21872_);
  or (_23432_, _23431_, _22142_);
  and (_23433_, _23075_, _21846_);
  and (_23434_, _23085_, _22518_);
  or (_23435_, _23434_, _23433_);
  and (_23436_, _23089_, _21873_);
  or (_23437_, _23436_, _23435_);
  or (_23438_, _23437_, _23432_);
  and (_23439_, _23101_, _21872_);
  or (_23440_, _23439_, _21868_);
  and (_23441_, _23096_, _21846_);
  and (_23442_, _23106_, _22518_);
  and (_23443_, _23110_, _21873_);
  or (_23444_, _23443_, _23442_);
  or (_23445_, _23444_, _23441_);
  or (_23446_, _23445_, _23440_);
  and (_23447_, _23446_, _23438_);
  and (_23448_, _23447_, _23024_);
  nand (_23449_, _23448_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_23450_, _23448_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_23451_, _23450_, _23449_);
  and (_23452_, _23045_, _21873_);
  or (_23453_, _23452_, _22142_);
  and (_23454_, _23041_, _21846_);
  and (_23455_, _23033_, _22518_);
  and (_23456_, _23037_, _21872_);
  or (_23457_, _23456_, _23455_);
  or (_23458_, _23457_, _23454_);
  or (_23459_, _23458_, _23453_);
  and (_23460_, _23061_, _21846_);
  or (_23461_, _23460_, _21868_);
  and (_23462_, _23057_, _21872_);
  and (_23463_, _23053_, _22518_);
  and (_23464_, _23065_, _21873_);
  or (_23465_, _23464_, _23463_);
  or (_23466_, _23465_, _23462_);
  or (_23467_, _23466_, _23461_);
  and (_23468_, _23467_, _23459_);
  and (_23469_, _23468_, _23024_);
  nor (_23470_, _23469_, _16479_);
  and (_23471_, _23469_, _16479_);
  or (_23472_, _23471_, _23470_);
  or (_23473_, _23472_, _23451_);
  or (_23474_, _23473_, _23430_);
  or (_23475_, _23474_, _23387_);
  or (_23476_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_23477_, _22262_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_23478_, _23477_, _23476_);
  and (_23479_, _22301_, _16487_);
  nor (_23480_, _22301_, _16487_);
  or (_23481_, _23480_, _23479_);
  or (_23482_, _23481_, _23478_);
  or (_23483_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_23484_, _22180_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_23485_, _23484_, _23483_);
  nor (_23486_, _22223_, _16495_);
  and (_23487_, _22223_, _16495_);
  or (_23488_, _23487_, _23486_);
  or (_23489_, _23488_, _23485_);
  or (_23490_, _23489_, _23482_);
  or (_23491_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_23492_, _22093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_23493_, _23492_, _23491_);
  nor (_23494_, _22138_, _16503_);
  and (_23495_, _22138_, _16503_);
  or (_23496_, _23495_, _23494_);
  or (_23497_, _23496_, _23493_);
  nor (_23498_, _21967_, _15859_);
  and (_23499_, _21967_, _15859_);
  or (_23500_, _23499_, _23498_);
  and (_23501_, _22048_, _16511_);
  nor (_23502_, _22048_, _16511_);
  or (_23503_, _23502_, _23501_);
  or (_23504_, _23503_, _23500_);
  or (_23505_, _23504_, _23497_);
  or (_23506_, _23505_, _23490_);
  or (_23507_, _23506_, _23475_);
  nor (_23508_, _23274_, _23072_);
  not (_23509_, _22718_);
  and (_23510_, _23509_, _22632_);
  and (_23511_, _22805_, _23510_);
  and (_23512_, _23511_, _22674_);
  and (_23513_, _23512_, _23508_);
  and (_23514_, _23513_, _23030_);
  and (property_invalid_ljmp, _23514_, _23507_);
  and (_23515_, _22348_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_23516_, _22348_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  or (_23517_, _22356_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_23518_, _22356_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_23519_, _23518_, _23517_);
  or (_23520_, _22364_, _16507_);
  nand (_23521_, _22364_, _16507_);
  and (_23522_, _23521_, _23520_);
  or (_23523_, _22371_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_23524_, _22371_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_23525_, _23524_, _23523_);
  and (_23526_, _22381_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_23527_, _22381_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_23528_, _22389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_23529_, _22389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_23531_, _22421_, _16479_);
  nor (_23532_, _22421_, _16479_);
  nor (_23533_, _22427_, _16475_);
  and (_23534_, _22427_, _16475_);
  and (_23535_, _22435_, _16471_);
  nor (_23536_, _22435_, _16471_);
  and (_23537_, _22441_, _16467_);
  nor (_23538_, _22441_, _16467_);
  and (_23539_, _22465_, _16463_);
  or (_23540_, _22449_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_23541_, _22449_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_23542_, _23541_, _23540_);
  or (_23543_, _23542_, _23189_);
  nor (_23544_, _22465_, _16463_);
  or (_23545_, _23544_, _23543_);
  or (_23546_, _23545_, _23539_);
  or (_23547_, _23546_, _23538_);
  or (_23548_, _23547_, _23537_);
  or (_23549_, _23548_, _23536_);
  or (_23550_, _23549_, _23535_);
  or (_23551_, _23550_, _23534_);
  or (_23552_, _23551_, _23533_);
  or (_23553_, _23552_, _23532_);
  or (_23554_, _23553_, _23531_);
  or (_23555_, _23554_, _22415_);
  or (_23556_, _23555_, _22408_);
  or (_23557_, _23556_, _23529_);
  or (_23558_, _23557_, _23528_);
  nor (_23559_, _22485_, _16495_);
  and (_23560_, _22485_, _16495_);
  or (_23561_, _23560_, _23559_);
  or (_23562_, _23561_, _23558_);
  or (_23563_, _23562_, _23527_);
  or (_23564_, _23563_, _23526_);
  or (_23565_, _23564_, _23525_);
  or (_23566_, _23565_, _23522_);
  or (_23567_, _23566_, _23519_);
  or (_23568_, _23567_, _23516_);
  or (_23569_, _23568_, _23515_);
  not (_23570_, _23072_);
  and (_23571_, _23274_, _23570_);
  and (_23572_, _23571_, _23230_);
  and (_23573_, _23572_, _22720_);
  and (_23574_, _23573_, _23030_);
  and (property_invalid_sjmp, _23574_, _23569_);
  and (_23575_, _22961_, _21850_);
  and (_23576_, _23575_, _21854_);
  and (_23577_, _23576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_23578_, _23577_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_23579_, _23578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_23580_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_23581_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_23582_, _23581_, _23580_);
  not (_23583_, _23582_);
  nor (_23584_, _23583_, _23579_);
  and (_23585_, _23583_, _23579_);
  not (_23586_, _23577_);
  nor (_23587_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_23588_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_23589_, _23588_, _23587_);
  nor (_23590_, _23589_, _23586_);
  and (_23591_, _23575_, _21852_);
  and (_23592_, _23575_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_23593_, _23592_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_23594_, _23593_, _23591_);
  and (_23595_, _23594_, _16491_);
  and (_23596_, _22961_, _21849_);
  and (_23597_, _22961_, _21848_);
  nor (_23598_, _23597_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_23599_, _23598_, _23596_);
  nor (_23600_, _23599_, _16479_);
  or (_23601_, _23600_, _23595_);
  nor (_23602_, _23594_, _16491_);
  and (_23603_, _23599_, _16479_);
  or (_23604_, _23603_, _23602_);
  or (_23605_, _23604_, _23601_);
  or (_23606_, _23605_, _23590_);
  nor (_23607_, _23596_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_23608_, _23607_, _23575_);
  nand (_23609_, _23608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_23610_, _23608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_23611_, _23610_, _23609_);
  and (_23612_, _23589_, _23586_);
  or (_23613_, _23612_, _23611_);
  or (_23614_, _23613_, _23606_);
  or (_23615_, _23614_, _23585_);
  or (_23616_, _23615_, _23584_);
  nor (_23617_, _23578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_23618_, _23617_, _23579_);
  and (_23619_, _23618_, _16511_);
  nor (_23620_, _23618_, _16511_);
  nor (_23621_, _23576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_23622_, _23621_, _23577_);
  and (_23623_, _23622_, _16503_);
  nor (_23624_, _23622_, _16503_);
  and (_23625_, _23575_, _21853_);
  nor (_23626_, _23591_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_23627_, _23626_, _23625_);
  and (_23628_, _23627_, _16495_);
  and (_23629_, _22961_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_23630_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_23631_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_23632_, _23631_, _23630_);
  not (_23633_, _23632_);
  nor (_23634_, _23633_, _23629_);
  and (_23635_, _22963_, _16467_);
  and (_23636_, _23633_, _23629_);
  or (_23637_, _23636_, _23635_);
  or (_23638_, _23637_, _23634_);
  and (_23639_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_23640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_23641_, _23640_, _23639_);
  nand (_23642_, _23641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_23643_, _23641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23644_, _23643_, _23642_);
  nand (_23645_, _22966_, _16463_);
  nand (_23646_, _23645_, _23644_);
  nor (_23647_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_23648_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_23649_, _23648_, _23647_);
  not (_23650_, _23649_);
  nor (_23651_, _23650_, _22961_);
  nor (_23652_, _22966_, _16463_);
  or (_23653_, _23652_, _23651_);
  or (_23654_, _23653_, _23646_);
  nor (_23655_, _22963_, _16467_);
  and (_23656_, _23650_, _22961_);
  or (_23657_, _23656_, _22456_);
  or (_23658_, _23657_, _23655_);
  or (_23659_, _23658_, _23654_);
  or (_23660_, _23659_, _23638_);
  nor (_23661_, _23575_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_23662_, _23661_, _23592_);
  nor (_23663_, _23662_, _16487_);
  and (_23664_, _23662_, _16487_);
  or (_23665_, _23664_, _23663_);
  or (_23666_, _23665_, _23660_);
  or (_23667_, _23666_, _23628_);
  nor (_23668_, _23627_, _16495_);
  nor (_23669_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_23670_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_23671_, _23670_, _23669_);
  or (_23672_, _23671_, _23625_);
  nand (_23673_, _23671_, _23625_);
  and (_23674_, _23673_, _23672_);
  or (_23675_, _23674_, _23668_);
  or (_23676_, _23675_, _23667_);
  or (_23677_, _23676_, _23624_);
  or (_23678_, _23677_, _23623_);
  or (_23679_, _23678_, _23620_);
  or (_23680_, _23679_, _23619_);
  or (_23681_, _23680_, _23616_);
  not (_23682_, _22762_);
  nor (_23683_, _22673_, _22588_);
  and (_23684_, _23683_, _22631_);
  and (_23685_, _23684_, _22718_);
  and (_23686_, _23685_, _23682_);
  and (_23687_, _23686_, _22805_);
  or (_23688_, _23687_, _22807_);
  and (_23689_, _23688_, _23571_);
  and (_23690_, _23685_, _22804_);
  and (_23691_, _23690_, _22762_);
  and (_23692_, _23298_, _22673_);
  nand (_23693_, _22804_, _22761_);
  and (_23694_, _23693_, _23692_);
  or (_23695_, _23694_, _23691_);
  and (_23696_, _23695_, _23117_);
  or (_23697_, _23696_, _23689_);
  and (_23698_, _23697_, _23030_);
  and (property_invalid_pcp3, _23698_, _23681_);
  not (_23699_, _22717_);
  and (_23700_, _23684_, _23699_);
  and (_23701_, _22674_, _22631_);
  and (_23702_, _23701_, _22762_);
  and (_23703_, _23702_, _22804_);
  or (_23704_, _23703_, _23700_);
  and (_23705_, _23704_, _23116_);
  or (_23706_, _23705_, _23686_);
  and (_23707_, _23706_, _23072_);
  or (_23708_, _23512_, _23072_);
  or (_23709_, _23690_, _23511_);
  and (_23710_, _23709_, _23274_);
  and (_23711_, _23710_, _23708_);
  and (_23712_, _23684_, _22806_);
  not (_23713_, _22761_);
  or (_23714_, _23701_, _22589_);
  and (_23715_, _23714_, _23713_);
  or (_23716_, _23715_, _23712_);
  and (_23717_, _23716_, _23571_);
  not (_23718_, _23274_);
  and (_23719_, _23685_, _22805_);
  and (_23720_, _23071_, _22588_);
  and (_23721_, _23720_, _22804_);
  and (_23722_, _23721_, _22761_);
  or (_23723_, _23722_, _23719_);
  and (_23724_, _23723_, _23718_);
  and (_23725_, _23571_, _22803_);
  and (_23726_, _23117_, _22674_);
  or (_23727_, _23726_, _23725_);
  and (_23728_, _23727_, _23510_);
  and (_23729_, _23508_, _22804_);
  and (_23730_, _23729_, _23684_);
  or (_23731_, _23730_, _23728_);
  or (_23732_, _23731_, _23724_);
  or (_23733_, _23732_, _23717_);
  or (_23734_, _23733_, _23711_);
  or (_23735_, _23734_, _23707_);
  and (_23736_, _21997_, _16491_);
  or (_23737_, _22051_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_23738_, _22051_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_23739_, _23738_, _23737_);
  nor (_23740_, _21997_, _16491_);
  or (_23741_, _23740_, _23739_);
  or (_23742_, _23741_, _23736_);
  and (_23743_, _21874_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_23744_, _21874_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_23745_, _23744_, _23743_);
  or (_23746_, _23649_, _21847_);
  nand (_23747_, _23649_, _21847_);
  and (_23748_, _23747_, _23746_);
  nand (_23749_, _23641_, _22456_);
  or (_23750_, _23749_, _23748_);
  or (_23751_, _23750_, _23745_);
  or (_23752_, _23632_, _22094_);
  nand (_23753_, _23632_, _22094_);
  and (_23754_, _23753_, _23752_);
  or (_23755_, _21868_, _16467_);
  nand (_23756_, _21868_, _16467_);
  and (_23757_, _23756_, _23755_);
  or (_23758_, _23757_, _23754_);
  or (_23759_, _23758_, _23751_);
  or (_23760_, _23759_, _22401_);
  or (_23761_, _23760_, _22398_);
  or (_23762_, _23761_, _23273_);
  nor (_23763_, _21991_, _16495_);
  and (_23764_, _21991_, _16495_);
  or (_23765_, _23764_, _23763_);
  or (_23766_, _23765_, _23762_);
  or (_23767_, _23766_, _23742_);
  or (_23768_, _23767_, _23255_);
  and (_23769_, _23768_, _23030_);
  and (property_invalid_pcp2, _23769_, _23735_);
  and (_23770_, _22806_, _22588_);
  and (_23771_, _23230_, _22719_);
  and (_23772_, _23699_, _22631_);
  and (_23773_, _23772_, _22805_);
  or (_23774_, _23773_, _23771_);
  and (_23775_, _23774_, _23718_);
  and (_23776_, _23700_, _23230_);
  or (_23777_, _23776_, _23692_);
  or (_23778_, _23777_, _23775_);
  or (_23779_, _23778_, _23770_);
  and (_23780_, _23779_, _23570_);
  and (_23781_, _23115_, _23699_);
  and (_23782_, _23781_, _22804_);
  or (_23783_, _23782_, _23715_);
  and (_23784_, _22718_, _22674_);
  or (_23785_, _23772_, _23784_);
  nor (_23786_, _23116_, _22589_);
  and (_23787_, _23786_, _23785_);
  or (_23788_, _23787_, _23783_);
  and (_23789_, _23788_, _23072_);
  and (_23790_, _23684_, _23682_);
  and (_23791_, _23725_, _23790_);
  nor (_23792_, _23115_, _22803_);
  and (_23793_, _23792_, _22589_);
  and (_23794_, _23721_, _23274_);
  or (_23795_, _23794_, _23793_);
  or (_23796_, _23795_, _23791_);
  nor (_23797_, _22804_, _22589_);
  and (_23798_, _23797_, _23702_);
  and (_23799_, _23714_, _23508_);
  or (_23800_, _23799_, _23798_);
  or (_23801_, _23800_, _23796_);
  or (_23802_, _23801_, _23789_);
  or (_23803_, _23802_, _23780_);
  and (_23804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _16515_);
  and (_23805_, _21975_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23806_, _23805_, _23804_);
  nor (_23807_, _23806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_23808_, _21857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23809_, _23808_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_23810_, _23808_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_23811_, _23810_, _23809_);
  and (_23812_, _23811_, _16511_);
  and (_23813_, _23806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_23814_, _23813_, _23812_);
  or (_23815_, _23814_, _23807_);
  or (_23816_, _16547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_23817_, _21997_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23818_, _23817_, _23816_);
  and (_23819_, _23818_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_23820_, _23818_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_23821_, _21847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_23822_, _23821_, _21850_);
  and (_23823_, _23822_, _21853_);
  or (_23824_, _23823_, _23671_);
  nand (_23825_, _23823_, _23671_);
  and (_23826_, _23825_, _23824_);
  nor (_23827_, _21877_, _16463_);
  and (_23828_, _21877_, _16463_);
  or (_23829_, _23828_, _23827_);
  not (_23830_, _23822_);
  nor (_23831_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_23832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_23833_, _23832_, _23831_);
  nor (_23834_, _23833_, _23830_);
  and (_23835_, _23833_, _23830_);
  or (_23836_, _23835_, _23834_);
  or (_23837_, _23836_, _23829_);
  and (_23838_, _22004_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23839_, _23838_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_23840_, _23839_, _23822_);
  and (_23841_, _23840_, _16483_);
  nor (_23842_, _23821_, _23650_);
  and (_23843_, _23821_, _23650_);
  or (_23844_, _23843_, _22456_);
  or (_23845_, _23844_, _23842_);
  or (_23846_, _23845_, _23644_);
  or (_23847_, _23846_, _23841_);
  or (_23848_, _23847_, _23837_);
  or (_23849_, _23848_, _23826_);
  not (_23850_, _22050_);
  nor (_23851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23852_, _23851_, _23838_);
  and (_23853_, _23852_, _23850_);
  or (_23854_, _23853_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_23855_, _23853_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_23856_, _23855_, _23854_);
  nor (_23857_, _23840_, _16483_);
  nor (_23858_, _21870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_23859_, _21870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_23860_, _23859_, _23858_);
  or (_23861_, _23860_, _23857_);
  or (_23862_, _23861_, _23856_);
  or (_23863_, _23862_, _23849_);
  or (_23864_, _23863_, _23820_);
  or (_23865_, _23864_, _23819_);
  nor (_23866_, _23811_, _16511_);
  and (_23867_, _23822_, _21854_);
  and (_23868_, _23867_, _16558_);
  nor (_23869_, _23867_, _16558_);
  or (_23870_, _23869_, _23868_);
  nand (_23871_, _23870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_23872_, _23870_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_23873_, _23872_, _23871_);
  and (_23874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _16515_);
  and (_23875_, _22096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_23876_, _23875_, _23874_);
  or (_23877_, _23876_, _16475_);
  nand (_23878_, _23876_, _16475_);
  and (_23879_, _23878_, _23877_);
  or (_23880_, _23879_, _23873_);
  nor (_23881_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_23882_, _23881_, _23823_);
  nor (_23883_, _23882_, _21990_);
  nor (_23884_, _23883_, _16495_);
  and (_23885_, _23883_, _16495_);
  or (_23886_, _23885_, _23884_);
  or (_23887_, _23886_, _23880_);
  or (_23888_, _23887_, _23866_);
  or (_23889_, _23888_, _23865_);
  nor (_23890_, _23809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_23891_, _23809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_23892_, _23891_, _23890_);
  and (_23893_, _23892_, _15859_);
  nor (_23894_, _23892_, _15859_);
  or (_23895_, _23894_, _23893_);
  or (_23896_, _23895_, _23889_);
  or (_23897_, _23896_, _23815_);
  and (_23898_, _23897_, _23030_);
  and (property_invalid_pcp1, _23898_, _23803_);
  buf (_00587_, _27357_);
  buf (_02706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7]);
  buf (_10034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0]);
  buf (_10038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1]);
  buf (_10042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2]);
  buf (_10046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3]);
  buf (_10050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4]);
  buf (_10054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5]);
  buf (_10058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6]);
  buf (_24407_, _24307_);
  buf (_24409_, _24308_);
  buf (_24421_, _24307_);
  buf (_24422_, _24308_);
  buf (_24739_, _24328_);
  buf (_24740_, _24329_);
  buf (_24741_, _24330_);
  buf (_24743_, _24331_);
  buf (_24744_, _24333_);
  buf (_24745_, _24334_);
  buf (_24746_, _24335_);
  buf (_24747_, _24336_);
  buf (_24748_, _24337_);
  buf (_24749_, _24339_);
  buf (_24750_, _24340_);
  buf (_24751_, _24341_);
  buf (_24752_, _24342_);
  buf (_24754_, _24343_);
  buf (_24805_, _24328_);
  buf (_24806_, _24329_);
  buf (_24807_, _24330_);
  buf (_24809_, _24331_);
  buf (_24810_, _24333_);
  buf (_24811_, _24334_);
  buf (_24812_, _24335_);
  buf (_24813_, _24336_);
  buf (_24814_, _24337_);
  buf (_24815_, _24339_);
  buf (_24816_, _24340_);
  buf (_24817_, _24341_);
  buf (_24818_, _24342_);
  buf (_24820_, _24343_);
  buf (_25393_, _25154_);
  buf (_25569_, _25154_);
  dff (cy_reg, _00000_);
  dff (pc_log_change_r, pc_log_change);
  dff (first_instr, _00001_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _28202_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _28202_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _28202_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _28202_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _28202_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _28202_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _28202_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _28202_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _25625_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _25629_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _25634_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _25640_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _25647_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _25655_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _25663_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _25673_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _25683_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _28201_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _28201_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _28201_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _28201_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _28201_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _28201_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _25618_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _28209_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _28209_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _28209_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _28209_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _28209_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _28209_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _28209_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _28209_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _28210_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _28210_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _28210_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _28210_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _28210_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _28210_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _28210_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _28210_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _28211_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _28211_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _28211_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _28211_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _28211_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _28211_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _28211_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _28211_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _28212_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _28212_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _28212_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _28212_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _28212_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _28212_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _28212_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _28212_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _28213_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _28213_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _28213_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _28213_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _28213_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _28213_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _28213_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _28213_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _28214_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _28214_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _28214_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _28214_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _28214_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _28214_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _28214_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _28214_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _28215_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _28215_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _28215_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _28215_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _28215_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _28215_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _28215_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _28215_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _28216_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _28216_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _28216_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _28216_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _28216_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _28216_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _28216_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _28216_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _28217_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _28217_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _28217_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _28217_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _28217_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _28217_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _28217_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _28217_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _28203_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _28203_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _28203_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _28203_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _28203_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _28203_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _28203_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _28203_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _28204_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _28204_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _28204_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _28204_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _28204_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _28204_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _28204_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _28204_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _28205_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _28205_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _28205_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _28205_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _28205_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _28205_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _28205_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _28205_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _28206_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _28206_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _28206_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _28206_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _28206_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _28206_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _28206_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _28206_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _28207_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _28207_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _28207_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _28207_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _28207_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _28207_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _28207_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _28207_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _28208_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _28208_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _28208_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _28208_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _28208_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _28208_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _28208_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _25622_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03039_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03049_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03068_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03084_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03100_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00985_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03108_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00958_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03117_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03125_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03132_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03141_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03149_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03158_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03166_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _01001_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02784_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _23530_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02984_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _03157_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03302_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03443_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03584_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03782_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03985_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04190_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04293_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04397_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04499_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04604_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04707_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04810_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04914_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _23899_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _24320_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _24321_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _24322_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _24323_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _24324_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _24325_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _24327_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _24306_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _24328_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _24329_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _24330_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _24331_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _24333_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _24334_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _24335_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _24307_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _24336_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _24337_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _24339_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _24340_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _24341_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _24342_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _24343_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _24308_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _23904_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _18908_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _23905_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _23906_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _18911_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _23907_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _23908_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18914_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _23909_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _18917_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _23910_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _23911_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _23912_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _18920_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _23913_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _18923_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _18926_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _18984_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _18986_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _18890_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _18989_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _18992_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _18893_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _18995_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _18896_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _18998_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _19001_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _19004_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _19007_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _19010_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _19013_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _19016_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _18899_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _18902_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _19019_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18905_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _25154_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _25261_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _25262_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _25263_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _25264_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _25265_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _25267_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _25268_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _25156_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _25269_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _25270_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _25271_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _25272_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _25273_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _25274_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _25275_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _25157_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _25276_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _25278_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _25279_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _25280_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _25281_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _25282_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _25283_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _25158_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _25284_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _25285_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _25286_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _25287_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _25289_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _25290_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _25291_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _25159_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _25292_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _25293_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _25294_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _25295_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _25296_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _25297_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _25298_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _25160_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _25300_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _25301_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _25302_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _25303_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _25304_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _25305_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _25306_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _25161_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _25307_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _25308_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _25309_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _25311_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _25312_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _25313_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _25314_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _25162_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _25315_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _25316_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _25317_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _25318_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _25319_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _25320_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _25322_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _25163_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _24692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _24693_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _24695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _24696_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _24405_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _24470_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _24472_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _24473_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _24474_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _24475_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _24476_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _24477_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _24478_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _24479_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _24480_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _24481_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _24483_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _24484_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _24485_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _24486_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _24370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _24490_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _24491_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _24492_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _24493_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _24494_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _24495_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _24497_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _24498_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _24499_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _24500_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _24501_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _24502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _24503_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _24504_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _24505_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _24372_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _24697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _24698_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _24699_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _24700_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _24701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _24702_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _24703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _24704_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _24706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _24707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _24708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _24709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _24710_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _24711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _24712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _24713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _24714_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _24715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _24717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _24718_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _24719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _24720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _24721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _24722_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _24723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _24724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _24725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _24726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _24728_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _24729_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _24730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _24429_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _24404_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _24731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _24732_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _24733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _24735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _24736_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _24737_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _24738_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _24406_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _24739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _24740_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _24741_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _24743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _24744_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _24745_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _24746_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _24407_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _24747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _24748_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _24749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _24750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _24751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _24752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _24754_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _24409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _24410_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _24411_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _24755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _24756_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _24757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _24758_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _24759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _24760_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _24761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _24412_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _24762_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _24763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _24765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _24766_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _24767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _24768_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _24769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _24770_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _24771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _24772_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _24773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _24774_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _24776_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _24777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _24778_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _24414_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _24779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _24780_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _24781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _24782_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _24783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _24784_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _24785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _24787_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _24788_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _24789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _24790_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _24791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _24792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _24793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _24794_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _24415_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _24416_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _24418_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _24417_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _24795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _24796_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _24798_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _24799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _24800_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _24801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _24802_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _24419_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _24803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _24804_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _24420_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _24805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _24806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _24807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _24809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _24810_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _24811_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _24812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _24421_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _24813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _24814_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _24815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _24816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _24817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _24818_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _24820_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _24422_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _24423_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _24821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _24822_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _24823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _24824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _24825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _24826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _24827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _24424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _24426_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _24427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _24828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _24829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _24831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _24428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _24832_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _24833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _24834_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _24835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _24836_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _24837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _24838_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _24839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _24840_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _24842_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _24843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _24844_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _24845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _24846_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _24847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _24848_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _24849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _24850_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _24851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _24853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _24854_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _24855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _24856_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _24857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _24858_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _24859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _24860_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _24861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _24862_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _24864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _24865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _24430_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _24866_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _24867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _24868_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _24869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _24870_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _24871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _24872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _24431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _24433_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _24434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _24873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _24875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _24876_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _24877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _24878_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _24879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _24880_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _24881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _24882_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _24883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _24884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _24886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _24887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _24888_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _24889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _24435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _24436_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _24437_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _24438_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _24890_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _24891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _24892_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _24893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _24894_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _24895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _24897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _24898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _24899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _24900_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _24901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _24902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _24903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _24904_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _24905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _24439_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _24440_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _25567_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _25586_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _25587_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _25588_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _25589_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _25590_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _25591_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _25592_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _25568_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25569_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _25593_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _25594_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _25571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _04005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _04008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _04011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _04014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _04017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _04021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _04024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _04026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _03999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _04030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _04033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _04036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _04039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _04042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _04045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _04049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _04051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _04055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _04058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _04061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _04064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _04067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _04070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _04073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _04076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _04278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _04281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _04284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _04287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _04290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _04294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _04297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _04300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _04253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _04256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _04259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _04262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _04266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _04269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _04272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _04274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _04228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _04231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _04234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _04238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _04241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _04244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _04247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _04249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _04855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _04858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _04861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _04864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _04867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _04870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _04873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _04876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _04830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _04834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _04837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _04840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _04843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _04846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _04849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _04851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _04805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _04808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _04812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _04815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _04818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _04821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _04824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _04826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _04779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _04782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _04785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _04788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _04791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _04794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _04797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _04799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _04754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _04757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _04760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _04763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _04766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _04769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _04772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _04775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _04730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _04733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _04736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _04739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _04742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _04745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _04748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _04750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _04704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _04708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _04711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _04714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _04717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _04720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _04723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _04726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _04679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _04682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _04685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _04688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _04691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _04694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _04698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _04700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _04655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _04658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _04661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _04664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _04667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _04670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _04673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _04676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _04630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _04633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _04636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _04639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _04642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _04646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _04649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _04651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _04605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _04608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _04611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _04614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _04618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _04621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _04624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _04626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _06067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _06070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _06073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _06076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _06079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _06082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _06085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _06088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _06043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _06046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _06049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _06052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _06055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _06058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _06061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _06064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _06018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _06021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _06024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _06027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _06030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _06033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _06037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _06039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _05993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _05996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _05999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _06002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _06005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _06009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _06012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _06014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _05968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _05971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _05974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _05977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _05980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _05984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _05987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _05989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _05943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _05946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _05949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _05952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _05956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _05959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _05962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _05964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _05919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _05922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _05925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _05928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _05931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _05934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _05937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _05940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _05894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _05897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _05900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _05904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _05907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _05910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _05913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _05915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _06314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _06317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _06320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _06323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _06326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _06329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _06333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _06335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _06289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _06292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _06295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _06298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _06301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _06305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _06308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _06310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _06264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _06267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _06270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _06273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _06277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _06280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _06283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _06286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _06239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _06242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _06245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _06249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _06252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _06255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _06258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _06260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _06339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _06342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _06345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _06348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _06351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _06354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _06357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _06360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _06487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _06490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _06493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _06496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _06499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _06502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _06505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _06508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _06462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _06466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _06469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _06472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _06475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _06478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _06481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _06483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _06438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _06441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _06447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _06450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _06453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _06456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _06458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0], _10034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1], _10038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2], _10042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3], _10046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4], _10050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5], _10054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6], _10058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7], _02706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _09997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _10001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _10005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _10009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _10013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _10017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _10021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _10024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _09965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _09969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _09973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _09977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _09981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _09985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _09989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _09992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _09933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _09937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _09941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _09945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _09949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _09953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _09957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _09960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _09901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _09905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _09909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _09913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _09917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _09921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _09925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _09928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _09869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _09873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _09877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _09881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _09885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _09889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _09893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _09896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _05475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _05478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _05481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _05484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _05487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _05490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _05493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _05495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _09837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _09841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _09845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _09849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _09853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _09857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _09861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _09864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _09805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _09809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _09813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _09817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _09821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _09825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _09829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _09832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _09773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _09777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _09781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _09785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _09789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _09793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _09797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _09800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _09741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _09745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _09749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _09753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _09757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _09761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _09765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _09768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _09709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _09713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _09717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _09721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _09725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _09729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _09733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _09736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _09684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _09687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _09690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _09693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _09696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _09699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _09702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _09704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _09659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _09662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _09665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _09668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _09671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _09674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _09677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _09680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _09635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _09638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _09641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _09644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _09647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _09650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _09653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _09656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _09610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _09613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _09616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _09619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _09622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _09625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _09629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _09631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _09585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _09588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _09591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _09594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _09597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _09601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _09604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _09606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _09561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _09564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _09567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _09570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _09573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _09576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _09579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _09582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _09535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _09538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _09541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _09544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _09548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _09551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _09554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _09556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _09511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _09514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _09517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _09520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _09523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _09526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _09529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _09532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _09485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _09488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _09491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _09495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _09499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _09502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _09505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _09507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _05426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _05429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _05432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _05435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _05438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _05441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _05444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _05446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _09459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _09462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _09466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _09469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _09472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _09476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _09479_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _09481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _05450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _05453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _05456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _05459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _05462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _05465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _05468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _05471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _09435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _09438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _09441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _09444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _09447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _09450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _09453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _09456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _09410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _09414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _09417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _09420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _09423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _09426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _09429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _09431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _09386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _09389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _09392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _09395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _09398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _09401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _09404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _09406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _09361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _09364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _09367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _09370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _09373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _09376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _09379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _09382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _09337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _09340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _09343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _09346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _09349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _09352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _09355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _09357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _09312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _09315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _09318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _09321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _09324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _09327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _09330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _09333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _05401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _05404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _05407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _05410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _05413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _05416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _05419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _05422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _05376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _05379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _05382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _05385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _05388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _05391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _05395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _05397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _05327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _05330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _05333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _05336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _05339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _05342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _05345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _05348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _05302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _05305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _05308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _05311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _05315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _05318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _05321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _05323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _05277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _05280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _05283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _05287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _05290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _05293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _05296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _05298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _03613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _03616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _03619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _03622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _03626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _03629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _03632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _03634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _05228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _05231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _05235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _05238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _05241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _05244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _05247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _05249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _03577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _03581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _03587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _03591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _03595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _03600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _03605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _03607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _03694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _03697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _03700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _03704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _03707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _03710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _03713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _03716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _03667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _03670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _03673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _03676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _03679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _03682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _03685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _03688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _03641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _03644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _03647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _03650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _03653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _03656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _03659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _03662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _03745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _03748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _03720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _03723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _03726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _03729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _03733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _03736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _03739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _03741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _05253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _05256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _05259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _05262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _05265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _05268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _05271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _05274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _09287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _09290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _09293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _09296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _09299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _09302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _09306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _09308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _09262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _09265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _09268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _09271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _09274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _09278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _09281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _09284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _09238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _09241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _09244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _09247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _09250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _09253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _09256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _09259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _09213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _09216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _09219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _09222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _09226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _09229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _09232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _09234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _09188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _09191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _09194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _09198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _09201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _09204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _09207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _09209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _09164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _09167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _09170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _09173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _09176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _09179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _09182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _09185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _09138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _09141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _09145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _09148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _09151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _09154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _09157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _09159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _09114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _09117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _09120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _09123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _09126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _09129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _09132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _09135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _09089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _09093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _09096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _09099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _09102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _09105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _09108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _09110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _09065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _09068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _09071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _09074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _09077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _09080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _09083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _09085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _09040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _09043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _09046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _09049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _09052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _09055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _09058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _09061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _09016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _09019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _09022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _09025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _09028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _09031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _09034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _09036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _08991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _08994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _08997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _09000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _09003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _09006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _09009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _09012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _08966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _08969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _08972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _08975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _08978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _08981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _08985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _08987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _08942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _08945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _08948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _08951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _08954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _08957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _08960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _08963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _08917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _08920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _08923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _08926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _08929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _08933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _08936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _08938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _08890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _08893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _08896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _08900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _08904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _08907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _08911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _08913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _08863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _08867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _08870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _08873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _08877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _08880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _08883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _08886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _08836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _08839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _08843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _08847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _08850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _08854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _08857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _08859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _08811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _08814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _08818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _08821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _08824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _08827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _08830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _08832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _08786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _08790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _08793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _08796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _08799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _08802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _08805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _08807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _08762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _08765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _08768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _08771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _08774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _08777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _08780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _08783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _08737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _08740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _08743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _08746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _08749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _08752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _08755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _08757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _08712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _08715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _08718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _08721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _08724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _08727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _08730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _08733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _08688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _08691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _08694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _08697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _08700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _08703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _08706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _08708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _08663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _08666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _08669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _08672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _08675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _08678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _08681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _08684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _08638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _08641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _08644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _08647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _08650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _08653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _08657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _08659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _08614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _08617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _08620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _08623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _08626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _08629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _08632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _08635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _08589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _08592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _08595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _08598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _08601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _08605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _08608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _08610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _08564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _08567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _08570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _08573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _08577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _08580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _08583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _08585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _08540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _08543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _08546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _08549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _08552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _08555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _08558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _08561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _08515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _08518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _08521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _08525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _08528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _08531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _08534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _08536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _08490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _08493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _08497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _08500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _08503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _08506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _08509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _08511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _08466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _08469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _08472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _08475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _08478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _08481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _08484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _08487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _08441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _08445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _08448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _08451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _08454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _08457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _08460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _08462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _08417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _08420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _08423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _08426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _08429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _08432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _08435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _08437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _08392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _08395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _08398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _08401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _08404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _08407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _08410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _08412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _08367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _08370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _08373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _08376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _08379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _08382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _08385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _08388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _08341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _08344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _08347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _08350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _08353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _08356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _08359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _08362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _08317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _08320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _08323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _08326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _08329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _08332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _08335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _08338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _08292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _08295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _08298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _08301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _08304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _08307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _08311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _08313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _08267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _08270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _08273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _08276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _08279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _08283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _08286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _08288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _06413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _06416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _06419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _06422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _06425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _06428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _06431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _06434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _06215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _06218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _06221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _06224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _06227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _06230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _06233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _06236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _05869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _05872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _05876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _05879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _05882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _05885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _05888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _05890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _05844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _05848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _05851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _05854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _05857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _05860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _05863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _05866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _05820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _05823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _05826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _05829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _05832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _05835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _05838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _05841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _05796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _05799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _05802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _05805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _05808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _05811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _05814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _05816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _05771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _05774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _05777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _05780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _05783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _05786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _05789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _05791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _05746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _05749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _05752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _05755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _05758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _05761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _05764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _05767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _05722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _05725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _05728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _05731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _05734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _05737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _05740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _05743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _05697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _05700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _05703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _05706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _05709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _05712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _05716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _05718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _05672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _05675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _05678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _05681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _05684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _05688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _05691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _05693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _05648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _05651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _05654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _05657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _05660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _05663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _05666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _05669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _05623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _05626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _05629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _05632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _05636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _05639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _05642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _05644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _05598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _05601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _05604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _05608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _05611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _05614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _05617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _05619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _05573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _05576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _05579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _05583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _05586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _05589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _05592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _05594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _05548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _05551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _05555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _05558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _05561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _05564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _05567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _05569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _05524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _05527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _05530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _05533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _05536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _05539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _05542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _05545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _05499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _05503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _05506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _05509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _05512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _05515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _05518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _05520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _04580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _04583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _04586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _04589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _04592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _04595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _04598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _04601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _04930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _04933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _04936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _04939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _04942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _04945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _04948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _04951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _04554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _04557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _04561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _04565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _04568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _04571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _04574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _04576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _04904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _04907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _04910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _04915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _04918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _04921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _04924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _04926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _04529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _04533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _04536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _04539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _04542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _04545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _04548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _04550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _04879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _04882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _04886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _04889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _04892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _04895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _04898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _04900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _04505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _04508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _04511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _04514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _04517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _04520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _04523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _04526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _04480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _04483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _04486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _04489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _04492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _04495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _04498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _04501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _04455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _04458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _04461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _04464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _04467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _04470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _04473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _04475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _04430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _04433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _04436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _04439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _04442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _04445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _04448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _04451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _04406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _04409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _04412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _04415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _04418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _04421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _04424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _04427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _04377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _04380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _04383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _04386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _04389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _04392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _04395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _04399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _04353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _04356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _04359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _04362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _04365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _04368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _04371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _04374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _04328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _04331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _04334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _04337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _04340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _04343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _04347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _04349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _04303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _04306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _04309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _04312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _04315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _04319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _04322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _04324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _04204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _04207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _04210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _04213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _04216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _04219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _04222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _04225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _06117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _06120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _06123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _06126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _06129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _06132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _06135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _06137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _07946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _07949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _07952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _07955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _07958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _07962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _07965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _07967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _07675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _07678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _07681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _07684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _07687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _07690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _07694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _07696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _07651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _07654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _07657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _07660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _07663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _07666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _07669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _07672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _06935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _06938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _06941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _06944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _06947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _06950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _06953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _06956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _06984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _06987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _06990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _06993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _06996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _07000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _07003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _07005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _06959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _06962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _06965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _06968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _06972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _06975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _06978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _06980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _06685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _06688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _06691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _06694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _06697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _06700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _06703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _06706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _06660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _06663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _06666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _06669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _06672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _06675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _06679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _06681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _06092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _06095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _06098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _06101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _06104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _06107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _06110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _06112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _06141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _06144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _06147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _06150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _06153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _06156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _06159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _06162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _05351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _05354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _05357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _05360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _05363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _05367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _05370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _05372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _05203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _05207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _05210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _05213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _05216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _05219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _05222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _05224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _05053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _05056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _05059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _05062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _05065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _05068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _05071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _05074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _05176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _05179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _05183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _05186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _05189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _05192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _05195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _05197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _05151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _05155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _05158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _05161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _05164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _05167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _05170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _05172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _05127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _05130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _05133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _05136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _05139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _05142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _05145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _05148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _05103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _05106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _05109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _05112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _05115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _05118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _05121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _05123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _05078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _05081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _05084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _05087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _05090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _05093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _05096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _05098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _05029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _05032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _05035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _05038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _05041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _05044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _05047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _05050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _05004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _05007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _05010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _05013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _05016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _05019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _05023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _05025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _04979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _04982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _04985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _04988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _04991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _04995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _04998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _05000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _04954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _04957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _04960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _04963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _04967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _04970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _04973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _04975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _04178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _04181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _04185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _04188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _04192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _04195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _04198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _04200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _04153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _04157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _04160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _04163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _04166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _04169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _04172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _04174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _04129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _04132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _04135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _04138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _04141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _04144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _04147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _04150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _04104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _04107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _04110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _04113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _04116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _04119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _04122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _04124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _04079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _04082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _04085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _04088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _04091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _04094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _04097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _04100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _08243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _08246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _08249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _08252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _08255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _08258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _08261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _08264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _08218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _08221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _08224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _08227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _08231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _08234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _08237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _08239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _08193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _08196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _08199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _08203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _08206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _08209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _08212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _08214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _08169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _08172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _08175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _08178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _08181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _08184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _08187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _08190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _08144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _08147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _08151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _08154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _08157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _08160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _08163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _08165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _08119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _08123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _08126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _08129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _08132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _08135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _08138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _08140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _08095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _08098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _08101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _08104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _08107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _08110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _08113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _08116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _08071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _08074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _08077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _08080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _08083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _08086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _08089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _08091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _07921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _07924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _07927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _07930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _07934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _07937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _07940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _07942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _08046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _08049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _08052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _08055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _08058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _08061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _08064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _08066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _08021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _08024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _08027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _08030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _08033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _08036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _08039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _08042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _07971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _07974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _07977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _07980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _07983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _07987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _07991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _07993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _07997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _08000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _08003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _08006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _08009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _08012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _08015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _08018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _07897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _07900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _07903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _07906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _07909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _07912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _07915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _07918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _07872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _07875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _07878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _07882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _07885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _07888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _07891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _07893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _07823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _07826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _07829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _07832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _07835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _07838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _07841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _07844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _07847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _07850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _07854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _07857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _07860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _07863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _07866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _07868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _07798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _07802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _07805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _07808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _07811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _07814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _07817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _07819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _07774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _07777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _07780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _07783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _07786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _07789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _07792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _07794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _07749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _07752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _07755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _07758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _07761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _07764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _07767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _07770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _07725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _07728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _07731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _07734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _07737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _07740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _07743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _07745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _07700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _07703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _07706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _07709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _07712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _07715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _07718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _07721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _07626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _07629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _07632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _07635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _07638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _07642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _07645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _07647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _07601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _07604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _07607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _07610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _07614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _07617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _07620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _07622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _07551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _07554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _07557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _07561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _07564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _07567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _07570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _07572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _07577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _07580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _07583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _07586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _07589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _07592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _07595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _07598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _07502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _07505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _07508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _07511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _07514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _07517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _07520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _07523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _07526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _07529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _07533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _07536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _07539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _07542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _07545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _07547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _07477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _07481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _07484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _07487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _07490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _07493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _07496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _07498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _07453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _07456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _07459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _07462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _07465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _07468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _07471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _07473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _07428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _07431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _07434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _07437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _07440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _07443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _07446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _07449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _07379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _07382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _07385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _07388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _07391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _07394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _07397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _07400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _07404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _07407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _07410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _07413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _07416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _07419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _07422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _07424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _07354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _07357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _07360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _07363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _07366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _07369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _07373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _07375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _07330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _07333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _07336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _07339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _07342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _07345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _07348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _07351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _07305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _07308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _07311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _07314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _07317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _07321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _07324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _07326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _07256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _07259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _07262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _07265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _07268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _07271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _07274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _07277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _07280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _07283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _07286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _07289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _07293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _07296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _07299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _07301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _07231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _07234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _07237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _07241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _07244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _07247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _07250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _07252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _07206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _07209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _07213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _07216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _07219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _07222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _07225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _07227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _07182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _07185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _07188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _07191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _07194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _07197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _07200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _07203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _07132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _07135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _07138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _07141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _07144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _07147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _07150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _07153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _07156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _07160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _07163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _07166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _07169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _07172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _07175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _07177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _07107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _07110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _07113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _07116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _07119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _07122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _07125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _07128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _07083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _07086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _07089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _07092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _07095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _07098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _07101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _07103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _07058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _07061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _07064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _07067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _07070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _07073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _07079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _07033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _07036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _07039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _07042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _07045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _07048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _07052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _07054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _07009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _07012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _07015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _07018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _07021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _07024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _07027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _07030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _06885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _06888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _06892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _06895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _06898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _06901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _06904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _06906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _06910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _06913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _06916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _06920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _06923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _06926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _06931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _06861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _06864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _06867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _06870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _06873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _06876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _06879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _06882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _06836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _06840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _06843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _06846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _06849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _06852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _06855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _06857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _06812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _06815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _06818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _06821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _06824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _06827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _06830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _06832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _06759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _06762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _06765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _06768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _06771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _06774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _06777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _06780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _06787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _06790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _06793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _06796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _06799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _06802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _06805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _06808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _06735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _06738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _06741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _06744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _06747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _06750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _06753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _06755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _06710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _06713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _06716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _06719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _06722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _06725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _06728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _06730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _06511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _06514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _06518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _06521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _06525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _06528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _06531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _06533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _06636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _06639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _06642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _06645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _06648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _06651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _06654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _06657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _06611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _06614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _06617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _06620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _06623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _06627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _06630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _06632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _06586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _06589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _06592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _06595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _06599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _06602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _06605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _06607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _06537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _06540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _06543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _06547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _06550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _06553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _06556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _06558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _06562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _06565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _06568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _06571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _06574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _06577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _06580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _06583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _06363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _06366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _06369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _06372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _06375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _06378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _06381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _06384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _06389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _06392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _06395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _06398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _06401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _06404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _06407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _06409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _06190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _06193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _06197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _06200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _06203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _06206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _06209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _06211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _06165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _06169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _06172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _06175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _06178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _06181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _06184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _06186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _15236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _15238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _15240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _15242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _15244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _15246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _15248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02715_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _25387_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _25485_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _25486_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _25487_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _25388_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _25389_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _25391_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _25488_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _25489_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _25490_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _25492_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _25493_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _25494_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _25495_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _25392_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _25393_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19498_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19508_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19518_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19528_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17824_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08864_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08876_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08887_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08898_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06524_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13716_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13738_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12743_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13760_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13771_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13782_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _27359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _27357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _27355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _27353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _27351_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _27349_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _27347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _27345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _27343_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _27341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _27307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _27305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _27303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _27301_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _27298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00176_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00182_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00188_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _27296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00190_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00192_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00194_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00196_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00198_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00200_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00202_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _27294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _24987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _24989_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _24991_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _24993_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _24995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _24997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _24999_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _23900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _25001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _25003_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _25005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _25007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _25009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _25011_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _25013_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _23901_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _25015_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _25017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _25019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _25021_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _25023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _25025_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _25027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _23902_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _25029_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _25031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _25033_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _25035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _25037_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _25039_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _25041_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _23903_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17315_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15222_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09474_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10773_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10784_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09496_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _25436_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _25439_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _26040_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _26042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _26044_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _26046_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _26048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _26050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _26052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _25442_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _26054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _26056_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _26058_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _26060_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _26062_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _26064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _26066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _25445_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _25448_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _25451_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _26068_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _26070_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _26072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _26074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _26076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _26078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _26080_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _25454_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _26082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _26084_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _26086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _26088_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _26090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _26092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _26094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _25457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _25460_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _26096_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _26098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _26100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _26102_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _26104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _26106_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _26108_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _25463_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02205_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02207_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02223_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02227_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02229_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01661_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02251_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02253_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01667_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02259_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02265_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02267_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01241_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00598_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01260_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00604_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01262_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01267_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01269_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01277_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00617_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01286_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01299_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01301_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00632_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00637_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
