
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jnc, ABINPUT, ABINPUT000, ABINPUT000000);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  input [8:0] ABINPUT;
  input [16:0] ABINPUT000;
  input [16:0] ABINPUT000000;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [16:0] \oc8051_top_1.ABINPUT000 ;
  wire [16:0] \oc8051_top_1.ABINPUT000000 ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT000 ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire \oc8051_top_1.oc8051_alu1.divOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.mulOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jnc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_05110_, rst);
  not (_05111_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_05112_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  not (_05113_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05114_, _05113_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_05115_, _05114_, _05112_);
  or (_05116_, _05115_, _05111_);
  not (_05117_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_05118_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_05119_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _05113_);
  nand (_05120_, _05119_, _05118_);
  or (_05121_, _05120_, _05117_);
  and (_05122_, _05121_, _05116_);
  not (_05123_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_05124_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_05125_, _05124_, _05113_);
  nor (_05126_, _05125_, _05123_);
  and (_05127_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_05128_, _05127_, _05112_);
  not (_05129_, _05128_);
  and (_05130_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_05131_, _05130_, _05126_);
  and (_05132_, _05131_, _05122_);
  nor (_05133_, _05124_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_05134_, _05133_);
  not (_05135_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_05136_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05135_);
  or (_05137_, _05136_, ABINPUT[5]);
  nand (_05138_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05135_);
  or (_05139_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_05140_, _05139_, _05137_);
  or (_05141_, _05140_, _05134_);
  not (_05142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_05143_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_05144_, _05143_, _05113_);
  nor (_05145_, _05144_, _05142_);
  and (_05146_, _05127_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_05147_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_05148_, _05147_, _05145_);
  and (_05149_, _05148_, _05141_);
  and (_05150_, _05149_, _05132_);
  not (_05151_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_05152_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05151_);
  and (_05153_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05151_);
  nor (_05154_, _05153_, _05152_);
  and (_05155_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _05151_);
  and (_05156_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _05151_);
  nor (_05157_, _05156_, _05155_);
  and (_05158_, _05157_, _05154_);
  not (_05159_, _05158_);
  not (_05160_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not (_05162_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_05163_, _05152_, _05162_);
  nand (_05164_, _05163_, _05160_);
  nand (_05165_, _05154_, _05156_);
  and (_05166_, _05165_, _05164_);
  and (_05167_, _05166_, _05159_);
  and (_05168_, _05153_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  nand (_05169_, _05168_, _05160_);
  not (_05170_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_05171_, _05153_, _05170_);
  and (_05172_, _05171_, _05155_);
  not (_05174_, _05172_);
  and (_05175_, _05174_, _05169_);
  and (_05176_, _05175_, _05167_);
  nor (_05177_, _05176_, _05150_);
  not (_05178_, _05177_);
  and (_05180_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_05181_, _05180_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_05182_, _05181_);
  or (_05183_, _05136_, ABINPUT[0]);
  or (_05184_, _05138_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_05185_, _05184_, _05183_);
  or (_05186_, _05185_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_05187_, _05186_, _05182_);
  not (_05188_, _05187_);
  not (_05189_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_05190_, _05115_, _05189_);
  not (_05191_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or (_05192_, _05120_, _05191_);
  and (_05193_, _05192_, _05190_);
  nand (_05194_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_05195_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_05196_, _05125_, _05195_);
  and (_05197_, _05196_, _05194_);
  and (_05198_, _05197_, _05193_);
  or (_05199_, _05136_, ABINPUT[4]);
  or (_05200_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_05201_, _05200_, _05199_);
  or (_05202_, _05201_, _05134_);
  nand (_05203_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not (_05204_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_05206_, _05144_, _05204_);
  and (_05207_, _05206_, _05203_);
  and (_05209_, _05207_, _05202_);
  and (_05210_, _05209_, _05198_);
  not (_05211_, _05210_);
  not (_05212_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_05213_, _05115_, _05212_);
  not (_05214_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or (_05215_, _05120_, _05214_);
  and (_05217_, _05215_, _05213_);
  not (_05218_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_05219_, _05125_, _05218_);
  not (_05220_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_05221_, _05128_, _05220_);
  and (_05222_, _05221_, _05219_);
  and (_05223_, _05222_, _05217_);
  or (_05224_, _05136_, ABINPUT[3]);
  or (_05225_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_05226_, _05225_, _05224_);
  or (_05227_, _05226_, _05134_);
  not (_05228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_05229_, _05144_, _05228_);
  nand (_05230_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and (_05231_, _05230_, _05229_);
  and (_05232_, _05231_, _05227_);
  and (_05233_, _05232_, _05223_);
  not (_05234_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or (_05235_, _05115_, _05234_);
  not (_05236_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  or (_05237_, _05120_, _05236_);
  and (_05238_, _05237_, _05235_);
  nand (_05239_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_05240_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_05241_, _05125_, _05240_);
  and (_05242_, _05241_, _05239_);
  and (_05243_, _05242_, _05238_);
  or (_05244_, _05136_, ABINPUT[1]);
  or (_05245_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_05246_, _05245_, _05244_);
  or (_05247_, _05246_, _05134_);
  nand (_05248_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not (_05249_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_05250_, _05144_, _05249_);
  and (_05251_, _05250_, _05248_);
  and (_05252_, _05251_, _05247_);
  and (_05253_, _05252_, _05243_);
  or (_05254_, _05136_, ABINPUT[2]);
  or (_05255_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_05256_, _05255_, _05254_);
  or (_05257_, _05256_, _05134_);
  not (_05258_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_05259_, _05115_, _05258_);
  not (_05260_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or (_05261_, _05120_, _05260_);
  and (_05262_, _05261_, _05259_);
  and (_05263_, _05262_, _05257_);
  not (_05264_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_05265_, _05125_, _05264_);
  not (_05266_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_05267_, _05128_, _05266_);
  and (_05268_, _05267_, _05265_);
  not (_05269_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_05270_, _05144_, _05269_);
  nand (_05271_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_05272_, _05271_, _05270_);
  and (_05273_, _05272_, _05268_);
  and (_05274_, _05273_, _05263_);
  and (_05275_, _05274_, _05253_);
  nand (_05276_, _05275_, _05233_);
  or (_05277_, _05276_, _05211_);
  or (_05278_, _05277_, _05188_);
  not (_05279_, _05233_);
  nand (_05280_, _05252_, _05243_);
  nand (_05281_, _05273_, _05263_);
  and (_05282_, _05281_, _05280_);
  nand (_05283_, _05282_, _05279_);
  or (_05284_, _05283_, _05210_);
  or (_05285_, _05284_, _05187_);
  and (_05286_, _05285_, _05278_);
  or (_05287_, _05286_, _05150_);
  not (_05288_, _05155_);
  nor (_05290_, _05288_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_05291_, _05168_, _05290_);
  nand (_05292_, _05286_, _05150_);
  and (_05293_, _05292_, _05291_);
  nand (_05294_, _05293_, _05287_);
  and (_05295_, _05171_, _05157_);
  nor (_05296_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not (_05297_, _05296_);
  nor (_05298_, _05297_, _05140_);
  not (_05299_, _05298_);
  and (_05300_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05301_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_05302_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_05303_, _05302_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05304_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_05305_, _05304_, _05301_);
  and (_05306_, _05305_, _05299_);
  nor (_05307_, _05306_, _05150_);
  and (_05308_, _05306_, _05150_);
  nor (_05309_, _05308_, _05307_);
  nand (_05310_, _05309_, _05295_);
  and (_05311_, _05155_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_05312_, _05311_, _05163_);
  and (_05313_, _05312_, _05307_);
  and (_05314_, _05290_, _05163_);
  and (_05316_, _05314_, _05150_);
  nor (_05317_, _05316_, _05313_);
  and (_05318_, _05188_, _05150_);
  not (_05319_, _05318_);
  and (_05320_, _05168_, _05311_);
  not (_05321_, _05320_);
  and (_05322_, _05306_, _05187_);
  nor (_05323_, _05322_, _05321_);
  and (_05324_, _05323_, _05319_);
  and (_05325_, _05156_, _05160_);
  and (_05326_, _05171_, _05325_);
  not (_05327_, _05326_);
  nor (_05328_, _05327_, _05308_);
  nor (_05329_, _05328_, _05324_);
  and (_05330_, _05329_, _05317_);
  and (_05332_, _05330_, _05310_);
  and (_05333_, _05332_, _05294_);
  and (_05334_, _05333_, _05178_);
  not (_05335_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_05336_, \oc8051_top_1.oc8051_decoder1.wr , _05151_);
  and (_05337_, _05336_, _05335_);
  not (_05338_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05339_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05151_);
  and (_05340_, _05339_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_05341_, _05340_, _05338_);
  and (_05343_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_05344_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_05345_, _05344_, _05343_);
  and (_05346_, _05345_, _05341_);
  and (_05347_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05151_);
  nor (_05348_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05349_, _05348_, _05347_);
  and (_05350_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_05351_, _05350_, _05346_);
  not (_05352_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_05353_, _05339_, _05352_);
  nand (_05354_, _05353_, _05338_);
  or (_05355_, _05354_, _05258_);
  and (_05356_, _05353_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nand (_05357_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nor (_05358_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor (_05359_, _05358_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_05361_, _05359_, _05339_);
  nand (_05362_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_05363_, _05362_, _05357_);
  and (_05364_, _05363_, _05355_);
  and (_05365_, _05364_, _05351_);
  and (_05366_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_05367_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_05368_, _05367_, _05366_);
  not (_05369_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_05370_, _05341_, _05369_);
  or (_05371_, _05354_, _05234_);
  nand (_05372_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nand (_05373_, _05372_, _05371_);
  nor (_05374_, _05373_, _05370_);
  and (_05375_, _05374_, _05368_);
  and (_05376_, _05375_, _05365_);
  nand (_05377_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or (_05378_, _05354_, _05189_);
  and (_05379_, _05378_, _05377_);
  and (_05380_, _05343_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nand (_05381_, _05380_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  or (_05382_, _05380_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_05383_, _05382_, _05381_);
  nand (_05384_, _05383_, _05341_);
  nand (_05385_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nand (_05386_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and (_05387_, _05386_, _05385_);
  and (_05388_, _05387_, _05384_);
  and (_05389_, _05388_, _05379_);
  not (_05390_, _05389_);
  nor (_05391_, _05343_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_05392_, _05391_, _05380_);
  and (_05393_, _05392_, _05341_);
  and (_05394_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_05395_, _05394_, _05393_);
  or (_05396_, _05354_, _05212_);
  nand (_05397_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  nand (_05398_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  and (_05399_, _05398_, _05397_);
  and (_05400_, _05399_, _05396_);
  and (_05401_, _05400_, _05395_);
  and (_05402_, _05401_, _05390_);
  and (_05403_, _05402_, _05376_);
  and (_05404_, _05380_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_05405_, _05404_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_05406_, _05404_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nand (_05407_, _05406_, _05341_);
  or (_05408_, _05407_, _05405_);
  nand (_05409_, _05356_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nand (_05410_, _05340_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nand (_05411_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  and (_05412_, _05411_, _05410_);
  and (_05413_, _05412_, _05409_);
  or (_05414_, _05354_, _05111_);
  nand (_05415_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_05416_, _05415_, _05414_);
  and (_05417_, _05416_, _05413_);
  and (_05418_, _05417_, _05408_);
  not (_05419_, _05418_);
  nand (_05420_, _05405_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  or (_05421_, _05405_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_05422_, _05421_, _05341_);
  nand (_05423_, _05422_, _05420_);
  nand (_05424_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  not (_05425_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_05426_, _05354_, _05425_);
  nand (_05427_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_05429_, _05427_, _05410_);
  and (_05431_, _05429_, _05426_);
  and (_05432_, _05431_, _05424_);
  and (_05433_, _05432_, _05423_);
  and (_05434_, _05433_, _05419_);
  and (_05435_, _05405_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand (_05436_, _05435_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or (_05437_, _05435_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_05438_, _05437_, _05341_);
  nand (_05439_, _05438_, _05436_);
  nand (_05440_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_05441_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  or (_05442_, _05354_, _05441_);
  nand (_05443_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_05444_, _05443_, _05410_);
  and (_05445_, _05444_, _05442_);
  and (_05446_, _05445_, _05440_);
  and (_05447_, _05446_, _05439_);
  not (_05448_, _05447_);
  nand (_05449_, _05436_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or (_05450_, _05436_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_05451_, _05450_, _05449_);
  nand (_05452_, _05451_, _05341_);
  nand (_05453_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  not (_05454_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or (_05455_, _05354_, _05454_);
  nand (_05456_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_05457_, _05456_, _05410_);
  and (_05458_, _05457_, _05455_);
  and (_05459_, _05458_, _05453_);
  nand (_05460_, _05459_, _05452_);
  nor (_05461_, _05460_, _05448_);
  and (_05462_, _05461_, _05434_);
  and (_05463_, _05462_, _05403_);
  and (_05464_, _05463_, _05337_);
  not (_05465_, _05464_);
  nor (_05466_, _05465_, _05334_);
  not (_05467_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_05468_, _05464_, _05467_);
  or (_05469_, _05468_, _05466_);
  and (_05161_, _05469_, _05110_);
  not (_05470_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor (_05471_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_05472_, _05471_, _05470_);
  nor (_05473_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_05474_, _05473_, _05151_);
  and (_05475_, _05474_, _05472_);
  and (pc_log_change, _05475_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_05476_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not (_05478_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_05479_, pc_log_change, _05478_);
  and (_05480_, _05479_, _05110_);
  and (_06782_, _05480_, _05476_);
  and (_05481_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_05482_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_05483_, pc_log_change, _05482_);
  or (_05484_, _05483_, _05481_);
  and (_06919_, _05484_, _05110_);
  not (_05485_, _05401_);
  not (_05486_, _05365_);
  and (_05487_, _05375_, _05486_);
  and (_05488_, _05487_, _05485_);
  and (_05489_, _05325_, _05154_);
  not (_05490_, _05489_);
  nor (_05491_, _05115_, _05454_);
  not (_05492_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_05493_, _05120_, _05492_);
  nor (_05494_, _05493_, _05491_);
  and (_05495_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_05496_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_05497_, _05125_, _05496_);
  nor (_05498_, _05497_, _05495_);
  and (_05499_, _05498_, _05494_);
  nor (_05500_, _05136_, ABINPUT[8]);
  nor (_05501_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor (_05502_, _05501_, _05500_);
  and (_05503_, _05502_, _05133_);
  not (_05504_, _05503_);
  and (_05505_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  not (_05506_, _05144_);
  and (_05507_, _05506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_05508_, _05507_, _05505_);
  and (_05509_, _05508_, _05504_);
  and (_05510_, _05509_, _05499_);
  and (_05511_, _05502_, _05296_);
  not (_05512_, _05511_);
  and (_05514_, _05300_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_05515_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_05516_, _05515_, _05514_);
  and (_05517_, _05516_, _05512_);
  nor (_05518_, _05517_, _05510_);
  not (_05519_, _05518_);
  and (_05520_, _05517_, _05510_);
  or (_05521_, _05297_, _05201_);
  and (_05522_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_05523_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_05524_, _05523_, _05522_);
  and (_05526_, _05524_, _05521_);
  nor (_05527_, _05526_, _05210_);
  and (_05528_, _05526_, _05210_);
  nor (_05529_, _05528_, _05527_);
  or (_05530_, _05297_, _05226_);
  and (_05531_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_05532_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_05533_, _05532_, _05531_);
  and (_05534_, _05533_, _05530_);
  nor (_05535_, _05534_, _05233_);
  not (_05536_, _05535_);
  and (_05537_, _05534_, _05233_);
  nor (_05538_, _05537_, _05535_);
  or (_05539_, _05297_, _05256_);
  nand (_05540_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand (_05541_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_05542_, _05541_, _05540_);
  nand (_05543_, _05542_, _05539_);
  and (_05544_, _05543_, _05281_);
  or (_05545_, _05297_, _05246_);
  nand (_05546_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand (_05547_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_05548_, _05547_, _05546_);
  and (_05549_, _05548_, _05545_);
  not (_05550_, _05549_);
  and (_05551_, _05550_, _05280_);
  and (_05552_, _05542_, _05539_);
  and (_05553_, _05552_, _05274_);
  nor (_05554_, _05553_, _05544_);
  and (_05555_, _05554_, _05551_);
  or (_05556_, _05555_, _05544_);
  nand (_05557_, _05556_, _05538_);
  nand (_05558_, _05557_, _05536_);
  nand (_05559_, _05558_, _05529_);
  or (_05560_, _05558_, _05529_);
  and (_05561_, _05560_, _05559_);
  and (_05562_, _05549_, _05253_);
  nor (_05563_, _05562_, _05551_);
  and (_05564_, _05563_, _05187_);
  and (_05566_, _05564_, _05554_);
  or (_05567_, _05556_, _05538_);
  and (_05568_, _05567_, _05557_);
  and (_05570_, _05568_, _05566_);
  and (_05571_, _05570_, _05561_);
  not (_05572_, _05528_);
  and (_05573_, _05558_, _05572_);
  or (_05574_, _05573_, _05527_);
  or (_05575_, _05574_, _05571_);
  nand (_05576_, _05575_, _05309_);
  nor (_05577_, _05115_, _05425_);
  not (_05578_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor (_05579_, _05120_, _05578_);
  nor (_05580_, _05579_, _05577_);
  not (_05581_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_05582_, _05125_, _05581_);
  not (_05583_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_05584_, _05128_, _05583_);
  nor (_05585_, _05584_, _05582_);
  and (_05586_, _05585_, _05580_);
  nor (_05587_, _05136_, ABINPUT[6]);
  nor (_05588_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor (_05589_, _05588_, _05587_);
  and (_05590_, _05589_, _05133_);
  not (_05591_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05592_, _05144_, _05591_);
  and (_05593_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nor (_05594_, _05593_, _05592_);
  not (_05595_, _05594_);
  nor (_05596_, _05595_, _05590_);
  and (_05597_, _05596_, _05586_);
  and (_05598_, _05589_, _05296_);
  not (_05599_, _05598_);
  and (_05600_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_05601_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05602_, _05601_, _05600_);
  and (_05603_, _05602_, _05599_);
  and (_05604_, _05603_, _05597_);
  nor (_05605_, _05603_, _05597_);
  nor (_05606_, _05605_, _05604_);
  not (_05607_, _05606_);
  or (_05608_, _05607_, _05576_);
  nor (_05609_, _05115_, _05441_);
  not (_05610_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_05611_, _05120_, _05610_);
  nor (_05612_, _05611_, _05609_);
  not (_05613_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_05614_, _05125_, _05613_);
  and (_05615_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_05616_, _05615_, _05614_);
  and (_05617_, _05616_, _05612_);
  nor (_05618_, _05136_, ABINPUT[7]);
  nor (_05619_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor (_05620_, _05619_, _05618_);
  and (_05621_, _05620_, _05133_);
  not (_05622_, _05621_);
  and (_05623_, _05506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_05624_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_05625_, _05624_, _05623_);
  and (_05626_, _05625_, _05622_);
  and (_05627_, _05626_, _05617_);
  and (_05628_, _05620_, _05296_);
  not (_05629_, _05628_);
  and (_05630_, _05300_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and (_05631_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_05632_, _05631_, _05630_);
  and (_05633_, _05632_, _05629_);
  nor (_05634_, _05633_, _05627_);
  and (_05635_, _05633_, _05627_);
  nor (_05636_, _05635_, _05634_);
  not (_05637_, _05636_);
  and (_05638_, _05606_, _05307_);
  nor (_05639_, _05638_, _05605_);
  nor (_05640_, _05639_, _05637_);
  and (_05641_, _05639_, _05637_);
  nor (_05642_, _05641_, _05640_);
  not (_05643_, _05642_);
  or (_05644_, _05643_, _05608_);
  nor (_05645_, _05640_, _05634_);
  and (_05646_, _05645_, _05644_);
  or (_05647_, _05646_, _05520_);
  and (_05648_, _05647_, _05519_);
  or (_05649_, _05648_, _05490_);
  and (_05650_, _05290_, _05154_);
  not (_05651_, _05650_);
  not (_05652_, _05517_);
  and (_05653_, _05652_, _05510_);
  nor (_05654_, _05520_, _05518_);
  not (_05655_, _05633_);
  nor (_05656_, _05655_, _05627_);
  not (_05658_, _05597_);
  and (_05659_, _05603_, _05658_);
  not (_05661_, _05306_);
  and (_05662_, _05661_, _05150_);
  nor (_05663_, _05606_, _05662_);
  nor (_05664_, _05663_, _05659_);
  nor (_05666_, _05664_, _05636_);
  nor (_05667_, _05666_, _05656_);
  and (_05668_, _05664_, _05636_);
  nor (_05669_, _05668_, _05666_);
  not (_05671_, _05669_);
  and (_05672_, _05606_, _05662_);
  nor (_05673_, _05672_, _05663_);
  not (_05674_, _05673_);
  not (_05675_, _05309_);
  and (_05676_, _05550_, _05253_);
  or (_05677_, _05676_, _05554_);
  or (_05678_, _05543_, _05274_);
  and (_05679_, _05678_, _05677_);
  or (_05681_, _05679_, _05538_);
  not (_05682_, _05534_);
  or (_05683_, _05682_, _05233_);
  and (_05684_, _05683_, _05681_);
  nor (_05685_, _05684_, _05529_);
  and (_05686_, _05684_, _05529_);
  or (_05687_, _05686_, _05685_);
  and (_05689_, _05679_, _05538_);
  not (_05690_, _05689_);
  nand (_05692_, _05690_, _05681_);
  and (_05693_, _05676_, _05554_);
  not (_05694_, _05693_);
  nand (_05696_, _05694_, _05677_);
  nor (_05697_, _05563_, _05188_);
  and (_05699_, _05697_, _05696_);
  and (_05700_, _05699_, _05692_);
  and (_05702_, _05700_, _05687_);
  not (_05703_, _05526_);
  or (_05705_, _05703_, _05210_);
  and (_05707_, _05703_, _05210_);
  or (_05708_, _05684_, _05707_);
  and (_05710_, _05708_, _05705_);
  or (_05711_, _05710_, _05702_);
  and (_05713_, _05711_, _05675_);
  and (_05714_, _05713_, _05674_);
  and (_05715_, _05714_, _05671_);
  nor (_05716_, _05715_, _05667_);
  nor (_05717_, _05716_, _05654_);
  nor (_05718_, _05717_, _05653_);
  or (_05719_, _05718_, _05651_);
  and (_05720_, _05627_, _05597_);
  not (_05722_, _05720_);
  not (_05723_, _05150_);
  and (_05725_, _05325_, _05163_);
  and (_05726_, _05274_, _05233_);
  nor (_05728_, _05726_, _05210_);
  and (_05729_, _05728_, _05725_);
  and (_05731_, _05729_, _05723_);
  nor (_05732_, _05731_, _05722_);
  nor (_05734_, _05732_, _05510_);
  nor (_05735_, _05734_, _05187_);
  not (_05736_, _05735_);
  not (_05737_, _05725_);
  nor (_05738_, _05510_, _05188_);
  not (_05739_, _05738_);
  nor (_05740_, _05739_, _05732_);
  nor (_05741_, _05740_, _05737_);
  and (_05742_, _05741_, _05736_);
  not (_05743_, _05729_);
  and (_05744_, _05168_, _05325_);
  and (_05746_, _05280_, _05744_);
  and (_05747_, _05185_, _05181_);
  and (_05749_, _05171_, _05290_);
  and (_05751_, _05312_, _05185_);
  nor (_05752_, _05751_, _05749_);
  nor (_05753_, _05752_, _05747_);
  nor (_05754_, _05753_, _05746_);
  nor (_05755_, _05187_, _05185_);
  not (_05756_, _05295_);
  and (_05758_, _05187_, _05185_);
  or (_05759_, _05758_, _05756_);
  and (_05760_, _05759_, _05327_);
  or (_05761_, _05760_, _05755_);
  and (_05762_, _05171_, _05311_);
  not (_05763_, _05762_);
  nor (_05764_, _05510_, _05763_);
  nor (_05765_, _05314_, _05187_);
  and (_05766_, _05168_, _05157_);
  not (_05767_, _05185_);
  nand (_05768_, _05767_, _05766_);
  and (_05769_, _05768_, _05159_);
  and (_05770_, _05769_, _05187_);
  nor (_05771_, _05770_, _05765_);
  nor (_05773_, _05771_, _05764_);
  and (_05774_, _05773_, _05761_);
  and (_05776_, _05774_, _05754_);
  and (_05777_, _05776_, _05743_);
  not (_05778_, _05777_);
  nor (_05779_, _05778_, _05742_);
  and (_05781_, _05779_, _05719_);
  nand (_05782_, _05781_, _05649_);
  and (_05784_, _05782_, _05488_);
  and (_05785_, _05401_, _05375_);
  or (_05786_, _05376_, _05785_);
  and (_05787_, _05786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_05788_, _05787_, _05784_);
  and (_05789_, _05447_, _05433_);
  not (_05790_, _05341_);
  not (_05791_, _05336_);
  nor (_05792_, _05349_, _05791_);
  and (_05793_, _05792_, _05790_);
  and (_05794_, _05793_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_05795_, _05794_, _05390_);
  and (_05796_, _05795_, _05418_);
  and (_05797_, _05796_, _05460_);
  and (_05798_, _05797_, _05789_);
  and (_05799_, _05798_, _05788_);
  nand (_05800_, _05798_, _05375_);
  and (_05801_, _05800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_05802_, _05433_, _05418_);
  and (_05803_, _05460_, _05447_);
  and (_05804_, _05803_, _05802_);
  and (_05805_, _05376_, _05401_);
  and (_05806_, _05793_, _05335_);
  and (_05807_, _05806_, _05390_);
  and (_05808_, _05807_, _05805_);
  and (_05809_, _05808_, _05804_);
  or (_05810_, _05809_, _05801_);
  or (_05811_, _05810_, _05799_);
  nor (_05812_, _05633_, _05188_);
  nor (_05813_, _05627_, _05187_);
  or (_05814_, _05813_, _05812_);
  and (_05815_, _05814_, _05320_);
  not (_05816_, _05627_);
  or (_05817_, _05277_, _05723_);
  or (_05818_, _05658_, _05817_);
  nand (_05819_, _05818_, _05187_);
  or (_05820_, _05597_, _05150_);
  nor (_05821_, _05820_, _05284_);
  or (_05822_, _05821_, _05187_);
  and (_05823_, _05822_, _05819_);
  nand (_05824_, _05823_, _05816_);
  or (_05825_, _05823_, _05816_);
  and (_05826_, _05825_, _05291_);
  and (_05827_, _05826_, _05824_);
  nor (_05828_, _05827_, _05815_);
  nor (_05829_, _05627_, _05176_);
  not (_05830_, _05829_);
  and (_05831_, _05636_, _05295_);
  not (_05832_, _05831_);
  nor (_05833_, _05635_, _05327_);
  not (_05834_, _05833_);
  and (_05835_, _05634_, _05312_);
  and (_05836_, _05627_, _05314_);
  nor (_05837_, _05836_, _05835_);
  and (_05838_, _05837_, _05834_);
  and (_05839_, _05838_, _05832_);
  and (_05840_, _05839_, _05830_);
  and (_05841_, _05840_, _05828_);
  nand (_05842_, _05841_, _05809_);
  and (_05843_, _05842_, _05110_);
  and (_07249_, _05843_, _05811_);
  not (_05844_, _05809_);
  nor (_05845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_05846_, _05845_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not (_05847_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_05848_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_05849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_05850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_05851_, _05850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_05852_, _05851_, _05849_);
  nor (_05853_, _05852_, _05848_);
  or (_05854_, _05853_, _05847_);
  and (_05855_, _05850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_05856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_05857_, _05856_, _05855_);
  nor (_05858_, _05857_, _05848_);
  and (_05859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_05860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _05850_);
  nor (_05861_, _05860_, _05859_);
  nand (_05862_, _05861_, _05858_);
  or (_05863_, _05862_, _05854_);
  and (_05864_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_05865_, _05864_, _05846_);
  nor (_05866_, _05375_, _05365_);
  and (_05867_, _05866_, _05485_);
  and (_05868_, _05867_, _05804_);
  and (_05869_, _05868_, _05795_);
  or (_05870_, _05869_, _05865_);
  and (_05871_, _05870_, _05844_);
  and (_05872_, _05781_, _05649_);
  nand (_05873_, _05869_, _05872_);
  and (_05874_, _05873_, _05871_);
  and (_05875_, _05821_, _05816_);
  and (_05876_, _05875_, _05188_);
  nor (_05877_, _05722_, _05817_);
  and (_05878_, _05877_, _05187_);
  nor (_05879_, _05878_, _05876_);
  and (_05880_, _05879_, _05510_);
  not (_05881_, _05880_);
  not (_05882_, _05291_);
  nor (_05883_, _05879_, _05510_);
  nor (_05884_, _05883_, _05882_);
  and (_05885_, _05884_, _05881_);
  and (_05886_, _05510_, _05188_);
  not (_05887_, _05886_);
  and (_05888_, _05517_, _05187_);
  nor (_05889_, _05888_, _05321_);
  and (_05890_, _05889_, _05887_);
  nor (_05891_, _05890_, _05885_);
  and (_05892_, _05518_, _05312_);
  and (_05893_, _05510_, _05314_);
  nor (_05894_, _05893_, _05892_);
  nor (_05895_, _05510_, _05176_);
  and (_05896_, _05654_, _05295_);
  nor (_05897_, _05520_, _05327_);
  or (_05898_, _05897_, _05896_);
  nor (_05899_, _05898_, _05895_);
  and (_05900_, _05899_, _05894_);
  and (_05901_, _05900_, _05891_);
  nor (_05902_, _05901_, _05844_);
  or (_05903_, _05902_, _05874_);
  and (_07357_, _05903_, _05110_);
  not (_05904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_05905_, _05853_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor (_05906_, _05861_, _05848_);
  or (_05907_, _05906_, _05858_);
  or (_05908_, _05907_, _05905_);
  and (_05909_, _05908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_05910_, _05909_, _05904_);
  not (_05911_, _05375_);
  and (_05912_, _05911_, _05365_);
  and (_05913_, _05912_, _05402_);
  and (_05914_, _05804_, _05913_);
  and (_05915_, _05914_, _05794_);
  or (_05916_, _05915_, _05910_);
  and (_05917_, _05916_, _05844_);
  nand (_05918_, _05915_, _05872_);
  and (_05919_, _05918_, _05917_);
  and (_05920_, _05543_, _05320_);
  nor (_05921_, _05282_, _05275_);
  or (_05922_, _05921_, _05187_);
  nand (_05923_, _05921_, _05187_);
  and (_05924_, _05923_, _05291_);
  and (_05925_, _05924_, _05922_);
  nor (_05926_, _05925_, _05920_);
  or (_05927_, _05553_, _05327_);
  or (_05928_, _05553_, _05544_);
  or (_05929_, _05928_, _05756_);
  and (_05930_, _05929_, _05927_);
  nand (_05931_, _05544_, _05312_);
  not (_05932_, _05314_);
  or (_05933_, _05932_, _05281_);
  and (_05934_, _05933_, _05931_);
  or (_05935_, _05274_, _05176_);
  and (_05936_, _05935_, _05934_);
  and (_05937_, _05936_, _05930_);
  and (_05938_, _05937_, _05926_);
  nor (_05939_, _05938_, _05844_);
  or (_05940_, _05939_, _05919_);
  and (_07655_, _05940_, _05110_);
  and (_05941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _05848_);
  not (_05942_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_05943_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_05944_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_05945_, _05944_, _05943_);
  and (_05946_, _05945_, _05942_);
  not (_05947_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_05948_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_05949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_05950_, _05949_, _05948_);
  and (_05951_, _05950_, _05947_);
  nor (_05952_, _05951_, _05946_);
  not (_05953_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_05954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_05955_, _05954_, _05953_);
  not (_05956_, _05955_);
  not (_05957_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_05958_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_05959_, _05958_, _05957_);
  not (_05960_, _05959_);
  not (_05961_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_05962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_05963_, _05962_, _05961_);
  not (_05964_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_05965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_05966_, _05965_, _05964_);
  nor (_05967_, _05966_, _05963_);
  and (_05968_, _05967_, _05960_);
  and (_05969_, _05968_, _05956_);
  nand (_05970_, _05969_, _05952_);
  nand (_05971_, _05970_, _05941_);
  nand (_05972_, _05945_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_05973_, _05950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_05974_, _05973_);
  and (_05975_, _05974_, _05972_);
  and (_05976_, _05958_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_05977_, _05962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_05978_, _05977_, _05976_);
  and (_05979_, _05965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_05980_, _05954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_05981_, _05980_, _05979_);
  and (_05982_, _05981_, _05978_);
  and (_05983_, _05982_, _05975_);
  and (_05984_, _05983_, _05848_);
  nand (_05985_, _05984_, _05971_);
  and (_05986_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_05987_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05850_);
  nand (_05988_, _05987_, _05986_);
  and (_05989_, _05988_, _05110_);
  and (_07918_, _05989_, _05985_);
  and (_05990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _05110_);
  and (_08055_, _05990_, _05986_);
  and (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _05110_);
  and (_05991_, _05401_, _05389_);
  and (_05992_, _05991_, _05376_);
  and (_05993_, _05802_, _05461_);
  and (_05994_, _05993_, _05992_);
  not (_05995_, _05337_);
  and (_05996_, _05991_, _05912_);
  and (_05997_, _05993_, _05996_);
  nor (_05998_, _05997_, _05994_);
  and (_05999_, _05992_, _05462_);
  not (_06000_, _05999_);
  and (_06001_, _05913_, _05993_);
  and (_06002_, _05993_, _05403_);
  nor (_06003_, _06002_, _06001_);
  and (_06004_, _06003_, _06000_);
  and (_06005_, _06004_, _05998_);
  or (_06006_, _06005_, _05995_);
  or (_06007_, _06006_, _05994_);
  and (_06008_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_06009_, _05938_, _06000_);
  not (_06010_, _05997_);
  nand (_06011_, _06003_, _06010_);
  and (_06012_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or (_06014_, _06012_, _06009_);
  and (_06015_, _06014_, _05337_);
  or (_06016_, _06015_, _06008_);
  and (_08933_, _06016_, _05110_);
  not (_06017_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_06018_, _06017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not (_06019_, _05906_);
  or (_06020_, _06019_, _05858_);
  or (_06021_, _06020_, _05854_);
  and (_06022_, _06021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_06023_, _06022_, _06018_);
  nor (_06024_, _05401_, _05389_);
  and (_06025_, _06024_, _05912_);
  and (_06026_, _06025_, _05804_);
  and (_06027_, _06026_, _05794_);
  or (_06028_, _06027_, _06023_);
  and (_06029_, _06028_, _05844_);
  nand (_06030_, _06027_, _05872_);
  and (_06031_, _06030_, _06029_);
  nor (_06032_, _05597_, _05187_);
  nor (_06033_, _05603_, _05188_);
  or (_06034_, _06033_, _06032_);
  and (_06035_, _06034_, _05320_);
  nand (_06036_, _05817_, _05285_);
  and (_06037_, _06036_, _05319_);
  or (_06038_, _06037_, _05658_);
  nand (_06040_, _06037_, _05658_);
  and (_06041_, _06040_, _05291_);
  and (_06042_, _06041_, _06038_);
  nor (_06043_, _06042_, _06035_);
  nor (_06044_, _05597_, _05176_);
  not (_06045_, _06044_);
  and (_06046_, _05606_, _05295_);
  nor (_06047_, _05604_, _05327_);
  nor (_06048_, _06047_, _06046_);
  and (_06049_, _05605_, _05312_);
  and (_06050_, _05597_, _05314_);
  nor (_06051_, _06050_, _06049_);
  and (_06052_, _06051_, _06048_);
  and (_06053_, _06052_, _06045_);
  and (_06054_, _06053_, _06043_);
  nor (_06055_, _06054_, _05844_);
  or (_06056_, _06055_, _06031_);
  and (_08980_, _06056_, _05110_);
  and (_06057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_06058_, _06020_, _05905_);
  and (_06059_, _06058_, _06057_);
  and (_06061_, _05866_, _05402_);
  and (_06062_, _06061_, _05804_);
  and (_06063_, _06062_, _05794_);
  or (_06064_, _06063_, _06059_);
  and (_06065_, _06064_, _05844_);
  nand (_06066_, _06063_, _05872_);
  and (_06067_, _06066_, _06065_);
  nor (_06068_, _05210_, _05176_);
  not (_06069_, _06068_);
  nand (_06070_, _05276_, _05187_);
  nand (_06071_, _05283_, _05188_);
  and (_06072_, _06071_, _06070_);
  or (_06073_, _06072_, _05211_);
  nand (_06074_, _06072_, _05211_);
  and (_06075_, _06074_, _05291_);
  nand (_06076_, _06075_, _06073_);
  nand (_06077_, _05529_, _05295_);
  or (_06078_, _05528_, _05327_);
  and (_06079_, _05527_, _05312_);
  not (_06080_, _06079_);
  nor (_06081_, _05526_, _05321_);
  and (_06082_, _05314_, _05210_);
  nor (_06083_, _06082_, _06081_);
  and (_06084_, _06083_, _06080_);
  and (_06085_, _06084_, _06078_);
  and (_06086_, _06085_, _06077_);
  and (_06087_, _06086_, _06076_);
  and (_06088_, _06087_, _06069_);
  nor (_06089_, _06088_, _05844_);
  or (_06091_, _06089_, _06067_);
  and (_09243_, _06091_, _05110_);
  nor (_06092_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_06093_, _06092_);
  and (_06094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _05850_);
  and (_06095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_06096_, _06095_, _06094_);
  and (_06097_, _06096_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_06098_, _06097_, _05848_);
  nor (_06099_, _06098_, _05983_);
  nor (_06100_, _06099_, _05971_);
  not (_06101_, _06100_);
  or (_06102_, _06101_, _05968_);
  not (_06103_, _05976_);
  nor (_06104_, _05979_, _05977_);
  and (_06105_, _06104_, _06103_);
  or (_06106_, _06098_, _06105_);
  and (_06107_, _06106_, _06102_);
  or (_06108_, _06107_, _06093_);
  not (_06109_, _05952_);
  and (_06110_, _06109_, _05941_);
  and (_06111_, _05955_, _05941_);
  or (_06112_, _06111_, _06110_);
  or (_06113_, _06112_, _06099_);
  not (_06114_, _05980_);
  and (_06115_, _06114_, _05975_);
  nand (_06116_, _06099_, _06115_);
  and (_06117_, _06116_, _06113_);
  and (_06118_, _06117_, _06092_);
  or (_06119_, _06118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_06120_, _06119_, _05110_);
  and (_10256_, _06120_, _06108_);
  not (_06121_, _05433_);
  and (_06122_, _05447_, _06121_);
  and (_06123_, _06122_, _05797_);
  and (_06124_, _06123_, _05867_);
  nand (_06125_, _06124_, _05872_);
  or (_06126_, _06124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_06127_, _06121_, _05418_);
  and (_06128_, _06127_, _05803_);
  and (_06129_, _06128_, _05808_);
  not (_06130_, _06129_);
  and (_06131_, _06130_, _06126_);
  and (_06132_, _06131_, _06125_);
  nor (_06134_, _06130_, _05901_);
  or (_06135_, _06134_, _06132_);
  and (_10306_, _06135_, _05110_);
  and (_06136_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_06137_, _05986_);
  and (_06138_, _06107_, _06137_);
  or (_06139_, _06138_, _06092_);
  and (_06140_, _06117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_06141_, _06140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_06142_, _06141_, _06139_);
  or (_06143_, _06142_, _06136_);
  and (_10385_, _06143_, _05110_);
  nor (_06144_, _05433_, _05418_);
  and (_06145_, _06144_, _05803_);
  and (_06146_, _05806_, _05389_);
  and (_06147_, _06146_, _05867_);
  and (_06148_, _06147_, _06145_);
  not (_06149_, _06148_);
  and (_06150_, _05794_, _05460_);
  nor (_06151_, _05418_, _05389_);
  and (_06152_, _06151_, _06150_);
  and (_06153_, _06152_, _06122_);
  and (_06154_, _06153_, _05867_);
  or (_06155_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_06156_, _06155_, _06149_);
  nand (_06157_, _06154_, _05872_);
  and (_06158_, _06157_, _06156_);
  nor (_06159_, _06149_, _05901_);
  or (_06160_, _06159_, _06158_);
  and (_10406_, _06160_, _05110_);
  or (_06161_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not (_06162_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_06163_, pc_log_change, _06162_);
  and (_06164_, _06163_, _05110_);
  and (_10427_, _06164_, _06161_);
  and (_06165_, _05913_, _05462_);
  not (_06166_, _06165_);
  nor (_06167_, _06166_, _05334_);
  not (_06168_, _05463_);
  and (_06169_, _05996_, _05462_);
  nor (_06170_, _05999_, _06169_);
  and (_06171_, _06170_, _06168_);
  and (_06172_, _06171_, _06166_);
  and (_06173_, _05401_, _05365_);
  and (_06174_, _05993_, _06173_);
  or (_06175_, _06174_, _05995_);
  nor (_06176_, _06175_, _06172_);
  nand (_06177_, _06176_, _06171_);
  and (_06178_, _06177_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_06179_, _06178_, _06167_);
  or (_06180_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_06182_, _06180_, _05110_);
  and (_12614_, _06182_, _06179_);
  not (_06183_, _06054_);
  and (_06184_, _06165_, _05337_);
  and (_06185_, _06184_, _06183_);
  or (_06186_, _06172_, _05995_);
  and (_06187_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand (_06188_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_06189_, _06188_, _06171_);
  or (_06190_, _06189_, _06187_);
  or (_06191_, _06190_, _06185_);
  and (_12886_, _06191_, _05110_);
  and (_06193_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  not (_06194_, _06088_);
  and (_06195_, _06184_, _06194_);
  nand (_06196_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_06197_, _06196_, _06171_);
  or (_06198_, _06197_, _06195_);
  or (_06199_, _06198_, _06193_);
  and (_12945_, _06199_, _05110_);
  not (_06200_, _05474_);
  not (_06201_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_06202_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_06203_, _06202_, _06201_);
  nor (_06204_, _06203_, _06200_);
  nor (_06205_, _06204_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_06206_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not (_06207_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_06208_, _06205_, _06207_);
  and (_06209_, _06208_, _05110_);
  and (_13108_, _06209_, _06206_);
  and (_06210_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_06211_, _05282_, _05187_);
  or (_06212_, _05275_, _05188_);
  and (_06213_, _06212_, _06211_);
  or (_06214_, _06213_, _05279_);
  nand (_06215_, _06213_, _05279_);
  and (_06216_, _06215_, _05291_);
  and (_06217_, _06216_, _06214_);
  nor (_06218_, _05534_, _05321_);
  nor (_06219_, _06218_, _06217_);
  and (_06220_, _05535_, _05312_);
  and (_06221_, _05314_, _05233_);
  nor (_06222_, _06221_, _06220_);
  nor (_06223_, _05233_, _05176_);
  and (_06224_, _05538_, _05295_);
  nor (_06225_, _05537_, _05327_);
  or (_06226_, _06225_, _06224_);
  nor (_06227_, _06226_, _06223_);
  and (_06228_, _06227_, _06222_);
  and (_06229_, _06228_, _06219_);
  not (_06230_, _06229_);
  and (_06231_, _06230_, _06184_);
  nand (_06232_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_06233_, _06232_, _06171_);
  or (_06234_, _06233_, _06231_);
  or (_06235_, _06234_, _06210_);
  and (_13173_, _06235_, _05110_);
  and (_06237_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_06238_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_06239_, \oc8051_top_1.oc8051_decoder1.state [0], _05151_);
  and (_06240_, _06239_, _06238_);
  not (_06241_, _05475_);
  nor (_06242_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_06243_, _06242_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_06244_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_06245_, _06202_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_06246_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_06247_, _06246_, _06244_);
  not (_06248_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  not (_06249_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_06250_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _06201_);
  nand (_06251_, _06250_, _06249_);
  or (_06252_, _06251_, _06248_);
  and (_06253_, _06252_, _06247_);
  not (_06254_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_06255_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_06256_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], _06255_);
  and (_06257_, _06256_, _06201_);
  nand (_06258_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_06259_, _06258_, _06254_);
  nor (_06260_, _06242_, _06201_);
  nand (_06261_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_06262_, _06242_, _06201_);
  nand (_06263_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_06264_, _06263_, _06261_);
  and (_06265_, _06264_, _06259_);
  nand (_06266_, _06265_, _06253_);
  or (_06267_, _06266_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_06268_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_06269_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  not (_06270_, _06269_);
  and (_06271_, _06270_, _06267_);
  or (_06272_, _06271_, _06241_);
  not (_06273_, _05472_);
  nor (_06274_, _05474_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_06275_, _06274_, _06273_);
  and (_06276_, _06275_, _06272_);
  not (_06277_, _06276_);
  nand (_06278_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_06279_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_06280_, _06279_, _06278_);
  nand (_06281_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_06282_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_06283_, _06282_, _06281_);
  nand (_06284_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  not (_06285_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_06286_, _06251_, _06285_);
  and (_06287_, _06286_, _06284_);
  and (_06288_, _06287_, _06283_);
  and (_06289_, _06288_, _06280_);
  or (_06290_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_06291_, _06290_, _06289_);
  and (_06292_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not (_06293_, _06292_);
  and (_06294_, _06293_, _06291_);
  nand (_06295_, _06294_, _05475_);
  nor (_06296_, _05474_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_06297_, _06296_, _06273_);
  and (_06298_, _06297_, _06295_);
  nand (_06300_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_06301_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_06302_, _06301_, _06300_);
  nand (_06303_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_06304_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_06305_, _06304_, _06303_);
  nand (_06306_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not (_06307_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_06308_, _06251_, _06307_);
  and (_06309_, _06308_, _06306_);
  and (_06310_, _06309_, _06305_);
  and (_06311_, _06310_, _06302_);
  or (_06312_, _06311_, _06290_);
  and (_06313_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_06314_, _06313_);
  and (_06315_, _06314_, _06312_);
  nand (_06316_, _06315_, _05475_);
  nor (_06317_, _05474_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_06318_, _06317_, _06273_);
  and (_06319_, _06318_, _06316_);
  not (_06320_, _06319_);
  and (_06321_, _06320_, _06298_);
  nor (_06322_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_06323_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_06324_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_06325_, _06324_, _06323_);
  nand (_06326_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_06327_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_06328_, _06327_, _06326_);
  nand (_06329_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not (_06330_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_06331_, _06251_, _06330_);
  and (_06332_, _06331_, _06329_);
  and (_06333_, _06332_, _06328_);
  nand (_06334_, _06333_, _06325_);
  nand (_06335_, _06334_, _06322_);
  and (_06336_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not (_06337_, _06336_);
  and (_06338_, _06337_, _06335_);
  nand (_06339_, _06338_, _05475_);
  nor (_06340_, _05474_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_06341_, _06340_, _06273_);
  and (_06342_, _06341_, _06339_);
  and (_06343_, _06342_, _06321_);
  and (_06344_, _06343_, _06277_);
  nand (_06345_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand (_06346_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_06347_, _06346_, _06345_);
  nand (_06348_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_06349_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_06350_, _06349_, _06348_);
  nand (_06351_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  not (_06352_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_06353_, _06251_, _06352_);
  and (_06354_, _06353_, _06351_);
  and (_06355_, _06354_, _06350_);
  nand (_06356_, _06355_, _06347_);
  nand (_06357_, _06356_, _06254_);
  nand (_06358_, _06357_, _06268_);
  nor (_06359_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  not (_06360_, _06359_);
  and (_06362_, _06360_, _06358_);
  or (_06363_, _06362_, _06241_);
  nor (_06364_, _05474_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_06365_, _06364_, _06273_);
  and (_06366_, _06365_, _06363_);
  nand (_06367_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_06368_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_06369_, _06368_, _06367_);
  not (_06370_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_06371_, _06251_, _06370_);
  and (_06373_, _06371_, _06369_);
  nand (_06374_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_06375_, _06374_, _06254_);
  nand (_06376_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_06377_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_06378_, _06377_, _06376_);
  and (_06379_, _06378_, _06375_);
  nand (_06380_, _06379_, _06373_);
  or (_06381_, _06380_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_06382_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  not (_06383_, _06382_);
  and (_06384_, _06383_, _06381_);
  or (_06385_, _06384_, _06241_);
  nor (_06386_, _05474_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_06387_, _06386_, _06273_);
  and (_06388_, _06387_, _06385_);
  nor (_06389_, _06388_, _06366_);
  nand (_06390_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand (_06391_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_06392_, _06391_, _06390_);
  nand (_06393_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_06394_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_06395_, _06394_, _06393_);
  nand (_06396_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  not (_06397_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_06398_, _06251_, _06397_);
  and (_06399_, _06398_, _06396_);
  and (_06400_, _06399_, _06395_);
  nand (_06401_, _06400_, _06392_);
  nand (_06402_, _06401_, _06254_);
  nand (_06403_, _06402_, _06268_);
  nor (_06404_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  not (_06405_, _06404_);
  and (_06406_, _06405_, _06403_);
  or (_06407_, _06406_, _06241_);
  nor (_06409_, _05474_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_06410_, _06409_, _06273_);
  and (_06411_, _06410_, _06407_);
  nand (_06412_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not (_06413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_06414_, _06251_, _06413_);
  and (_06415_, _06414_, _06412_);
  nand (_06416_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand (_06417_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_06418_, _06417_, _06416_);
  nand (_06419_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_06420_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_06421_, _06420_, _06419_);
  and (_06422_, _06421_, _06418_);
  and (_06423_, _06422_, _06415_);
  or (_06424_, _06423_, _06290_);
  and (_06425_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  not (_06426_, _06425_);
  and (_06427_, _06426_, _06424_);
  nand (_06428_, _06427_, _05475_);
  nor (_06429_, _05474_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_06430_, _06429_, _06273_);
  and (_06431_, _06430_, _06428_);
  not (_06432_, _06431_);
  and (_06433_, _06432_, _06411_);
  and (_06434_, _06433_, _06389_);
  and (_06435_, _06434_, _06344_);
  not (_06436_, _06342_);
  and (_06437_, _06436_, _06321_);
  and (_06438_, _06437_, _06277_);
  and (_06439_, _06438_, _06434_);
  nor (_06440_, _06439_, _06435_);
  not (_06442_, _06440_);
  and (_06443_, _06442_, _06240_);
  or (_06444_, _06443_, _06237_);
  not (_06445_, _06388_);
  nor (_06446_, _06411_, _06445_);
  and (_06447_, _06446_, _06432_);
  and (_06448_, _06447_, _06366_);
  and (_06449_, _06448_, _06344_);
  nor (_06450_, _06431_, _06411_);
  and (_06451_, _06450_, _06389_);
  and (_06452_, _06437_, _06276_);
  and (_06453_, _06452_, _06451_);
  or (_06454_, _06453_, _06449_);
  nor (_06455_, _06432_, _06276_);
  and (_06456_, _06436_, _06319_);
  and (_06457_, _06456_, _06455_);
  and (_06458_, _06457_, _06298_);
  and (_06459_, _06456_, _06298_);
  and (_06460_, _06433_, _06388_);
  and (_06461_, _06460_, _06459_);
  or (_06462_, _06461_, _06458_);
  and (_06463_, _06459_, _06277_);
  and (_06464_, _06433_, _06445_);
  and (_06465_, _06464_, _06463_);
  or (_06466_, _06465_, _06462_);
  or (_06467_, _06466_, _06454_);
  and (_06468_, _06467_, _05474_);
  or (_06469_, _06468_, _06444_);
  and (_01001_, _06469_, _05110_);
  and (_06470_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05151_);
  and (_06471_, _06470_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_06472_, _05785_, _05486_);
  and (_06473_, _05804_, _06472_);
  and (_06475_, _06473_, _06146_);
  nor (_06476_, _06475_, _06471_);
  not (_06477_, _06476_);
  or (_06478_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_06479_, _05697_, _05696_);
  nor (_06480_, _06479_, _05699_);
  nor (_06481_, _06480_, _05651_);
  not (_06482_, _06481_);
  or (_06483_, _05233_, _05169_);
  and (_06485_, _05157_, _05163_);
  and (_06486_, _06485_, ABINPUT000000[2]);
  and (_06487_, _05311_, _05154_);
  and (_06488_, _06487_, ABINPUT000[2]);
  nor (_06489_, _06488_, _06486_);
  and (_06490_, _06489_, _06483_);
  and (_06491_, _05281_, _05158_);
  and (_06492_, _05280_, _05172_);
  nor (_06493_, _06492_, _06491_);
  and (_06494_, _06493_, _06490_);
  and (_06495_, _06494_, _05934_);
  and (_06496_, _06495_, _05930_);
  and (_06497_, _06496_, _05926_);
  nor (_06498_, _05728_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_06499_, _06498_, _05281_);
  nor (_06500_, _06498_, _05281_);
  nor (_06501_, _06500_, _06499_);
  nor (_06502_, _06501_, _05737_);
  or (_06503_, _05549_, _05253_);
  and (_06504_, _05928_, _06503_);
  or (_06505_, _06504_, _05555_);
  and (_06506_, _06505_, _05564_);
  nor (_06507_, _06505_, _05564_);
  or (_06508_, _06507_, _06506_);
  and (_06509_, _06508_, _05489_);
  nor (_06510_, _06509_, _06502_);
  and (_06511_, _06510_, _06497_);
  and (_06512_, _06511_, _06482_);
  nand (_06513_, _06512_, _06477_);
  and (_06514_, _06513_, _05110_);
  and (_01593_, _06514_, _06478_);
  nor (_06515_, _05713_, _05674_);
  nor (_06516_, _06515_, _05714_);
  nor (_06517_, _06516_, _05651_);
  not (_06518_, _06517_);
  nor (_06519_, _05606_, _05307_);
  or (_06520_, _06519_, _05638_);
  and (_06521_, _06520_, _05576_);
  nor (_06522_, _06521_, _05490_);
  and (_06523_, _06522_, _05608_);
  nor (_06524_, _05597_, _05159_);
  and (_06525_, _06485_, ABINPUT000000[6]);
  nor (_06526_, _06525_, _06524_);
  and (_06528_, _06526_, _06052_);
  nor (_06529_, _05720_, _05510_);
  nor (_06530_, _06529_, _05187_);
  and (_06531_, _06530_, _05743_);
  nor (_06532_, _06531_, _05731_);
  and (_06533_, _06532_, _05597_);
  nor (_06534_, _06532_, _05597_);
  nor (_06535_, _06534_, _06533_);
  nor (_06536_, _06535_, _05737_);
  nor (_06537_, _05174_, _05150_);
  or (_06538_, _05627_, _05169_);
  and (_06539_, _06487_, ABINPUT000[6]);
  not (_06540_, _06539_);
  nand (_06541_, _06540_, _06538_);
  or (_06542_, _06541_, _06537_);
  nor (_06543_, _06542_, _06536_);
  and (_06544_, _06543_, _06528_);
  and (_06545_, _06544_, _06043_);
  not (_06546_, _06545_);
  nor (_06547_, _06546_, _06523_);
  and (_06548_, _06547_, _06518_);
  nand (_06549_, _06548_, _06477_);
  or (_06550_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_06551_, _06550_, _05110_);
  and (_01615_, _06551_, _06549_);
  not (_06552_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  not (_06553_, _06002_);
  and (_06554_, _06553_, _05998_);
  nor (_06555_, _06554_, _05995_);
  nor (_06556_, _06555_, _06552_);
  nand (_06557_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_06558_, _06557_, _05998_);
  not (_06559_, _05938_);
  and (_06560_, _06002_, _05337_);
  and (_06561_, _06560_, _06559_);
  or (_06562_, _06561_, _06558_);
  or (_06563_, _06562_, _06556_);
  and (_03222_, _06563_, _05110_);
  nand (_06564_, _05647_, _05519_);
  nor (_06565_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_06566_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05240_);
  nor (_06567_, _06566_, _06565_);
  and (_06568_, _06567_, _06564_);
  nor (_06569_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_06570_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05264_);
  nor (_06571_, _06570_, _06569_);
  and (_06572_, _06571_, _06568_);
  nor (_06573_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_06574_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05218_);
  nor (_06575_, _06574_, _06573_);
  and (_06576_, _06575_, _06572_);
  nor (_06577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06578_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05195_);
  nor (_06579_, _06578_, _06577_);
  or (_06580_, _06579_, _06576_);
  nand (_06581_, _06579_, _06576_);
  and (_06582_, _06581_, _05489_);
  nand (_06583_, _06582_, _06580_);
  and (_06584_, _05877_, _05510_);
  and (_06585_, _06584_, _05549_);
  and (_06586_, _06585_, _05552_);
  and (_06587_, _05534_, _05187_);
  and (_06588_, _06587_, _06586_);
  nor (_06589_, _05549_, _05510_);
  and (_06590_, _06589_, _05875_);
  and (_06591_, _06590_, _05543_);
  nor (_06592_, _05534_, _05187_);
  and (_06593_, _06592_, _06591_);
  nor (_06594_, _06593_, _06588_);
  and (_06595_, _06594_, _05526_);
  not (_06596_, _06595_);
  nor (_06597_, _06594_, _05526_);
  nor (_06598_, _06597_, _05882_);
  and (_06599_, _06598_, _06596_);
  and (_06600_, _06485_, ABINPUT000000[12]);
  and (_06601_, _06487_, ABINPUT000[12]);
  nor (_06602_, _06601_, _06600_);
  nor (_06603_, _05321_, _05210_);
  nor (_06604_, _05526_, _05159_);
  or (_06605_, _06604_, _06603_);
  nor (_06606_, _06605_, _05764_);
  and (_06607_, _06606_, _06602_);
  not (_06608_, _06607_);
  nor (_06609_, _06608_, _06599_);
  nand (_06610_, _06609_, _06583_);
  not (_06611_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_06612_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05151_);
  and (_06613_, _06612_, _06611_);
  nand (_06615_, _06613_, _06610_);
  not (_06616_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_06617_, _06470_, _06616_);
  and (_06618_, _05460_, _05448_);
  and (_06619_, _06618_, _06127_);
  and (_06620_, _06619_, _05992_);
  and (_06621_, _06620_, _05806_);
  nor (_06622_, _06621_, _06617_);
  not (_06623_, _06622_);
  and (_06624_, _05460_, _05389_);
  and (_06625_, _06624_, _05418_);
  nor (_06626_, _05447_, _05433_);
  and (_06627_, _06626_, _05794_);
  and (_06628_, _06627_, _06625_);
  nor (_06629_, _06628_, _05204_);
  nor (_06630_, _06629_, _06623_);
  and (_06631_, _05866_, _05401_);
  and (_06632_, _06631_, _05782_);
  nor (_06633_, _06631_, _05204_);
  or (_06634_, _06633_, _06632_);
  nand (_06635_, _06634_, _06628_);
  and (_06636_, _06635_, _06630_);
  not (_06637_, _06613_);
  and (_06638_, _06622_, _06637_);
  nor (_06639_, _05700_, _05687_);
  nor (_06640_, _06639_, _05702_);
  nor (_06641_, _06640_, _05651_);
  not (_06642_, _06641_);
  nor (_06643_, _05570_, _05561_);
  or (_06644_, _06643_, _05490_);
  nor (_06645_, _06644_, _05571_);
  not (_06646_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_06647_, _05726_, _06646_);
  nor (_06648_, _06647_, _05211_);
  nor (_06649_, _05728_, _05737_);
  not (_06650_, _06649_);
  nor (_06651_, _06650_, _06648_);
  nor (_06652_, _05233_, _05174_);
  and (_06653_, _06485_, ABINPUT000000[4]);
  and (_06654_, _06487_, ABINPUT000[4]);
  nor (_06655_, _06654_, _06653_);
  not (_06656_, _06655_);
  nor (_06657_, _06656_, _06652_);
  or (_06658_, _05169_, _05150_);
  nor (_06659_, _05210_, _05159_);
  not (_06660_, _06659_);
  and (_06661_, _06660_, _06658_);
  and (_06662_, _06661_, _06657_);
  not (_06663_, _06662_);
  nor (_06664_, _06663_, _06651_);
  and (_06665_, _06664_, _06087_);
  not (_06666_, _06665_);
  nor (_06667_, _06666_, _06645_);
  and (_06668_, _06667_, _06642_);
  nor (_06669_, _06668_, _06613_);
  nor (_06670_, _06669_, _06638_);
  or (_06671_, _06670_, _06636_);
  nand (_06672_, _06671_, _06615_);
  and (_03832_, _06672_, _05110_);
  and (_06673_, _05994_, _05337_);
  nand (_06674_, _06673_, _06088_);
  or (_06675_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_06676_, _06675_, _05110_);
  and (_03950_, _06676_, _06674_);
  nand (_06677_, _06673_, _06054_);
  or (_06678_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_06679_, _06678_, _05110_);
  and (_04296_, _06679_, _06677_);
  nor (_06680_, _06010_, _05334_);
  and (_06681_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_06682_, _06681_, _05995_);
  or (_06683_, _06682_, _06680_);
  or (_06685_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_06686_, _06685_, _05110_);
  and (_04377_, _06686_, _06683_);
  nand (_06687_, _06673_, _05334_);
  or (_06688_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_06689_, _06688_, _05110_);
  and (_05107_, _06689_, _06687_);
  nand (_06690_, _06560_, _06229_);
  or (_06691_, _06560_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_06692_, _06691_, _05110_);
  and (_05108_, _06692_, _06690_);
  and (_06693_, _06579_, _06576_);
  nor (_06694_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06695_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05581_);
  nor (_06696_, _06695_, _06694_);
  nor (_06697_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06698_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05123_);
  nor (_06699_, _06698_, _06697_);
  and (_06700_, _06699_, _06696_);
  and (_06701_, _06700_, _06693_);
  nor (_06702_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_06703_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05613_);
  nor (_06704_, _06703_, _06702_);
  or (_06705_, _06704_, _06701_);
  nand (_06706_, _06704_, _06701_);
  and (_06707_, _06706_, _05489_);
  nand (_06708_, _06707_, _06705_);
  not (_06709_, _05510_);
  and (_06710_, _05875_, _06709_);
  and (_06711_, _06710_, _05550_);
  and (_06712_, _06711_, _05543_);
  and (_06713_, _06712_, _05682_);
  and (_06714_, _06713_, _05703_);
  and (_06716_, _06714_, _05661_);
  nor (_06717_, _06716_, _05187_);
  and (_06718_, _06586_, _05534_);
  and (_06719_, _06718_, _05526_);
  and (_06720_, _06719_, _05306_);
  nor (_06721_, _06720_, _05188_);
  or (_06722_, _06721_, _06717_);
  and (_06723_, _05603_, _05188_);
  nor (_06724_, _06723_, _06033_);
  not (_06725_, _06724_);
  nor (_06726_, _06725_, _06722_);
  and (_06727_, _06726_, _05655_);
  or (_06728_, _06726_, _05655_);
  nand (_06729_, _06728_, _05291_);
  or (_06730_, _06729_, _06727_);
  and (_06731_, _06487_, ABINPUT000[15]);
  and (_06732_, _05627_, _05187_);
  not (_06733_, _06732_);
  and (_06734_, _05633_, _05188_);
  nor (_06735_, _06734_, _05321_);
  and (_06736_, _06735_, _06733_);
  nor (_06737_, _05233_, _05763_);
  nor (_06738_, _05633_, _05159_);
  and (_06739_, _06485_, ABINPUT000000[15]);
  or (_06740_, _06739_, _06738_);
  or (_06741_, _06740_, _06737_);
  or (_06742_, _06741_, _06736_);
  nor (_06743_, _06742_, _06731_);
  and (_06744_, _06743_, _06730_);
  nand (_06745_, _06744_, _06708_);
  and (_06746_, _06745_, _06613_);
  and (_06747_, _06628_, _05488_);
  nor (_06748_, _06747_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_06749_, _06748_);
  and (_06750_, _06749_, _06638_);
  nand (_06751_, _06747_, _05872_);
  and (_06752_, _06751_, _06750_);
  and (_06753_, _05643_, _05608_);
  not (_06754_, _06753_);
  and (_06755_, _05644_, _05489_);
  and (_06756_, _06755_, _06754_);
  not (_06757_, _06756_);
  nor (_06758_, _05714_, _05671_);
  nor (_06759_, _06758_, _05715_);
  nor (_06760_, _06759_, _05651_);
  nor (_06761_, _06533_, _05627_);
  and (_06762_, _06533_, _05627_);
  nor (_06763_, _06762_, _06761_);
  nor (_06764_, _06763_, _05737_);
  or (_06765_, _05510_, _05169_);
  and (_06766_, _06485_, ABINPUT000000[7]);
  and (_06767_, _06487_, ABINPUT000[7]);
  nor (_06768_, _06767_, _06766_);
  and (_06769_, _06768_, _06765_);
  nor (_06770_, _05627_, _05159_);
  nor (_06771_, _05597_, _05174_);
  nor (_06772_, _06771_, _06770_);
  and (_06773_, _06772_, _06769_);
  and (_06774_, _06773_, _05839_);
  not (_06775_, _06774_);
  nor (_06776_, _06775_, _06764_);
  and (_06777_, _06776_, _05828_);
  not (_06778_, _06777_);
  nor (_06779_, _06778_, _06760_);
  and (_06780_, _06779_, _06757_);
  nor (_06781_, _06780_, _06622_);
  or (_06783_, _06781_, _06752_);
  and (_06784_, _06783_, _06637_);
  or (_06785_, _06784_, _06746_);
  and (_05109_, _06785_, _05110_);
  or (_06786_, _05551_, _05756_);
  and (_06787_, _06786_, _05327_);
  or (_06788_, _06787_, _05562_);
  nand (_06789_, _05551_, _05312_);
  or (_06790_, _05932_, _05280_);
  and (_06791_, _06790_, _06789_);
  or (_06792_, _05549_, _05321_);
  or (_06793_, _05882_, _05280_);
  and (_06794_, _06793_, _06792_);
  or (_06795_, _05253_, _05176_);
  and (_06796_, _06795_, _06794_);
  and (_06797_, _06796_, _06791_);
  and (_06798_, _06797_, _06788_);
  not (_06799_, _06798_);
  and (_06800_, _06799_, _05463_);
  not (_06801_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_06802_, _05464_, _06801_);
  or (_06803_, _06802_, _06800_);
  or (_06804_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_06805_, _06804_, _05110_);
  and (_05173_, _06805_, _06803_);
  and (_06807_, \oc8051_top_1.oc8051_sfr1.wait_data , _05110_);
  and (_06808_, _06807_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_06809_, _06445_, _06366_);
  and (_06810_, _06809_, _06433_);
  and (_06811_, _06459_, _06276_);
  and (_06812_, _06811_, _06810_);
  nor (_06813_, _06319_, _06298_);
  and (_06814_, _06813_, _06436_);
  and (_06815_, _06814_, _06277_);
  and (_06816_, _06815_, _06434_);
  and (_06817_, _06815_, _06810_);
  or (_06818_, _06817_, _06816_);
  or (_06819_, _06818_, _06812_);
  and (_06820_, _06814_, _06276_);
  and (_06821_, _06820_, _06464_);
  or (_06822_, _06821_, _06819_);
  and (_06823_, _06814_, _06460_);
  and (_06824_, _06342_, _06276_);
  and (_06825_, _06824_, _06321_);
  and (_06826_, _06411_, _06388_);
  or (_06827_, _06826_, _06431_);
  and (_06828_, _06827_, _06825_);
  nor (_06829_, _06828_, _06823_);
  and (_06830_, _06431_, _06276_);
  or (_06831_, _06814_, _06459_);
  and (_06832_, _06831_, _06830_);
  and (_06833_, _06814_, _06455_);
  nor (_06834_, _06833_, _06832_);
  nand (_06835_, _06834_, _06829_);
  and (_06836_, _06825_, _06434_);
  and (_06837_, _06452_, _06434_);
  or (_06838_, _06837_, _06836_);
  or (_06839_, _06838_, _06454_);
  or (_06840_, _06839_, _06835_);
  or (_06841_, _06840_, _06822_);
  and (_06842_, _05474_, _05110_);
  and (_06843_, _06842_, _06841_);
  or (_05179_, _06843_, _06808_);
  and (_06844_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06845_, _06810_, _06438_);
  and (_06846_, _06845_, _05474_);
  or (_06847_, _06846_, _06844_);
  or (_06848_, _06847_, _06443_);
  and (_05205_, _06848_, _05110_);
  and (_06849_, _06448_, _06437_);
  not (_06850_, _06849_);
  and (_06851_, _06342_, _06319_);
  and (_06852_, _06851_, _06298_);
  and (_06853_, _06852_, _06451_);
  and (_06854_, _06853_, _06277_);
  and (_06856_, _06852_, _06277_);
  and (_06857_, _06856_, _06447_);
  nor (_06858_, _06857_, _06854_);
  nand (_06859_, _06858_, _06850_);
  and (_06860_, _06859_, _06240_);
  or (_06861_, _06860_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06862_, _06448_, _06438_);
  nor (_06863_, _06431_, _06366_);
  and (_06864_, _06863_, _06446_);
  and (_06865_, _06864_, _06820_);
  and (_06866_, _06809_, _06450_);
  and (_06867_, _06866_, _06276_);
  or (_06868_, _06867_, _06865_);
  or (_06869_, _06868_, _06862_);
  or (_06870_, _05473_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_06871_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_06872_, \oc8051_top_1.oc8051_decoder1.state [1], _05151_);
  and (_06873_, _06872_, _06871_);
  and (_06874_, _06868_, _06873_);
  or (_06875_, _06874_, _06870_);
  and (_06876_, _06875_, _06869_);
  or (_06877_, _06876_, _06861_);
  or (_06878_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05151_);
  and (_06879_, _06878_, _05110_);
  and (_05208_, _06879_, _06877_);
  and (_06880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_06881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_06882_, _06881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_06883_, _06882_, _06880_);
  or (_06884_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not (_06885_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_06886_, _06883_, _06885_);
  and (_06887_, _06886_, _06884_);
  and (_06888_, _06618_, _05802_);
  and (_06889_, _05807_, _06472_);
  and (_06890_, _06889_, _06888_);
  or (_06891_, _06890_, _06887_);
  nand (_06892_, _06890_, _06798_);
  and (_06893_, _06892_, _06891_);
  and (_06894_, _06631_, _05807_);
  and (_06895_, _06894_, _06888_);
  or (_06896_, _06895_, _06893_);
  not (_06897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_06898_, _06895_, _06897_);
  and (_06899_, _06898_, _05110_);
  and (_05216_, _06899_, _06896_);
  and (_06901_, _05999_, _05337_);
  and (_06902_, _06183_, _06901_);
  and (_06903_, _06174_, _05337_);
  or (_06904_, _06903_, _06006_);
  and (_06905_, _06904_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_06906_, _06905_, _06902_);
  and (_05289_, _06906_, _05110_);
  and (_06907_, _05472_, _05151_);
  and (_06908_, _06907_, _06871_);
  not (_06909_, _06338_);
  and (_06910_, _06315_, _06294_);
  and (_06911_, _06910_, _06909_);
  not (_06912_, _06362_);
  not (_06913_, _06406_);
  and (_06914_, _06427_, _06384_);
  and (_06915_, _06914_, _06913_);
  and (_06916_, _06915_, _06912_);
  and (_06917_, _06916_, _06911_);
  not (_06918_, _06294_);
  and (_06920_, _06315_, _06918_);
  and (_06921_, _06920_, _06338_);
  and (_06922_, _06915_, _06362_);
  and (_06923_, _06922_, _06921_);
  not (_06924_, _06427_);
  nor (_06925_, _06924_, _06384_);
  and (_06926_, _06925_, _06406_);
  and (_06927_, _06926_, _06912_);
  not (_06928_, _06271_);
  and (_06929_, _06920_, _06928_);
  and (_06930_, _06929_, _06927_);
  or (_06931_, _06930_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_06932_, _06931_, _06923_);
  or (_06933_, _06932_, _06917_);
  and (_06934_, _06933_, _06908_);
  nor (_06935_, _06907_, _06871_);
  or (_06936_, _06935_, rst);
  or (_05315_, _06936_, _06934_);
  and (_06937_, _06807_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_06938_, _06864_, _06811_);
  and (_06939_, _06811_, _06448_);
  or (_06940_, _06939_, _06938_);
  and (_06941_, _06864_, _06343_);
  or (_06942_, _06941_, _06458_);
  or (_06943_, _06942_, _06940_);
  or (_06944_, _06832_, _06812_);
  or (_06945_, _06944_, _06449_);
  or (_06946_, _06820_, _06463_);
  and (_06947_, _06820_, _06434_);
  or (_06948_, _06810_, _06460_);
  or (_06949_, _06948_, _06947_);
  and (_06950_, _06949_, _06946_);
  or (_06951_, _06950_, _06945_);
  or (_06952_, _06951_, _06943_);
  and (_06953_, _06952_, _06842_);
  or (_05331_, _06953_, _06937_);
  not (_06954_, _06842_);
  nor (_06955_, _06853_, _06849_);
  or (_05342_, _06955_, _06954_);
  nor (_06956_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_06957_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05496_);
  nor (_06958_, _06957_, _06956_);
  or (_06959_, _06958_, _06706_);
  nand (_06960_, _06958_, _06706_);
  nand (_06962_, _06960_, _06959_);
  nand (_06963_, _06962_, _05489_);
  nor (_06964_, _06734_, _05812_);
  and (_06966_, _06964_, _06726_);
  and (_06967_, _06966_, _05517_);
  nor (_06968_, _06966_, _05517_);
  nor (_06969_, _06968_, _06967_);
  nor (_06970_, _06969_, _05882_);
  and (_06971_, _06487_, ABINPUT000[16]);
  nor (_06972_, _05517_, _05187_);
  nor (_06973_, _06972_, _05738_);
  nor (_06974_, _06973_, _05321_);
  nor (_06975_, _05210_, _05763_);
  nor (_06976_, _05517_, _05159_);
  and (_06977_, _06485_, ABINPUT000000[16]);
  or (_06978_, _06977_, _06976_);
  or (_06979_, _06978_, _06975_);
  or (_06980_, _06979_, _06974_);
  nor (_06981_, _06980_, _06971_);
  not (_06982_, _06981_);
  nor (_06983_, _06982_, _06970_);
  nand (_06984_, _06983_, _06963_);
  and (_06985_, _06984_, _06613_);
  and (_06986_, _06628_, _05867_);
  nor (_06987_, _06986_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_06988_, _06987_);
  and (_06989_, _06988_, _06638_);
  not (_06990_, _06989_);
  and (_06991_, _06986_, _05872_);
  nor (_06992_, _06991_, _06990_);
  not (_06993_, _05654_);
  and (_06994_, _05716_, _06993_);
  nor (_06996_, _05716_, _06993_);
  nor (_06997_, _06996_, _06994_);
  and (_06998_, _06997_, _05650_);
  not (_06999_, _06998_);
  nor (_07000_, _06993_, _05646_);
  and (_07001_, _06993_, _05646_);
  nor (_07002_, _07001_, _07000_);
  and (_07003_, _07002_, _05489_);
  and (_07004_, _05280_, _05766_);
  and (_07005_, _06487_, ABINPUT000[8]);
  or (_07006_, _07005_, _07004_);
  nor (_07007_, _05627_, _05174_);
  nor (_07008_, _05510_, _05159_);
  and (_07009_, _05187_, _05744_);
  and (_07010_, _06485_, ABINPUT000000[8]);
  or (_07011_, _07010_, _07009_);
  or (_07012_, _07011_, _07008_);
  nor (_07013_, _07012_, _07007_);
  nand (_07014_, _07013_, _05894_);
  or (_07015_, _07014_, _07006_);
  nor (_07016_, _06531_, _05732_);
  and (_07017_, _07016_, _05510_);
  nor (_07018_, _07016_, _05510_);
  nor (_07019_, _07018_, _07017_);
  nor (_07020_, _07019_, _05737_);
  not (_07021_, _07020_);
  nand (_07023_, _07021_, _05891_);
  or (_07024_, _07023_, _07015_);
  nor (_07025_, _07024_, _05898_);
  not (_07026_, _07025_);
  nor (_07027_, _07026_, _07003_);
  and (_07028_, _07027_, _06999_);
  nor (_07029_, _07028_, _06622_);
  or (_07030_, _07029_, _06992_);
  and (_07031_, _07030_, _06637_);
  or (_07032_, _07031_, _06985_);
  and (_05360_, _07032_, _05110_);
  and (_07033_, _06177_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_07034_, _06798_, _05995_);
  and (_07035_, _07034_, _06165_);
  or (_07037_, _07035_, _07033_);
  and (_05428_, _07037_, _05110_);
  and (_07038_, _06813_, _06342_);
  and (_07039_, _07038_, _06431_);
  and (_07040_, _06460_, _06276_);
  and (_07041_, _07040_, _06437_);
  or (_07043_, _07041_, _07039_);
  and (_07044_, _07038_, _06460_);
  and (_07045_, _06452_, _06431_);
  or (_07046_, _07045_, _07044_);
  and (_07048_, _07038_, _06464_);
  or (_07049_, _07048_, _07046_);
  or (_07050_, _07049_, _07043_);
  and (_07051_, _06810_, _06452_);
  or (_07052_, _07051_, _06837_);
  or (_07053_, _07052_, _06442_);
  or (_07054_, _07053_, _07050_);
  and (_07055_, _07054_, _06842_);
  nor (_07056_, _06870_, _06440_);
  and (_07057_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_07058_, _07057_, _07056_);
  and (_07059_, _07058_, _05110_);
  or (_05430_, _07059_, _07055_);
  and (_07060_, _06807_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_07061_, _07040_, _06459_);
  nor (_07062_, _06431_, _06276_);
  and (_07063_, _07062_, _06826_);
  and (_07064_, _07063_, _06459_);
  or (_07065_, _07064_, _07061_);
  not (_07066_, _06460_);
  not (_07067_, _06298_);
  and (_07068_, _06851_, _07067_);
  and (_07069_, _07068_, _06277_);
  and (_07070_, _06319_, _07067_);
  and (_07071_, _07070_, _06436_);
  and (_07072_, _07071_, _06277_);
  nor (_07073_, _07072_, _07069_);
  nor (_07074_, _07073_, _07066_);
  or (_07075_, _07074_, _07065_);
  and (_07076_, _07069_, _06447_);
  and (_07077_, _06451_, _06343_);
  and (_07078_, _07069_, _06464_);
  and (_07079_, _06456_, _07067_);
  and (_07080_, _07079_, _06277_);
  and (_07081_, _07080_, _06810_);
  or (_07082_, _07081_, _07078_);
  or (_07083_, _07082_, _07077_);
  or (_07084_, _07083_, _07076_);
  or (_07085_, _07084_, _07075_);
  and (_07086_, _07080_, _06447_);
  and (_07087_, _07068_, _06276_);
  and (_07088_, _07087_, _06864_);
  and (_07089_, _07080_, _06434_);
  or (_07090_, _07089_, _07088_);
  or (_07091_, _07090_, _07086_);
  not (_07092_, _06834_);
  and (_07093_, _06813_, _06448_);
  or (_07094_, _07093_, _07092_);
  and (_07095_, _07068_, _06455_);
  or (_07096_, _07095_, _06457_);
  or (_07097_, _06823_, _06465_);
  or (_07098_, _07097_, _07096_);
  or (_07099_, _07098_, _07094_);
  or (_07100_, _07099_, _06822_);
  or (_07101_, _07100_, _07091_);
  or (_07103_, _07101_, _07085_);
  and (_07104_, _07103_, _06842_);
  or (_05477_, _07104_, _07060_);
  and (_07105_, _06864_, _06814_);
  and (_07106_, _07105_, _06276_);
  and (_07107_, _06810_, _06276_);
  and (_07108_, _07107_, _06851_);
  or (_07109_, _06811_, _06452_);
  nand (_07110_, _07109_, _06864_);
  not (_07111_, _07110_);
  or (_07113_, _07111_, _07108_);
  or (_07114_, _07113_, _07106_);
  and (_07115_, _06831_, _06810_);
  and (_07116_, _06459_, _06451_);
  or (_07117_, _07116_, _06845_);
  or (_07118_, _07117_, _07115_);
  or (_07119_, _07118_, _07086_);
  and (_07120_, _06864_, _06463_);
  and (_07121_, _06941_, _06276_);
  or (_07122_, _07121_, _07120_);
  or (_07123_, _07122_, _07076_);
  or (_07124_, _07123_, _07119_);
  or (_07125_, _07124_, _07114_);
  and (_07126_, _06851_, _06830_);
  and (_07127_, _06455_, _06343_);
  or (_07128_, _07127_, _07126_);
  nor (_07129_, _07128_, _06462_);
  nand (_07130_, _07129_, _06834_);
  and (_07131_, _06851_, _07040_);
  and (_07132_, _07063_, _06343_);
  or (_07133_, _07132_, _06823_);
  or (_07134_, _07133_, _07131_);
  and (_07135_, _06455_, _06437_);
  or (_07136_, _07135_, _06867_);
  and (_07137_, _06460_, _06438_);
  and (_07138_, _07079_, _06276_);
  and (_07139_, _07138_, _06447_);
  or (_07140_, _07139_, _07137_);
  or (_07141_, _07140_, _07136_);
  or (_07142_, _07141_, _07134_);
  or (_07143_, _07142_, _07130_);
  or (_07144_, _07143_, _07125_);
  and (_07145_, _07144_, _05474_);
  and (_07146_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_07147_, _06820_, _06451_);
  and (_07148_, _07147_, _06873_);
  or (_07149_, _06874_, _06443_);
  or (_07150_, _07149_, _07148_);
  or (_07151_, _07150_, _07146_);
  or (_07152_, _07151_, _07145_);
  and (_05513_, _07152_, _05110_);
  not (_07153_, _05473_);
  or (_07154_, _06362_, _07153_);
  or (_07155_, _05473_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_07156_, _07155_, _05110_);
  and (_05525_, _07156_, _07154_);
  nor (_05565_, _06294_, rst);
  nor (_07157_, _05474_, _05492_);
  and (_07158_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_07159_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_07160_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_07161_, _07160_, _07159_);
  and (_07162_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_07163_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_07164_, _07163_, _07162_);
  and (_07165_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  not (_07167_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_07168_, _06251_, _07167_);
  nor (_07169_, _07168_, _07165_);
  and (_07170_, _07169_, _07164_);
  and (_07171_, _07170_, _07161_);
  nor (_07172_, _07171_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07173_, _07172_, _07158_);
  nor (_07174_, _07173_, _06200_);
  nor (_07176_, _07174_, _07157_);
  nor (_05569_, _07176_, rst);
  not (_07177_, _06471_);
  or (_07178_, _06699_, _06693_);
  nand (_07179_, _06699_, _06693_);
  and (_07180_, _07179_, _05489_);
  nand (_07181_, _07180_, _07178_);
  and (_07182_, _06588_, _05526_);
  and (_07183_, _06593_, _05703_);
  nor (_07184_, _07183_, _07182_);
  and (_07185_, _07184_, _05306_);
  nor (_07186_, _07184_, _05306_);
  nor (_07187_, _07186_, _07185_);
  and (_07188_, _07187_, _05291_);
  and (_07190_, _06487_, ABINPUT000[13]);
  nor (_07191_, _05306_, _05187_);
  nor (_07192_, _05188_, _05150_);
  or (_07193_, _07192_, _07191_);
  and (_07194_, _07193_, _05320_);
  and (_07195_, _05280_, _05762_);
  nor (_07196_, _05306_, _05159_);
  and (_07197_, _06485_, ABINPUT000000[13]);
  or (_07198_, _07197_, _07196_);
  or (_07199_, _07198_, _07195_);
  or (_07200_, _07199_, _07194_);
  nor (_07201_, _07200_, _07190_);
  not (_07202_, _07201_);
  nor (_07203_, _07202_, _07188_);
  nand (_07204_, _07203_, _07181_);
  or (_07205_, _07204_, _07177_);
  and (_07206_, _06146_, _05804_);
  and (_07207_, _07206_, _06631_);
  not (_07208_, _07207_);
  nor (_07209_, _05711_, _05309_);
  and (_07210_, _05711_, _05309_);
  nor (_07211_, _07210_, _07209_);
  and (_07212_, _07211_, _05650_);
  not (_07213_, _07212_);
  nor (_07214_, _05575_, _05309_);
  nor (_07215_, _07214_, _05490_);
  and (_07216_, _07215_, _05576_);
  nor (_07217_, _06649_, _05158_);
  nor (_07218_, _07217_, _05150_);
  not (_07219_, _07218_);
  and (_07220_, _05729_, _05150_);
  or (_07221_, _05597_, _05169_);
  nor (_07222_, _05210_, _05174_);
  and (_07223_, _06485_, ABINPUT000000[5]);
  and (_07224_, _06487_, ABINPUT000[5]);
  nor (_07225_, _07224_, _07223_);
  not (_07226_, _07225_);
  nor (_07227_, _07226_, _07222_);
  and (_07228_, _07227_, _07221_);
  not (_07229_, _07228_);
  nor (_07230_, _07229_, _07220_);
  and (_07231_, _07230_, _07219_);
  and (_07232_, _07231_, _05333_);
  not (_07233_, _07232_);
  nor (_07234_, _07233_, _07216_);
  and (_07235_, _07234_, _07213_);
  nor (_07236_, _07235_, _07208_);
  and (_07237_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_07238_, _07237_, _06471_);
  or (_07239_, _07238_, _07236_);
  and (_07240_, _07239_, _05110_);
  and (_05657_, _07240_, _07205_);
  or (_07241_, _06610_, _07177_);
  nand (_07242_, _07207_, _06668_);
  or (_07243_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_07244_, _07243_, _07242_);
  or (_07245_, _07244_, _06471_);
  and (_07246_, _07245_, _05110_);
  and (_05660_, _07246_, _07241_);
  or (_07247_, _06745_, _07177_);
  nor (_07248_, _07208_, _06780_);
  and (_07250_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_07251_, _07250_, _06471_);
  or (_07252_, _07251_, _07248_);
  and (_07253_, _07252_, _05110_);
  and (_05665_, _07253_, _07247_);
  not (_07254_, _06696_);
  nand (_07255_, _07179_, _07254_);
  nor (_07256_, _06701_, _05490_);
  nand (_07257_, _07256_, _07255_);
  and (_07258_, _06722_, _05603_);
  not (_07259_, _07258_);
  nor (_07260_, _06722_, _05603_);
  nor (_07261_, _07260_, _05882_);
  and (_07262_, _07261_, _07259_);
  and (_07263_, _05281_, _05762_);
  and (_07264_, _06487_, ABINPUT000[14]);
  nor (_07265_, _07264_, _07263_);
  and (_07266_, _05597_, _05187_);
  not (_07267_, _07266_);
  nor (_07268_, _06723_, _05321_);
  and (_07269_, _07268_, _07267_);
  nor (_07270_, _05603_, _05159_);
  and (_07271_, _06485_, ABINPUT000000[14]);
  or (_07272_, _07271_, _07270_);
  nor (_07273_, _07272_, _07269_);
  and (_07274_, _07273_, _07265_);
  not (_07275_, _07274_);
  nor (_07276_, _07275_, _07262_);
  nand (_07277_, _07276_, _07257_);
  or (_07278_, _07277_, _07177_);
  nor (_07279_, _07208_, _06548_);
  and (_07280_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_07281_, _07280_, _06471_);
  or (_07282_, _07281_, _07279_);
  and (_07283_, _07282_, _05110_);
  and (_05670_, _07283_, _07278_);
  or (_07284_, _06575_, _06572_);
  nor (_07285_, _06576_, _05490_);
  nand (_07286_, _07285_, _07284_);
  nor (_07287_, _06586_, _05188_);
  nor (_07288_, _06591_, _05187_);
  nor (_07289_, _07288_, _07287_);
  and (_07290_, _07289_, _05534_);
  nor (_07291_, _07289_, _05534_);
  nor (_07292_, _07291_, _07290_);
  nor (_07293_, _07292_, _05882_);
  nor (_07294_, _05627_, _05763_);
  nor (_07295_, _05534_, _05159_);
  and (_07296_, _06485_, ABINPUT000000[11]);
  or (_07297_, _07296_, _07295_);
  nor (_07298_, _07297_, _07294_);
  nor (_07299_, _05321_, _05233_);
  and (_07300_, _06487_, ABINPUT000[11]);
  nor (_07301_, _07300_, _07299_);
  and (_07302_, _07301_, _07298_);
  not (_07303_, _07302_);
  nor (_07304_, _07303_, _07293_);
  nand (_07305_, _07304_, _07286_);
  or (_07306_, _07305_, _07177_);
  or (_07307_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_07308_, _05699_, _05692_);
  nor (_07309_, _07308_, _05700_);
  nor (_07310_, _07309_, _05651_);
  and (_07311_, _05726_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_07312_, _06500_, _05233_);
  nor (_07313_, _07312_, _07311_);
  nor (_07314_, _07313_, _05737_);
  not (_07315_, _06226_);
  nor (_07316_, _05233_, _05159_);
  and (_07317_, _06487_, ABINPUT000[3]);
  nor (_07318_, _07317_, _07316_);
  or (_07319_, _05210_, _05169_);
  and (_07320_, _05281_, _05172_);
  and (_07321_, _06485_, ABINPUT000000[3]);
  nor (_07322_, _07321_, _07320_);
  and (_07323_, _07322_, _07319_);
  and (_07324_, _07323_, _07318_);
  and (_07325_, _07324_, _07315_);
  not (_07326_, _07325_);
  nor (_07327_, _07326_, _07314_);
  not (_07328_, _07327_);
  nor (_07329_, _07328_, _07310_);
  nor (_07330_, _05568_, _05566_);
  not (_07331_, _07330_);
  nor (_07332_, _05570_, _05490_);
  and (_07333_, _07332_, _07331_);
  and (_07334_, _06222_, _06219_);
  not (_07335_, _07334_);
  nor (_07336_, _07335_, _07333_);
  and (_07337_, _07336_, _07329_);
  nand (_07338_, _07337_, _07207_);
  and (_07339_, _07338_, _07307_);
  or (_07340_, _07339_, _06471_);
  and (_07341_, _07340_, _05110_);
  and (_05680_, _07341_, _07306_);
  or (_07342_, _06571_, _06568_);
  nor (_07343_, _06572_, _05490_);
  nand (_07344_, _07343_, _07342_);
  nor (_07345_, _06711_, _05187_);
  nor (_07346_, _06585_, _05188_);
  or (_07347_, _07346_, _07345_);
  nor (_07348_, _07347_, _05543_);
  and (_07349_, _07347_, _05543_);
  nor (_07350_, _07349_, _07348_);
  nor (_07351_, _07350_, _05882_);
  nor (_07352_, _05597_, _05763_);
  and (_07353_, _05543_, _05158_);
  and (_07354_, _06485_, ABINPUT000000[10]);
  or (_07355_, _07354_, _07353_);
  nor (_07356_, _07355_, _07352_);
  and (_07358_, _05320_, _05281_);
  and (_07359_, _06487_, ABINPUT000[10]);
  nor (_07360_, _07359_, _07358_);
  and (_07361_, _07360_, _07356_);
  not (_07362_, _07361_);
  nor (_07363_, _07362_, _07351_);
  nand (_07364_, _07363_, _07344_);
  or (_07365_, _07364_, _07177_);
  or (_07366_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand (_07367_, _07207_, _06512_);
  and (_07368_, _07367_, _07366_);
  or (_07369_, _07368_, _06471_);
  and (_07370_, _07369_, _05110_);
  and (_05688_, _07370_, _07365_);
  or (_07371_, _06567_, _06564_);
  nor (_07372_, _06568_, _05490_);
  nand (_07373_, _07372_, _07371_);
  nor (_07374_, _06584_, _05876_);
  nor (_07375_, _07374_, _05886_);
  nor (_07376_, _07375_, _05550_);
  and (_07377_, _07375_, _05550_);
  nor (_07378_, _07377_, _07376_);
  and (_07379_, _07378_, _05291_);
  nor (_07380_, _05763_, _05150_);
  nor (_07381_, _05549_, _05159_);
  and (_07382_, _06485_, ABINPUT000000[9]);
  or (_07383_, _07382_, _07381_);
  nor (_07384_, _07383_, _07380_);
  and (_07385_, _05320_, _05280_);
  and (_07386_, _06487_, ABINPUT000[9]);
  nor (_07387_, _07386_, _07385_);
  and (_07388_, _07387_, _07384_);
  not (_07389_, _07388_);
  nor (_07390_, _07389_, _07379_);
  nand (_07391_, _07390_, _07373_);
  or (_07392_, _07391_, _07177_);
  or (_07393_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nor (_07394_, _05563_, _05187_);
  nor (_07395_, _07394_, _05564_);
  not (_07396_, _07395_);
  nor (_07397_, _05489_, _05650_);
  nor (_07398_, _07397_, _07396_);
  not (_07399_, _07398_);
  and (_07400_, _06709_, _05749_);
  not (_07401_, _07400_);
  and (_07402_, _06794_, _07401_);
  or (_07403_, _05274_, _05169_);
  nor (_07404_, _05725_, _05158_);
  nor (_07405_, _07404_, _05253_);
  not (_07406_, _07405_);
  and (_07407_, _07406_, _07403_);
  and (_07408_, _05187_, _05762_);
  and (_07409_, _06485_, ABINPUT000000[1]);
  and (_07410_, _06487_, ABINPUT000[1]);
  nor (_07411_, _07410_, _07409_);
  not (_07412_, _07411_);
  nor (_07413_, _07412_, _07408_);
  and (_07414_, _07413_, _07407_);
  and (_07415_, _07414_, _06791_);
  and (_07416_, _07415_, _07402_);
  and (_07417_, _07416_, _06788_);
  and (_07418_, _07417_, _07399_);
  nand (_07419_, _07418_, _07207_);
  and (_07420_, _07419_, _07393_);
  or (_07421_, _07420_, _06471_);
  and (_07422_, _07421_, _05110_);
  and (_05691_, _07422_, _07392_);
  and (_05695_, _06362_, _05110_);
  and (_05698_, _06384_, _05110_);
  and (_05701_, _06406_, _05110_);
  nor (_05704_, _06427_, rst);
  and (_05706_, _06271_, _05110_);
  nor (_05709_, _06338_, rst);
  nor (_05712_, _06315_, rst);
  nor (_07423_, _05474_, _05258_);
  and (_07424_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  not (_07425_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_07426_, _06251_, _07425_);
  nor (_07427_, _07426_, _07424_);
  and (_07428_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_07429_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_07430_, _07429_, _07428_);
  and (_07431_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_07432_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_07433_, _07432_, _07431_);
  and (_07434_, _07433_, _07430_);
  and (_07435_, _07434_, _07427_);
  and (_07436_, _05474_, _06254_);
  not (_07437_, _07436_);
  nor (_07438_, _07437_, _07435_);
  nor (_07439_, _07438_, _07423_);
  nor (_05721_, _07439_, rst);
  nor (_07440_, _05474_, _05212_);
  and (_07441_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  not (_07442_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_07443_, _06251_, _07442_);
  nor (_07444_, _07443_, _07441_);
  and (_07445_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_07446_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_07447_, _07446_, _07445_);
  and (_07448_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_07449_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_07450_, _07449_, _07448_);
  and (_07451_, _07450_, _07447_);
  and (_07452_, _07451_, _07444_);
  nor (_07453_, _07452_, _07437_);
  nor (_07454_, _07453_, _07440_);
  nor (_05724_, _07454_, rst);
  nor (_07455_, _05474_, _05189_);
  and (_07456_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  not (_07457_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_07458_, _06251_, _07457_);
  nor (_07459_, _07458_, _07456_);
  and (_07460_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_07461_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_07462_, _07461_, _07460_);
  and (_07463_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_07464_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_07465_, _07464_, _07463_);
  and (_07466_, _07465_, _07462_);
  and (_07467_, _07466_, _07459_);
  nor (_07469_, _07467_, _07437_);
  nor (_07470_, _07469_, _07455_);
  nor (_05727_, _07470_, rst);
  nor (_07471_, _05474_, _05111_);
  and (_07473_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  not (_07474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_07475_, _06251_, _07474_);
  nor (_07477_, _07475_, _07473_);
  and (_07478_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_07479_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_07480_, _07479_, _07478_);
  and (_07482_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_07483_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_07485_, _07483_, _07482_);
  and (_07486_, _07485_, _07480_);
  and (_07487_, _07486_, _07477_);
  nor (_07489_, _07487_, _07437_);
  nor (_07490_, _07489_, _07471_);
  nor (_05730_, _07490_, rst);
  nor (_07492_, _05474_, _05425_);
  and (_07493_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not (_07494_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_07496_, _06251_, _07494_);
  nor (_07497_, _07496_, _07493_);
  and (_07498_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_07499_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_07500_, _07499_, _07498_);
  and (_07501_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_07502_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_07503_, _07502_, _07501_);
  and (_07504_, _07503_, _07500_);
  and (_07505_, _07504_, _07497_);
  nor (_07506_, _07505_, _07437_);
  nor (_07507_, _07506_, _07492_);
  nor (_05733_, _07507_, rst);
  nor (_07508_, _05474_, _05260_);
  and (_07509_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_07510_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_07511_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_07512_, _07511_, _07510_);
  and (_07513_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  not (_07514_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_07515_, _06251_, _07514_);
  nor (_07516_, _07515_, _07513_);
  and (_07517_, _07516_, _07512_);
  and (_07518_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_07519_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_07520_, _07519_, _07518_);
  and (_07521_, _07520_, _07517_);
  nor (_07522_, _07521_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07523_, _07522_, _07509_);
  nor (_07524_, _07523_, _06200_);
  nor (_07525_, _07524_, _07508_);
  nor (_05745_, _07525_, rst);
  nor (_07526_, _05474_, _05214_);
  and (_07527_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_07528_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_07529_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_07530_, _07529_, _07528_);
  and (_07531_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not (_07532_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_07533_, _06251_, _07532_);
  nor (_07534_, _07533_, _07531_);
  and (_07535_, _07534_, _07530_);
  and (_07536_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_07537_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_07538_, _07537_, _07536_);
  and (_07539_, _07538_, _07535_);
  nor (_07540_, _07539_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07541_, _07540_, _07527_);
  nor (_07542_, _07541_, _06200_);
  nor (_07543_, _07542_, _07526_);
  nor (_05748_, _07543_, rst);
  nor (_07544_, _05474_, _05191_);
  and (_07545_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_07546_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_07547_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_07548_, _07547_, _07546_);
  and (_07549_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_07550_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_07551_, _07550_, _07549_);
  and (_07552_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not (_07553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_07554_, _06251_, _07553_);
  nor (_07555_, _07554_, _07552_);
  and (_07556_, _07555_, _07551_);
  and (_07557_, _07556_, _07548_);
  nor (_07558_, _07557_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07559_, _07558_, _07545_);
  nor (_07560_, _07559_, _06200_);
  nor (_07561_, _07560_, _07544_);
  nor (_05750_, _07561_, rst);
  nor (_07562_, _05474_, _05610_);
  and (_07563_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_07564_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_07565_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_07566_, _07565_, _07564_);
  and (_07567_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_07568_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_07569_, _07568_, _07567_);
  and (_07570_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  not (_07571_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_07572_, _06251_, _07571_);
  nor (_07574_, _07572_, _07570_);
  and (_07575_, _07574_, _07569_);
  and (_07576_, _07575_, _07566_);
  nor (_07578_, _07576_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07579_, _07578_, _07563_);
  nor (_07580_, _07579_, _06200_);
  nor (_07582_, _07580_, _07562_);
  nor (_05757_, _07582_, rst);
  nand (_07583_, _07235_, _06477_);
  or (_07585_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_07586_, _07585_, _05110_);
  and (_05772_, _07586_, _07583_);
  nor (_07588_, _07418_, _06476_);
  and (_07589_, _06476_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_07591_, _07589_, _07588_);
  and (_05775_, _07591_, _05110_);
  nand (_07592_, _06668_, _06477_);
  or (_07594_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_07595_, _07594_, _05110_);
  and (_05780_, _07595_, _07592_);
  nand (_07596_, _06780_, _06477_);
  or (_07598_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_07599_, _07598_, _05110_);
  and (_05783_, _07599_, _07596_);
  nor (_07600_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not (_07601_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07602_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _07601_);
  nor (_07603_, _07602_, _07600_);
  not (_07604_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_07605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_07606_, _06205_, _07605_);
  and (_07607_, _07606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_07608_, _07606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_07609_, _07608_, _07607_);
  nor (_07610_, _07609_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07611_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _07601_);
  nor (_07612_, _07611_, _07610_);
  nor (_07613_, _07612_, _07604_);
  and (_07614_, _07612_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_07615_, _07614_, _07613_);
  nor (_07616_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_07617_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _07601_);
  nor (_07618_, _07617_, _07616_);
  and (_07619_, _06205_, _07605_);
  nor (_07620_, _07619_, _07606_);
  nor (_07621_, _07620_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_07622_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _07601_);
  nor (_07623_, _07622_, _07621_);
  nor (_07624_, _07623_, _07618_);
  not (_07625_, _07624_);
  nor (_07626_, _07625_, _07615_);
  not (_07627_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_07628_, _07612_, _07627_);
  nor (_07629_, _07612_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_07630_, _07629_, _07628_);
  not (_07631_, _07630_);
  not (_07632_, _07618_);
  and (_07633_, _07623_, _07632_);
  and (_07634_, _07633_, _07631_);
  nor (_07635_, _07634_, _07626_);
  nor (_07636_, _07623_, _07632_);
  not (_07637_, _07636_);
  not (_07638_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_07640_, _07612_, _07638_);
  and (_07641_, _07612_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_07642_, _07641_, _07640_);
  nor (_07643_, _07642_, _07637_);
  and (_07644_, _07623_, _07618_);
  not (_07645_, _07644_);
  nor (_07646_, _07612_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_07647_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_07649_, _07612_, _07647_);
  or (_07650_, _07649_, _07646_);
  nor (_07651_, _07650_, _07645_);
  nor (_07652_, _07651_, _07643_);
  and (_07654_, _07652_, _07635_);
  and (_07656_, _07654_, _07603_);
  and (_07657_, _07612_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_07658_, _07657_, _07636_);
  not (_07659_, _07612_);
  and (_07660_, _07659_, _07636_);
  and (_07661_, _07660_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_07662_, _07661_, _07603_);
  or (_07663_, _07662_, _07658_);
  and (_07664_, _07612_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not (_07666_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_07667_, _07612_, _07666_);
  nor (_07668_, _07667_, _07664_);
  nor (_07669_, _07668_, _07625_);
  and (_07670_, _07659_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_07671_, _07612_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_07672_, _07671_, _07670_);
  nor (_07673_, _07672_, _07645_);
  not (_07674_, _07633_);
  not (_07675_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_07676_, _07612_, _07675_);
  nor (_07677_, _07612_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_07678_, _07677_, _07676_);
  nor (_07679_, _07678_, _07674_);
  or (_07680_, _07679_, _07673_);
  or (_07681_, _07680_, _07669_);
  nor (_07682_, _07681_, _07663_);
  nor (_07683_, _07682_, _07656_);
  not (_07684_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_07685_, _07603_, _07684_);
  or (_07687_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_07688_, _07687_, _07685_);
  and (_07690_, _07688_, _07644_);
  not (_07691_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_07693_, _07603_, _07691_);
  or (_07694_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_07695_, _07694_, _07693_);
  and (_07696_, _07695_, _07636_);
  or (_07698_, _07696_, _07690_);
  not (_07699_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_07701_, _07603_, _07699_);
  or (_07702_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_07704_, _07702_, _07701_);
  and (_07705_, _07704_, _07633_);
  not (_07706_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_07707_, _07603_, _07706_);
  or (_07709_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_07710_, _07709_, _07707_);
  and (_07711_, _07710_, _07624_);
  or (_07712_, _07711_, _07705_);
  or (_07714_, _07712_, _07698_);
  and (_07715_, _07714_, _07612_);
  not (_07716_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_07717_, _07603_, _07716_);
  or (_07718_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_07719_, _07718_, _07717_);
  and (_07720_, _07719_, _07636_);
  not (_07721_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_07722_, _07603_, _07721_);
  or (_07723_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_07724_, _07723_, _07722_);
  and (_07725_, _07724_, _07644_);
  or (_07726_, _07725_, _07720_);
  not (_07727_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_07728_, _07603_, _07727_);
  or (_07729_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_07730_, _07729_, _07728_);
  and (_07731_, _07730_, _07633_);
  not (_07732_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_07733_, _07603_, _07732_);
  or (_07734_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_07735_, _07734_, _07733_);
  and (_07736_, _07735_, _07624_);
  or (_07737_, _07736_, _07731_);
  or (_07738_, _07737_, _07726_);
  and (_07739_, _07738_, _07659_);
  or (_07740_, _07739_, _07715_);
  and (_07741_, _07740_, _07683_);
  not (_07742_, _07683_);
  and (_07743_, _07742_, word_in[7]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07743_, _07741_);
  and (_07744_, _07632_, _07603_);
  not (_07745_, _07744_);
  and (_07746_, _07618_, _07603_);
  nor (_07747_, _07746_, _07623_);
  and (_07748_, _07746_, _07623_);
  nor (_07749_, _07748_, _07747_);
  not (_07750_, _07749_);
  nor (_07751_, _07750_, _07672_);
  nor (_07752_, _07748_, _07659_);
  not (_07753_, _07623_);
  nor (_07754_, _07612_, _07753_);
  and (_07755_, _07746_, _07754_);
  nor (_07756_, _07755_, _07752_);
  nor (_07757_, _07756_, _07749_);
  and (_07759_, _07757_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_07760_, _07756_, _07750_);
  and (_07761_, _07760_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_07762_, _07761_, _07759_);
  nor (_07763_, _07762_, _07751_);
  nor (_07764_, _07763_, _07745_);
  not (_07765_, _07764_);
  not (_07766_, _07746_);
  nor (_07767_, _07750_, _07678_);
  and (_07768_, _07760_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_07769_, _07768_, _07767_);
  or (_07770_, _07769_, _07766_);
  nand (_07771_, _07755_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_07772_, _07771_, _07770_);
  and (_07773_, _07772_, _07765_);
  not (_07774_, _07603_);
  and (_07775_, _07618_, _07774_);
  not (_07776_, _07775_);
  nor (_07777_, _07750_, _07650_);
  and (_07778_, _07757_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_07779_, _07760_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_07780_, _07779_, _07778_);
  nor (_07781_, _07780_, _07777_);
  nor (_07782_, _07781_, _07776_);
  nor (_07783_, _07618_, _07603_);
  not (_07784_, _07783_);
  nor (_07785_, _07750_, _07630_);
  and (_07786_, _07757_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_07787_, _07760_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_07788_, _07787_, _07786_);
  nor (_07789_, _07788_, _07785_);
  nor (_07790_, _07789_, _07784_);
  nor (_07791_, _07790_, _07782_);
  and (_07793_, _07791_, _07773_);
  or (_07794_, _07746_, _07783_);
  not (_07796_, _07794_);
  not (_07797_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_07799_, _07603_, _07797_);
  or (_07800_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_07801_, _07800_, _07799_);
  and (_07802_, _07801_, _07796_);
  not (_07804_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_07805_, _07603_, _07804_);
  or (_07806_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_07808_, _07806_, _07805_);
  and (_07809_, _07808_, _07794_);
  or (_07810_, _07809_, _07802_);
  and (_07811_, _07810_, _07757_);
  and (_07813_, _07749_, _07612_);
  not (_07814_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_07815_, _07603_, _07814_);
  or (_07816_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_07818_, _07816_, _07815_);
  and (_07819_, _07818_, _07796_);
  not (_07820_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_07821_, _07603_, _07820_);
  or (_07823_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_07824_, _07823_, _07821_);
  and (_07825_, _07824_, _07794_);
  or (_07826_, _07825_, _07819_);
  and (_07827_, _07826_, _07813_);
  or (_07828_, _07827_, _07811_);
  not (_07829_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_07830_, _07603_, _07829_);
  or (_07831_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_07832_, _07831_, _07830_);
  and (_07833_, _07832_, _07794_);
  not (_07834_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_07835_, _07603_, _07834_);
  or (_07836_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_07837_, _07836_, _07835_);
  and (_07838_, _07837_, _07796_);
  or (_07839_, _07838_, _07833_);
  and (_07840_, _07839_, _07760_);
  and (_07841_, _07749_, _07659_);
  not (_07842_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_07843_, _07603_, _07842_);
  or (_07844_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_07845_, _07844_, _07843_);
  and (_07846_, _07845_, _07794_);
  not (_07847_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_07848_, _07603_, _07847_);
  or (_07849_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_07850_, _07849_, _07848_);
  and (_07851_, _07850_, _07796_);
  or (_07852_, _07851_, _07846_);
  and (_07853_, _07852_, _07841_);
  or (_07854_, _07853_, _07840_);
  nor (_07855_, _07854_, _07828_);
  nor (_07856_, _07855_, _07793_);
  and (_07857_, _07793_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07857_, _07856_);
  nor (_07858_, _07644_, _07624_);
  not (_07859_, _07858_);
  nor (_07860_, _07859_, _07630_);
  and (_07861_, _07644_, _07612_);
  nor (_07862_, _07644_, _07612_);
  nor (_07863_, _07862_, _07861_);
  and (_07865_, _07863_, _07859_);
  and (_07866_, _07865_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_07868_, _07863_, _07858_);
  and (_07869_, _07868_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_07870_, _07869_, _07866_);
  nor (_07871_, _07870_, _07860_);
  nor (_07872_, _07871_, _07766_);
  and (_07873_, _07868_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_07874_, _07873_);
  nor (_07875_, _07859_, _07650_);
  and (_07876_, _07865_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_07877_, _07876_, _07875_);
  and (_07879_, _07877_, _07874_);
  nor (_07880_, _07879_, _07745_);
  nor (_07881_, _07880_, _07872_);
  and (_07882_, _07868_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_07883_, _07882_);
  nor (_07884_, _07859_, _07672_);
  and (_07885_, _07865_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_07886_, _07885_, _07884_);
  and (_07887_, _07886_, _07883_);
  nor (_07888_, _07887_, _07784_);
  nor (_07889_, _07859_, _07678_);
  and (_07890_, _07865_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_07891_, _07868_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_07892_, _07891_, _07890_);
  nor (_07893_, _07892_, _07889_);
  nor (_07894_, _07893_, _07776_);
  nor (_07895_, _07894_, _07888_);
  and (_07896_, _07895_, _07881_);
  and (_07897_, _07896_, word_in[23]);
  and (_07898_, _07730_, _07636_);
  and (_07899_, _07719_, _07624_);
  or (_07901_, _07899_, _07898_);
  and (_07902_, _07724_, _07633_);
  and (_07903_, _07735_, _07644_);
  or (_07904_, _07903_, _07902_);
  or (_07905_, _07904_, _07901_);
  or (_07906_, _07905_, _07863_);
  not (_07907_, _07863_);
  and (_07908_, _07688_, _07633_);
  and (_07909_, _07710_, _07659_);
  or (_07910_, _07909_, _07908_);
  and (_07912_, _07704_, _07636_);
  and (_07913_, _07695_, _07624_);
  or (_07914_, _07913_, _07912_);
  or (_07916_, _07914_, _07910_);
  or (_07917_, _07916_, _07907_);
  nand (_07920_, _07917_, _07906_);
  nor (_07921_, _07920_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07921_, _07897_);
  and (_07923_, _07748_, _07612_);
  and (_07925_, _07923_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_07926_, _07784_, _07623_);
  not (_07927_, _07926_);
  nand (_07929_, _07784_, _07623_);
  and (_07930_, _07929_, _07927_);
  not (_07931_, _07930_);
  nor (_07933_, _07672_, _07931_);
  nor (_07935_, _07929_, _07612_);
  and (_07936_, _07929_, _07612_);
  nor (_07937_, _07936_, _07935_);
  nor (_07938_, _07937_, _07930_);
  and (_07939_, _07938_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_07940_, _07939_, _07933_);
  nor (_07941_, _07940_, _07766_);
  nor (_07942_, _07678_, _07931_);
  and (_07943_, _07938_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_07944_, _07937_, _07931_);
  and (_07945_, _07944_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_07946_, _07945_, _07943_);
  nor (_07947_, _07946_, _07942_);
  nor (_07948_, _07947_, _07745_);
  or (_07949_, _07948_, _07941_);
  nor (_07950_, _07949_, _07925_);
  and (_07951_, _07930_, _07631_);
  and (_07952_, _07944_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_07953_, _07938_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_07954_, _07953_, _07952_);
  nor (_07955_, _07954_, _07951_);
  nor (_07956_, _07955_, _07776_);
  nor (_07957_, _07931_, _07650_);
  and (_07958_, _07938_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_07959_, _07958_, _07957_);
  nor (_07960_, _07959_, _07784_);
  and (_07961_, _07926_, _07640_);
  or (_07962_, _07961_, _07960_);
  nor (_07963_, _07962_, _07956_);
  and (_07964_, _07963_, _07950_);
  and (_07965_, _07808_, _07796_);
  and (_07966_, _07801_, _07794_);
  or (_07967_, _07966_, _07965_);
  and (_07968_, _07967_, _07938_);
  and (_07969_, _07832_, _07796_);
  and (_07970_, _07837_, _07794_);
  or (_07971_, _07970_, _07969_);
  and (_07972_, _07971_, _07944_);
  and (_07973_, _07930_, _07659_);
  and (_07974_, _07845_, _07796_);
  and (_07975_, _07850_, _07794_);
  or (_07976_, _07975_, _07974_);
  and (_07977_, _07976_, _07973_);
  and (_07978_, _07824_, _07796_);
  and (_07979_, _07818_, _07794_);
  or (_07980_, _07979_, _07978_);
  and (_07981_, _07936_, _07927_);
  and (_07982_, _07981_, _07980_);
  or (_07983_, _07982_, _07977_);
  or (_07984_, _07983_, _07972_);
  nor (_07985_, _07984_, _07968_);
  nor (_07986_, _07985_, _07964_);
  and (_07987_, _07964_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _07987_, _07986_);
  and (_07988_, _07612_, _07623_);
  nor (_07989_, _07861_, _07647_);
  or (_07990_, _07989_, _07988_);
  and (_06013_, _07990_, _05110_);
  and (_07992_, _07858_, _07612_);
  and (_07993_, _07896_, _05110_);
  and (_07995_, _07993_, _07744_);
  and (_07996_, _07995_, _07992_);
  not (_07998_, _07996_);
  and (_07999_, _07793_, _05110_);
  and (_08001_, _07999_, _07775_);
  and (_08002_, _08001_, _07813_);
  and (_08004_, _07656_, _05110_);
  and (_08005_, _08004_, _07618_);
  nor (_08007_, _07683_, rst);
  and (_08008_, _08007_, _07988_);
  and (_08010_, _08008_, _08005_);
  and (_08011_, _08007_, word_in[7]);
  and (_08013_, _08011_, _08010_);
  nor (_08014_, _08010_, _07684_);
  nor (_08015_, _08014_, _08013_);
  nor (_08016_, _08015_, _08002_);
  and (_08017_, _08002_, word_in[15]);
  or (_08018_, _08017_, _08016_);
  and (_08019_, _08018_, _07998_);
  and (_08020_, _07988_, _07783_);
  and (_08021_, _07964_, _05110_);
  and (_08022_, _08021_, _08020_);
  and (_08023_, _07993_, word_in[23]);
  and (_08024_, _08023_, _07996_);
  or (_08025_, _08024_, _08022_);
  or (_08026_, _08025_, _08019_);
  not (_08027_, _08022_);
  and (_08028_, _08021_, word_in[31]);
  or (_08029_, _08028_, _08027_);
  and (_06039_, _08029_, _08026_);
  or (_08030_, _07944_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_06060_, _08030_, _05110_);
  and (_08031_, _07624_, _07659_);
  or (_08032_, _08031_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08033_, _08032_, _07861_);
  and (_06090_, _08033_, _05110_);
  nor (_08034_, _08031_, _07923_);
  or (_08035_, _07745_, _07623_);
  nor (_08036_, _08035_, _07612_);
  and (_08037_, _07775_, _07973_);
  nor (_08038_, _08037_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08039_, _08038_, _08036_);
  nand (_08040_, _08039_, _08034_);
  and (_06133_, _08040_, _05110_);
  not (_08041_, _07760_);
  and (_08042_, _07746_, _07973_);
  or (_08043_, _08042_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_08044_, _08043_, _08041_);
  and (_08045_, _07624_, _07640_);
  or (_08046_, _08045_, _08037_);
  or (_08047_, _08046_, _08044_);
  and (_08048_, _08047_, _08034_);
  and (_08049_, _08043_, _07923_);
  or (_08050_, _08049_, _08031_);
  or (_08051_, _08050_, _08048_);
  and (_06181_, _08051_, _05110_);
  not (_08052_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_08053_, _06001_, _05337_);
  nor (_08054_, _08053_, _08052_);
  not (_08056_, _08053_);
  nor (_08057_, _08056_, _06088_);
  or (_08058_, _08057_, _08054_);
  and (_06192_, _08058_, _05110_);
  and (_08059_, _07754_, _07783_);
  or (_08060_, _08059_, _08042_);
  or (_08061_, _08060_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_08062_, _08061_, _08041_);
  and (_08063_, _07926_, _07659_);
  or (_08064_, _08063_, _07923_);
  and (_08065_, _08064_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08066_, _08065_, _08036_);
  or (_08067_, _08066_, _08062_);
  or (_08068_, _08067_, _08037_);
  and (_06236_, _08068_, _05110_);
  nor (_08069_, _08063_, _07973_);
  not (_08070_, _07862_);
  or (_08071_, _08070_, _08060_);
  and (_08072_, _08071_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08073_, _08037_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08074_, _07744_, _07754_);
  and (_08075_, _08031_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08076_, _08075_, _08074_);
  or (_08078_, _08076_, _08073_);
  or (_08079_, _08078_, _08072_);
  and (_08081_, _08079_, _08069_);
  and (_08082_, _08063_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08083_, _08036_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08085_, _08083_, _08037_);
  or (_08086_, _08085_, _08082_);
  or (_08087_, _08086_, _08059_);
  or (_08088_, _08087_, _08042_);
  or (_08090_, _08088_, _08081_);
  and (_06299_, _08090_, _05110_);
  or (_08092_, _07752_, _07935_);
  and (_08093_, _07644_, _07659_);
  or (_08095_, _07752_, _08093_);
  and (_08096_, _07775_, _07754_);
  or (_08097_, _08096_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08099_, _08097_, _08095_);
  and (_08100_, _08060_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08101_, _08100_, _08074_);
  or (_08102_, _08101_, _08099_);
  and (_08104_, _08102_, _08092_);
  and (_08105_, _08097_, _07923_);
  and (_08106_, _07670_, _07747_);
  or (_08107_, _08106_, _08042_);
  or (_08108_, _08107_, _08059_);
  or (_08109_, _08108_, _08105_);
  or (_08110_, _08109_, _08104_);
  and (_06361_, _08110_, _05110_);
  not (_08111_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_08112_, _08053_, _08111_);
  nor (_08113_, _08056_, _06229_);
  or (_08114_, _08113_, _08112_);
  and (_06372_, _08114_, _05110_);
  and (_08115_, _08053_, _06559_);
  not (_08116_, _06903_);
  or (_08117_, _08116_, _06555_);
  and (_08118_, _08117_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_08119_, _08118_, _08115_);
  and (_06408_, _08119_, _05110_);
  or (_08120_, _07748_, _07612_);
  or (_08121_, _07755_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08122_, _08121_, _08120_);
  and (_08123_, _07973_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08124_, _08063_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_08125_, _08124_, _08059_);
  or (_08126_, _08125_, _08123_);
  or (_08127_, _08126_, _08096_);
  or (_08128_, _08127_, _08074_);
  or (_08129_, _08128_, _08122_);
  and (_06441_, _08129_, _05110_);
  nor (_08130_, _06628_, _05591_);
  and (_08131_, _06625_, _05794_);
  and (_08132_, _08131_, _06626_);
  and (_08133_, _05912_, _05485_);
  and (_08134_, _08133_, _05782_);
  nor (_08135_, _08133_, _05591_);
  or (_08136_, _08135_, _08134_);
  nand (_08137_, _08136_, _08132_);
  nand (_08138_, _08137_, _06622_);
  or (_08139_, _08138_, _08130_);
  and (_08140_, _06623_, _06548_);
  nor (_08141_, _08140_, _06613_);
  nand (_08142_, _08141_, _08139_);
  nand (_08143_, _07277_, _06613_);
  nand (_08144_, _08143_, _08142_);
  and (_06474_, _08144_, _05110_);
  nor (_08145_, _07418_, _06622_);
  nor (_08146_, _08145_, _06613_);
  and (_08147_, _08132_, _05805_);
  nand (_08148_, _08147_, _05872_);
  nor (_08149_, _08147_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not (_08150_, _08149_);
  and (_08151_, _08150_, _06638_);
  nand (_08152_, _08151_, _08148_);
  nand (_08153_, _08152_, _08146_);
  or (_08154_, _07391_, _06637_);
  and (_08155_, _08154_, _08153_);
  and (_06484_, _08155_, _05110_);
  and (_08156_, _07926_, _07612_);
  or (_08157_, _08156_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08158_, _08157_, _07612_);
  or (_08159_, _08031_, _07660_);
  and (_08160_, _08159_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08161_, _08059_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08162_, _08074_, _07755_);
  or (_08163_, _08162_, _08161_);
  or (_08164_, _08163_, _08160_);
  or (_08165_, _08164_, _08096_);
  or (_08166_, _08165_, _08158_);
  and (_06527_, _08166_, _05110_);
  and (_08167_, _07752_, _07927_);
  nor (_08168_, _08035_, _07659_);
  or (_08169_, _08168_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08170_, _08169_, _08167_);
  or (_08172_, _08170_, _08156_);
  and (_08173_, _07862_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08174_, _08169_, _07923_);
  or (_08176_, _08174_, _08093_);
  or (_08177_, _08176_, _08173_);
  or (_08178_, _08177_, _08172_);
  and (_06614_, _08178_, _05110_);
  not (_08179_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_08180_, _08053_, _08179_);
  nor (_08181_, _08056_, _05334_);
  or (_08182_, _08181_, _08180_);
  and (_06684_, _08182_, _05110_);
  and (_08183_, _07752_, _07625_);
  or (_08184_, _08183_, _07923_);
  and (_08186_, _07796_, _07973_);
  and (_08187_, _08186_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08188_, _08156_, _07755_);
  and (_08189_, _08188_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08190_, _07775_, _07936_);
  and (_08191_, _08063_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08192_, _08191_, _08190_);
  and (_08193_, _07841_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_08194_, _08035_, _07747_);
  and (_08195_, _08194_, _07657_);
  or (_08196_, _08195_, _08193_);
  or (_08197_, _08196_, _08192_);
  or (_08198_, _08197_, _08189_);
  or (_08199_, _08198_, _08187_);
  and (_08200_, _08199_, _08184_);
  or (_08201_, _08189_, _08168_);
  or (_08202_, _08201_, _08200_);
  and (_08203_, _08202_, _08167_);
  and (_08204_, _08199_, _07923_);
  or (_08205_, _08204_, _07755_);
  not (_08206_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_08207_, _08120_, _08206_);
  or (_08208_, _08207_, _08156_);
  or (_08209_, _08208_, _08205_);
  or (_08210_, _08209_, _08203_);
  and (_06715_, _08210_, _05110_);
  and (_08211_, _07746_, _07936_);
  and (_08212_, _07988_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08213_, _08212_, _08211_);
  or (_08214_, _08186_, _07755_);
  and (_08215_, _08214_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08216_, _07841_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08217_, _07926_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08218_, _08217_, _08156_);
  or (_08219_, _08218_, _08216_);
  or (_08220_, _08219_, _08215_);
  or (_08221_, _08220_, _08168_);
  or (_08222_, _08221_, _08190_);
  or (_08223_, _08222_, _08213_);
  and (_06806_, _08223_, _05110_);
  not (_08224_, _05841_);
  and (_08225_, _06184_, _08224_);
  not (_08226_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_08227_, _06184_, _08226_);
  or (_08228_, _08227_, _08225_);
  and (_06855_, _08228_, _05110_);
  or (_08229_, _07926_, _07659_);
  and (_08230_, _08229_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08231_, _07988_, _07784_);
  and (_08232_, _08231_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_08233_, _08232_, _07981_);
  or (_08234_, _08233_, _08230_);
  and (_06900_, _08234_, _05110_);
  nor (_08235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_08236_, _08235_);
  nor (_08237_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_08238_, _08237_, _08236_);
  and (_08239_, _08238_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_08240_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_08241_, _08238_, _08240_);
  or (_08242_, _08241_, _08239_);
  and (_08243_, _06152_, _05789_);
  or (_08244_, _08243_, _08242_);
  and (_08245_, _06472_, _05782_);
  or (_08246_, _06472_, _08240_);
  nand (_08248_, _08246_, _08243_);
  or (_08249_, _08248_, _08245_);
  and (_08251_, _08249_, _08244_);
  and (_08252_, _05803_, _05434_);
  and (_08253_, _08252_, _05808_);
  or (_08254_, _08253_, _08251_);
  nand (_08255_, _08253_, _06229_);
  and (_08256_, _08255_, _05110_);
  and (_06961_, _08256_, _08254_);
  and (_08257_, _07206_, _05867_);
  or (_08258_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_08259_, _08258_, _05110_);
  nand (_08260_, _08257_, _05334_);
  and (_06965_, _08260_, _08259_);
  or (_08261_, _07992_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_06995_, _08261_, _05110_);
  and (_08262_, _05806_, _05403_);
  and (_08263_, _08252_, _08262_);
  and (_08264_, _08243_, _08133_);
  nand (_08265_, _08264_, _05872_);
  or (_08266_, _08264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_08267_, _08266_, _08265_);
  or (_08268_, _08267_, _08263_);
  nand (_08269_, _08253_, _06054_);
  and (_08270_, _08269_, _05110_);
  and (_07022_, _08270_, _08268_);
  and (_08272_, _06173_, _05911_);
  and (_08273_, _05807_, _08272_);
  and (_08274_, _08273_, _08252_);
  and (_08276_, _08274_, _08236_);
  and (_08277_, _08276_, _06799_);
  and (_08278_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_08280_, _08278_, _08235_);
  and (_08281_, _08236_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_08282_, _08281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_08283_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_08285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_08286_, _08285_, _08283_);
  and (_08287_, _08286_, _08282_);
  nor (_08288_, _08287_, _08280_);
  not (_08290_, _08288_);
  and (_08291_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_08292_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_08293_, _08292_, _08291_);
  nor (_08296_, _08293_, _08274_);
  and (_08297_, _08274_, _08235_);
  and (_08298_, _08297_, _06559_);
  or (_08300_, _08298_, _08296_);
  or (_08301_, _08300_, _08277_);
  and (_07036_, _08301_, _05110_);
  and (_08302_, _07305_, _06613_);
  nor (_08303_, _07337_, _06622_);
  and (_08304_, _08132_, _06472_);
  nand (_08305_, _08304_, _05872_);
  nor (_08306_, _08304_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_08307_, _08306_);
  and (_08308_, _08307_, _06638_);
  and (_08309_, _08308_, _08305_);
  or (_08310_, _08309_, _08303_);
  and (_08311_, _08310_, _06637_);
  or (_08312_, _08311_, _08302_);
  and (_07042_, _08312_, _05110_);
  and (_08313_, _08243_, _05488_);
  nand (_08314_, _08313_, _05872_);
  or (_08315_, _08313_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_08316_, _08315_, _08314_);
  or (_08317_, _08316_, _08263_);
  nand (_08318_, _08253_, _05841_);
  and (_08319_, _08318_, _05110_);
  and (_07047_, _08319_, _08317_);
  nor (_08320_, _05901_, _05465_);
  not (_08321_, _06174_);
  and (_08322_, _08321_, _06170_);
  and (_08323_, _08322_, _06168_);
  or (_08324_, _08323_, _05995_);
  not (_08325_, _06001_);
  nand (_08326_, _08325_, _06170_);
  nand (_08327_, _08326_, _05337_);
  nand (_08328_, _08327_, _06554_);
  or (_08329_, _08328_, _08324_);
  and (_08330_, _08329_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_08331_, _08330_, _08320_);
  and (_07102_, _08331_, _05110_);
  or (_08332_, _07813_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_07112_, _08332_, _05110_);
  nor (_08333_, _06229_, _06010_);
  not (_08334_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_08335_, _05997_, _08334_);
  or (_08336_, _08335_, _05995_);
  or (_08337_, _08336_, _08333_);
  or (_08338_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_08339_, _08338_, _05110_);
  and (_07166_, _08339_, _08337_);
  and (_08340_, _08282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  or (_08341_, _08340_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_08342_, _08340_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_08343_, _08342_, rst);
  nand (_08344_, _08343_, _08341_);
  nor (_07175_, _08344_, _08274_);
  or (_08345_, _08282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_08346_, _08340_, rst);
  nand (_08347_, _08346_, _08345_);
  nor (_07189_, _08347_, _08274_);
  and (_08348_, _07999_, _07923_);
  not (_08349_, _08348_);
  not (_08350_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_08351_, _08007_, _07618_);
  nor (_08352_, _08351_, _08004_);
  and (_08353_, _08007_, _07623_);
  and (_08354_, _08007_, _07612_);
  nor (_08355_, _08354_, _08353_);
  and (_08356_, _08355_, _08007_);
  and (_08357_, _08356_, _08352_);
  nor (_08358_, _08357_, _08350_);
  and (_08359_, _08357_, word_in[0]);
  or (_08360_, _08359_, _08358_);
  and (_08361_, _08360_, _08349_);
  and (_08362_, _08348_, word_in[8]);
  or (_08363_, _08362_, _08361_);
  and (_08364_, _07988_, _07775_);
  and (_08365_, _07993_, _08364_);
  not (_08366_, _08365_);
  and (_08367_, _08366_, _08363_);
  and (_08368_, _07988_, _07744_);
  and (_08369_, _08021_, _08368_);
  and (_08370_, _07993_, word_in[16]);
  and (_08371_, _08370_, _08364_);
  or (_08372_, _08371_, _08369_);
  or (_08373_, _08372_, _08367_);
  not (_08375_, _08369_);
  or (_08376_, _08375_, word_in[24]);
  and (_07468_, _08376_, _08373_);
  or (_08378_, _08357_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  not (_08379_, word_in[1]);
  nand (_08381_, _08357_, _08379_);
  and (_08383_, _08381_, _08349_);
  and (_08384_, _08383_, _08378_);
  and (_08385_, _07923_, word_in[9]);
  and (_08387_, _08385_, _07999_);
  or (_08388_, _08387_, _08365_);
  or (_08390_, _08388_, _08384_);
  nor (_08391_, _08366_, word_in[17]);
  nor (_08393_, _08391_, _08369_);
  and (_08394_, _08393_, _08390_);
  and (_08395_, _08021_, word_in[25]);
  and (_08397_, _08395_, _08369_);
  or (_07472_, _08397_, _08394_);
  not (_08398_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_08400_, _08357_, _08398_);
  and (_08401_, _08007_, word_in[2]);
  and (_08402_, _08401_, _08357_);
  or (_08403_, _08402_, _08400_);
  or (_08404_, _08403_, _08348_);
  or (_08405_, _08349_, word_in[10]);
  and (_08406_, _08405_, _08404_);
  or (_08407_, _08406_, _08365_);
  nor (_08408_, _08366_, word_in[18]);
  nor (_08409_, _08408_, _08369_);
  and (_08410_, _08409_, _08407_);
  and (_08411_, _08021_, word_in[26]);
  and (_08412_, _08411_, _08369_);
  or (_07476_, _08412_, _08410_);
  not (_08413_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_08414_, _08357_, _08413_);
  and (_08415_, _08007_, word_in[3]);
  and (_08416_, _08415_, _08357_);
  or (_08417_, _08416_, _08414_);
  or (_08418_, _08417_, _08348_);
  or (_08419_, _08349_, word_in[11]);
  and (_08420_, _08419_, _08418_);
  or (_08421_, _08420_, _08365_);
  nor (_08422_, _08366_, word_in[19]);
  nor (_08423_, _08422_, _08369_);
  and (_08424_, _08423_, _08421_);
  and (_08425_, _08021_, word_in[27]);
  and (_08426_, _08425_, _08369_);
  or (_07481_, _08426_, _08424_);
  not (_08427_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_08428_, _08357_, _08427_);
  and (_08429_, _08007_, word_in[4]);
  and (_08430_, _08429_, _08357_);
  or (_08431_, _08430_, _08428_);
  and (_08432_, _08431_, _08349_);
  and (_08433_, _08348_, word_in[12]);
  or (_08434_, _08433_, _08432_);
  or (_08435_, _08434_, _08365_);
  nor (_08436_, _08366_, word_in[20]);
  nor (_08437_, _08436_, _08369_);
  and (_08438_, _08437_, _08435_);
  and (_08439_, _08021_, word_in[28]);
  and (_08440_, _08439_, _08369_);
  or (_07484_, _08440_, _08438_);
  not (_08441_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_08442_, _08357_, _08441_);
  and (_08443_, _08007_, word_in[5]);
  and (_08444_, _08443_, _08357_);
  or (_08445_, _08444_, _08442_);
  or (_08446_, _08445_, _08348_);
  or (_08447_, _08349_, word_in[13]);
  and (_08448_, _08447_, _08446_);
  or (_08449_, _08448_, _08365_);
  nor (_08450_, _08366_, word_in[21]);
  nor (_08451_, _08450_, _08369_);
  and (_08452_, _08451_, _08449_);
  and (_08453_, _08021_, word_in[29]);
  and (_08454_, _08453_, _08369_);
  or (_07488_, _08454_, _08452_);
  not (_08455_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_08456_, _08357_, _08455_);
  and (_08457_, _08007_, word_in[6]);
  and (_08458_, _08457_, _08357_);
  or (_08459_, _08458_, _08456_);
  or (_08460_, _08459_, _08348_);
  or (_08461_, _08349_, word_in[14]);
  and (_08462_, _08461_, _08460_);
  or (_08463_, _08462_, _08365_);
  nor (_08464_, _08366_, word_in[22]);
  nor (_08466_, _08464_, _08369_);
  and (_08467_, _08466_, _08463_);
  and (_08469_, _08021_, word_in[30]);
  and (_08470_, _08469_, _08369_);
  or (_07491_, _08470_, _08467_);
  and (_08471_, _08369_, word_in[31]);
  nor (_08473_, _08357_, _07829_);
  and (_08474_, _08357_, word_in[7]);
  or (_08476_, _08474_, _08473_);
  and (_08478_, _08476_, _08349_);
  and (_08480_, _08348_, word_in[15]);
  or (_08481_, _08480_, _08478_);
  or (_08483_, _08481_, _08365_);
  nor (_08484_, _08366_, word_in[23]);
  nor (_08486_, _08484_, _08369_);
  and (_08487_, _08486_, _08483_);
  or (_07495_, _08487_, _08471_);
  and (_08488_, _08021_, _08364_);
  not (_08489_, _08488_);
  and (_08490_, _07993_, _07746_);
  and (_08491_, _08490_, _07868_);
  and (_08492_, _08491_, _08370_);
  and (_08493_, _07999_, _07783_);
  and (_08494_, _08493_, _07760_);
  and (_08495_, _08007_, word_in[0]);
  and (_08496_, _08004_, _07632_);
  and (_08497_, _08496_, _08355_);
  and (_08498_, _08497_, _08495_);
  not (_08499_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_08500_, _08497_, _08499_);
  or (_08501_, _08500_, _08498_);
  or (_08502_, _08501_, _08494_);
  not (_08503_, _08491_);
  not (_08504_, _08494_);
  or (_08505_, _08504_, word_in[8]);
  and (_08506_, _08505_, _08503_);
  and (_08507_, _08506_, _08502_);
  or (_08508_, _08507_, _08492_);
  and (_08509_, _08508_, _08489_);
  and (_08510_, _08488_, word_in[24]);
  or (_07573_, _08510_, _08509_);
  and (_08511_, _07993_, word_in[17]);
  and (_08512_, _08491_, _08511_);
  and (_08513_, _08007_, word_in[1]);
  and (_08514_, _08497_, _08513_);
  not (_08515_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_08516_, _08497_, _08515_);
  nor (_08517_, _08516_, _08514_);
  nor (_08518_, _08517_, _08494_);
  and (_08519_, _08494_, word_in[9]);
  or (_08520_, _08519_, _08518_);
  and (_08521_, _08520_, _08503_);
  or (_08522_, _08521_, _08512_);
  and (_08523_, _08522_, _08489_);
  and (_08524_, _08488_, word_in[25]);
  or (_07577_, _08524_, _08523_);
  and (_08525_, _07993_, word_in[18]);
  and (_08526_, _08491_, _08525_);
  and (_08527_, _08497_, _08401_);
  not (_08528_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_08529_, _08497_, _08528_);
  or (_08530_, _08529_, _08527_);
  or (_08531_, _08530_, _08494_);
  or (_08532_, _08504_, word_in[10]);
  and (_08533_, _08532_, _08503_);
  and (_08534_, _08533_, _08531_);
  or (_08535_, _08534_, _08526_);
  and (_08536_, _08535_, _08489_);
  and (_08537_, _08488_, word_in[26]);
  or (_07581_, _08537_, _08536_);
  not (_08538_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_08539_, _08497_, _08538_);
  and (_08540_, _08497_, _08415_);
  or (_08541_, _08540_, _08539_);
  or (_08542_, _08541_, _08494_);
  or (_08543_, _08504_, word_in[11]);
  and (_08544_, _08543_, _08542_);
  or (_08545_, _08544_, _08491_);
  and (_08546_, _07993_, word_in[19]);
  or (_08547_, _08503_, _08546_);
  and (_08548_, _08547_, _08489_);
  and (_08549_, _08548_, _08545_);
  and (_08551_, _08488_, word_in[27]);
  or (_07584_, _08551_, _08549_);
  not (_08553_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_08554_, _08497_, _08553_);
  and (_08555_, _08497_, _08429_);
  or (_08557_, _08555_, _08554_);
  or (_08558_, _08557_, _08494_);
  or (_08560_, _08504_, word_in[12]);
  and (_08561_, _08560_, _08558_);
  or (_08563_, _08561_, _08491_);
  and (_08564_, _07993_, word_in[20]);
  or (_08565_, _08503_, _08564_);
  and (_08567_, _08565_, _08489_);
  and (_08569_, _08567_, _08563_);
  and (_08570_, _08488_, word_in[28]);
  or (_07587_, _08570_, _08569_);
  and (_08572_, _07993_, word_in[21]);
  and (_08573_, _08491_, _08572_);
  and (_08574_, _08497_, _08443_);
  not (_08575_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_08576_, _08497_, _08575_);
  nor (_08577_, _08576_, _08574_);
  nor (_08578_, _08577_, _08494_);
  and (_08579_, _08494_, word_in[13]);
  or (_08580_, _08579_, _08578_);
  and (_08581_, _08580_, _08503_);
  or (_08582_, _08581_, _08573_);
  and (_08583_, _08582_, _08489_);
  and (_08584_, _08488_, word_in[29]);
  or (_07590_, _08584_, _08583_);
  not (_08585_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_08586_, _08497_, _08585_);
  and (_08587_, _08497_, _08457_);
  or (_08588_, _08587_, _08586_);
  or (_08589_, _08588_, _08494_);
  or (_08590_, _08504_, word_in[14]);
  and (_08591_, _08590_, _08589_);
  or (_08592_, _08591_, _08491_);
  and (_08593_, _07993_, word_in[22]);
  or (_08594_, _08503_, _08593_);
  and (_08595_, _08594_, _08489_);
  and (_08596_, _08595_, _08592_);
  and (_08597_, _08488_, word_in[30]);
  or (_07593_, _08597_, _08596_);
  and (_08598_, _08491_, _08023_);
  and (_08599_, _08497_, _08011_);
  nor (_08600_, _08497_, _07732_);
  or (_08601_, _08600_, _08599_);
  or (_08602_, _08601_, _08494_);
  or (_08603_, _08504_, word_in[15]);
  and (_08604_, _08603_, _08503_);
  and (_08605_, _08604_, _08602_);
  or (_08606_, _08605_, _08598_);
  and (_08607_, _08606_, _08489_);
  and (_08608_, _08488_, word_in[31]);
  or (_07597_, _08608_, _08607_);
  and (_08609_, _06559_, _05464_);
  and (_08610_, _08329_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  or (_08611_, _08610_, _08609_);
  and (_07639_, _08611_, _05110_);
  not (_08612_, _06004_);
  nand (_08613_, _05998_, _05337_);
  or (_08614_, _08613_, _08322_);
  or (_08615_, _08614_, _08612_);
  and (_08616_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_08617_, _06169_, _05337_);
  and (_08618_, _08617_, _06194_);
  or (_08619_, _08618_, _08616_);
  and (_07648_, _08619_, _05110_);
  and (_08620_, _08614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_08621_, _08617_, _06559_);
  nand (_08622_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_08623_, _08622_, _06004_);
  or (_08624_, _08623_, _08621_);
  or (_08625_, _08624_, _08620_);
  and (_07653_, _08625_, _05110_);
  not (_08626_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_08627_, _05464_, _08626_);
  nor (_08628_, _06088_, _05465_);
  or (_08629_, _08628_, _08627_);
  and (_07665_, _08629_, _05110_);
  and (_08630_, _07999_, _07744_);
  and (_08631_, _08630_, _07760_);
  not (_08632_, _08004_);
  and (_08633_, _08351_, _08632_);
  and (_08634_, _08633_, _08355_);
  and (_08635_, _08634_, _08495_);
  not (_08637_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_08638_, _08634_, _08637_);
  or (_08639_, _08638_, _08635_);
  or (_08641_, _08639_, _08631_);
  and (_08642_, _07993_, _07783_);
  and (_08643_, _08642_, _07868_);
  not (_08644_, _08643_);
  not (_08646_, _08631_);
  or (_08647_, _08646_, word_in[8]);
  and (_08648_, _08647_, _08644_);
  and (_08649_, _08648_, _08641_);
  and (_08651_, _08021_, _07746_);
  and (_08652_, _08651_, _07944_);
  and (_08653_, _08643_, _08370_);
  or (_08654_, _08653_, _08652_);
  or (_08655_, _08654_, _08649_);
  not (_08656_, _08652_);
  or (_08657_, _08656_, word_in[24]);
  and (_07686_, _08657_, _08655_);
  and (_08658_, _08634_, _08513_);
  not (_08659_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_08660_, _08634_, _08659_);
  or (_08661_, _08660_, _08658_);
  or (_08662_, _08661_, _08631_);
  or (_08663_, _08646_, word_in[9]);
  and (_08664_, _08663_, _08644_);
  and (_08665_, _08664_, _08662_);
  and (_08666_, _08643_, _08511_);
  or (_08667_, _08666_, _08652_);
  or (_08668_, _08667_, _08665_);
  or (_08669_, _08656_, word_in[25]);
  and (_07689_, _08669_, _08668_);
  and (_08670_, _08634_, _08401_);
  not (_08671_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_08672_, _08634_, _08671_);
  or (_08673_, _08672_, _08670_);
  or (_08674_, _08673_, _08631_);
  or (_08675_, _08646_, word_in[10]);
  and (_08676_, _08675_, _08644_);
  and (_08677_, _08676_, _08674_);
  and (_08678_, _08643_, _08525_);
  or (_08679_, _08678_, _08652_);
  or (_08680_, _08679_, _08677_);
  or (_08681_, _08656_, word_in[26]);
  and (_07692_, _08681_, _08680_);
  and (_08682_, _08634_, _08415_);
  not (_08683_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_08684_, _08634_, _08683_);
  or (_08685_, _08684_, _08682_);
  or (_08686_, _08685_, _08631_);
  or (_08687_, _08646_, word_in[11]);
  and (_08688_, _08687_, _08644_);
  and (_08689_, _08688_, _08686_);
  and (_08690_, _08643_, _08546_);
  or (_08691_, _08690_, _08652_);
  or (_08692_, _08691_, _08689_);
  or (_08693_, _08656_, word_in[27]);
  and (_07697_, _08693_, _08692_);
  and (_08694_, _08643_, _08564_);
  and (_08695_, _08634_, _08429_);
  not (_08696_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_08697_, _08634_, _08696_);
  nor (_08698_, _08697_, _08695_);
  nor (_08699_, _08698_, _08631_);
  and (_08700_, _08631_, word_in[12]);
  or (_08701_, _08700_, _08699_);
  and (_08702_, _08701_, _08644_);
  or (_08703_, _08702_, _08694_);
  and (_08704_, _08703_, _08656_);
  and (_08705_, _08652_, word_in[28]);
  or (_07700_, _08705_, _08704_);
  and (_08706_, _08643_, _08572_);
  and (_08707_, _08634_, _08443_);
  not (_08708_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_08709_, _08634_, _08708_);
  or (_08710_, _08709_, _08707_);
  or (_08711_, _08710_, _08631_);
  or (_08712_, _08646_, word_in[13]);
  and (_08713_, _08712_, _08644_);
  and (_08714_, _08713_, _08711_);
  or (_08715_, _08714_, _08706_);
  and (_08716_, _08715_, _08656_);
  and (_08717_, _08652_, word_in[29]);
  or (_07703_, _08717_, _08716_);
  not (_08718_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_08719_, _08634_, _08718_);
  and (_08720_, _08634_, _08457_);
  or (_08721_, _08720_, _08719_);
  or (_08722_, _08721_, _08631_);
  or (_08723_, _08646_, word_in[14]);
  and (_08724_, _08723_, _08722_);
  or (_08725_, _08724_, _08643_);
  nor (_08726_, _08644_, _08593_);
  nor (_08727_, _08726_, _08652_);
  and (_08728_, _08727_, _08725_);
  and (_08729_, _08652_, word_in[30]);
  or (_07708_, _08729_, _08728_);
  and (_08730_, _08643_, _08023_);
  and (_08731_, _08634_, _08011_);
  nor (_08732_, _08634_, _07834_);
  or (_08733_, _08732_, _08731_);
  or (_08734_, _08733_, _08631_);
  or (_08735_, _08646_, word_in[15]);
  and (_08736_, _08735_, _08644_);
  and (_08737_, _08736_, _08734_);
  or (_08738_, _08737_, _08730_);
  and (_08739_, _08738_, _08656_);
  and (_08740_, _08652_, word_in[31]);
  or (_07713_, _08740_, _08739_);
  not (_08741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_08742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_08743_, _08235_, _08742_);
  and (_08745_, _08743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_08746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_08748_, _08746_, _08236_);
  nor (_08749_, _08748_, _08745_);
  or (_08750_, _08749_, _08741_);
  and (_08751_, _08750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_08752_, _08745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_08753_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_08754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_08755_, _08754_, _08753_);
  and (_08756_, _08755_, _08752_);
  or (_08757_, _08756_, _08751_);
  and (_07758_, _08757_, _05110_);
  and (_08758_, _08021_, _08063_);
  not (_08759_, _08758_);
  and (_08760_, _07995_, _07868_);
  and (_08761_, _08760_, _08370_);
  and (_08762_, _08001_, _07760_);
  and (_08763_, _08355_, _08005_);
  and (_08764_, _08763_, _08495_);
  not (_08765_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_08766_, _08763_, _08765_);
  or (_08767_, _08766_, _08764_);
  or (_08768_, _08767_, _08762_);
  not (_08769_, _08760_);
  not (_08770_, _08762_);
  or (_08771_, _08770_, word_in[8]);
  and (_08772_, _08771_, _08769_);
  and (_08773_, _08772_, _08768_);
  or (_08774_, _08773_, _08761_);
  and (_08775_, _08774_, _08759_);
  and (_08776_, _08758_, word_in[24]);
  or (_07792_, _08776_, _08775_);
  and (_08777_, _08760_, _08511_);
  and (_08778_, _08763_, _08513_);
  not (_08779_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_08780_, _08763_, _08779_);
  or (_08781_, _08780_, _08778_);
  or (_08782_, _08781_, _08762_);
  or (_08783_, _08770_, word_in[9]);
  and (_08784_, _08783_, _08769_);
  and (_08785_, _08784_, _08782_);
  or (_08786_, _08785_, _08777_);
  and (_08787_, _08786_, _08759_);
  and (_08788_, _08758_, word_in[25]);
  or (_07795_, _08788_, _08787_);
  and (_08789_, _08760_, _08525_);
  and (_08790_, _08763_, _08401_);
  not (_08791_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_08792_, _08763_, _08791_);
  or (_08793_, _08792_, _08790_);
  or (_08794_, _08793_, _08762_);
  or (_08795_, _08770_, word_in[10]);
  and (_08796_, _08795_, _08769_);
  and (_08797_, _08796_, _08794_);
  or (_08798_, _08797_, _08789_);
  and (_08799_, _08798_, _08759_);
  and (_08800_, _08758_, word_in[26]);
  or (_07798_, _08800_, _08799_);
  and (_08801_, _08760_, _08546_);
  and (_08802_, _08763_, _08415_);
  not (_08803_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_08804_, _08763_, _08803_);
  or (_08805_, _08804_, _08802_);
  or (_08806_, _08805_, _08762_);
  or (_08807_, _08770_, word_in[11]);
  and (_08808_, _08807_, _08769_);
  and (_08809_, _08808_, _08806_);
  or (_08810_, _08809_, _08801_);
  and (_08811_, _08810_, _08759_);
  and (_08812_, _08758_, word_in[27]);
  or (_07803_, _08812_, _08811_);
  and (_08813_, _08760_, _08564_);
  and (_08814_, _08763_, _08429_);
  not (_08815_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_08816_, _08763_, _08815_);
  or (_08817_, _08816_, _08814_);
  or (_08818_, _08817_, _08762_);
  or (_08819_, _08770_, word_in[12]);
  and (_08820_, _08819_, _08769_);
  and (_08821_, _08820_, _08818_);
  or (_08822_, _08821_, _08813_);
  and (_08824_, _08822_, _08759_);
  and (_08825_, _08758_, word_in[28]);
  or (_07807_, _08825_, _08824_);
  and (_08827_, _08760_, _08572_);
  and (_08828_, _08763_, _08443_);
  not (_08830_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_08831_, _08763_, _08830_);
  or (_08833_, _08831_, _08828_);
  or (_08834_, _08833_, _08762_);
  or (_08836_, _08770_, word_in[13]);
  and (_08837_, _08836_, _08769_);
  and (_08838_, _08837_, _08834_);
  or (_08840_, _08838_, _08827_);
  and (_08841_, _08840_, _08759_);
  and (_08842_, _08758_, word_in[29]);
  or (_07812_, _08842_, _08841_);
  and (_08844_, _08758_, word_in[30]);
  and (_08845_, _08763_, _08457_);
  not (_08847_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_08848_, _08763_, _08847_);
  nor (_08849_, _08848_, _08845_);
  nor (_08850_, _08849_, _08762_);
  and (_08851_, _08762_, word_in[14]);
  or (_08852_, _08851_, _08850_);
  or (_08853_, _08852_, _08760_);
  or (_08854_, _08769_, _08593_);
  and (_08855_, _08854_, _08759_);
  and (_08856_, _08855_, _08853_);
  or (_07817_, _08856_, _08844_);
  and (_08857_, _08758_, word_in[31]);
  and (_08858_, _08763_, _08011_);
  nor (_08859_, _08763_, _07716_);
  nor (_08860_, _08859_, _08858_);
  nor (_08861_, _08860_, _08762_);
  and (_08862_, _08762_, word_in[15]);
  or (_08863_, _08862_, _08861_);
  or (_08864_, _08863_, _08760_);
  or (_08865_, _08769_, _08023_);
  and (_08866_, _08865_, _08759_);
  and (_08867_, _08866_, _08864_);
  or (_07822_, _08867_, _08857_);
  nand (_08868_, _06890_, _06054_);
  and (_08869_, _06061_, _05806_);
  and (_08870_, _08869_, _06888_);
  not (_08871_, _08870_);
  not (_08872_, _06883_);
  and (_08873_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_08874_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_08875_, _08874_, _08873_);
  or (_08876_, _08875_, _06890_);
  and (_08877_, _08876_, _08871_);
  and (_08878_, _08877_, _08868_);
  and (_08879_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_08880_, _08879_, _08878_);
  and (_07864_, _08880_, _05110_);
  nand (_08881_, _07337_, _06477_);
  or (_08882_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_08883_, _08882_, _05110_);
  and (_07867_, _08883_, _08881_);
  nor (_08884_, _06890_, _08872_);
  or (_08885_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  not (_08886_, _08884_);
  or (_08887_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_08888_, _08887_, _08885_);
  or (_08889_, _08888_, _08870_);
  nand (_08890_, _08870_, _06229_);
  and (_08891_, _08890_, _05110_);
  and (_07878_, _08891_, _08889_);
  nand (_08892_, _08870_, _06054_);
  or (_08893_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or (_08894_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_08895_, _08894_, _08893_);
  or (_08896_, _08895_, _08870_);
  and (_08897_, _08896_, _05110_);
  and (_07900_, _08897_, _08892_);
  and (_08898_, _08021_, _07930_);
  and (_08899_, _08898_, _07937_);
  and (_08900_, _08899_, _07744_);
  not (_08901_, _08900_);
  and (_08902_, _07993_, _08037_);
  not (_08903_, _08902_);
  and (_08904_, _07999_, _08042_);
  not (_08905_, _08904_);
  not (_08907_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_08908_, _08007_, _07754_);
  and (_08910_, _08908_, _08352_);
  nor (_08911_, _08910_, _08907_);
  and (_08912_, _08910_, word_in[0]);
  or (_08914_, _08912_, _08911_);
  and (_08915_, _08914_, _08905_);
  and (_08917_, _08904_, word_in[8]);
  or (_08918_, _08917_, _08915_);
  and (_08919_, _08918_, _08903_);
  and (_08921_, _08902_, word_in[16]);
  or (_08922_, _08921_, _08919_);
  and (_08924_, _08922_, _08901_);
  and (_08925_, _08021_, word_in[24]);
  and (_08927_, _08900_, _08925_);
  or (_07911_, _08927_, _08924_);
  or (_08928_, _08903_, word_in[17]);
  not (_08929_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_08930_, _08910_, _08929_);
  and (_08931_, _08910_, word_in[1]);
  or (_08932_, _08931_, _08930_);
  or (_08934_, _08932_, _08904_);
  or (_08935_, _08905_, word_in[9]);
  and (_08936_, _08935_, _08934_);
  or (_08937_, _08936_, _08902_);
  and (_08938_, _08937_, _08928_);
  or (_08939_, _08938_, _08900_);
  or (_08940_, _08901_, _08395_);
  and (_07915_, _08940_, _08939_);
  not (_08941_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_08942_, _08910_, _08941_);
  and (_08943_, _08910_, word_in[2]);
  or (_08944_, _08943_, _08942_);
  and (_08945_, _08944_, _08905_);
  and (_08946_, _08904_, word_in[10]);
  or (_08947_, _08946_, _08945_);
  and (_08948_, _08947_, _08903_);
  and (_08949_, _08902_, word_in[18]);
  or (_08950_, _08949_, _08900_);
  or (_08951_, _08950_, _08948_);
  or (_08952_, _08901_, _08411_);
  and (_07919_, _08952_, _08951_);
  not (_08953_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_08954_, _08910_, _08953_);
  and (_08955_, _08910_, word_in[3]);
  or (_08956_, _08955_, _08954_);
  and (_08957_, _08956_, _08905_);
  and (_08958_, _08904_, word_in[11]);
  or (_08959_, _08958_, _08957_);
  and (_08960_, _08959_, _08903_);
  and (_08961_, _08902_, word_in[19]);
  or (_08962_, _08961_, _08960_);
  and (_08963_, _08962_, _08901_);
  and (_08964_, _08900_, _08425_);
  or (_07922_, _08964_, _08963_);
  not (_08965_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_08966_, _08910_, _08965_);
  and (_08967_, _08910_, word_in[4]);
  or (_08968_, _08967_, _08966_);
  or (_08969_, _08968_, _08904_);
  or (_08970_, _08905_, word_in[12]);
  and (_08971_, _08970_, _08969_);
  or (_08972_, _08971_, _08902_);
  or (_08973_, _08903_, word_in[20]);
  and (_08974_, _08973_, _08972_);
  or (_08975_, _08974_, _08900_);
  or (_08976_, _08901_, _08439_);
  and (_07924_, _08976_, _08975_);
  not (_08977_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_08978_, _08910_, _08977_);
  and (_08979_, _08910_, word_in[5]);
  or (_08981_, _08979_, _08978_);
  or (_08982_, _08981_, _08904_);
  or (_08983_, _08905_, word_in[13]);
  and (_08984_, _08983_, _08982_);
  or (_08985_, _08984_, _08902_);
  nor (_08986_, _08903_, word_in[21]);
  nor (_08987_, _08986_, _08900_);
  and (_08988_, _08987_, _08985_);
  and (_08989_, _08900_, _08453_);
  or (_07928_, _08989_, _08988_);
  not (_08990_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_08991_, _08910_, _08990_);
  and (_08992_, _08910_, word_in[6]);
  or (_08993_, _08992_, _08991_);
  and (_08994_, _08993_, _08905_);
  and (_08995_, _08904_, word_in[14]);
  or (_08996_, _08995_, _08994_);
  and (_08997_, _08996_, _08903_);
  and (_08998_, _08902_, word_in[22]);
  or (_08999_, _08998_, _08900_);
  or (_09000_, _08999_, _08997_);
  or (_09001_, _08901_, _08469_);
  and (_07932_, _09001_, _09000_);
  nor (_09002_, _08910_, _07842_);
  and (_09003_, _08910_, word_in[7]);
  or (_09004_, _09003_, _09002_);
  and (_09005_, _09004_, _08905_);
  and (_09006_, _08904_, word_in[15]);
  or (_09007_, _09006_, _09005_);
  and (_09008_, _09007_, _08903_);
  and (_09009_, _08902_, _08023_);
  or (_09010_, _09009_, _08900_);
  or (_09011_, _09010_, _09008_);
  or (_09012_, _08901_, _08028_);
  and (_07934_, _09012_, _09011_);
  and (_09013_, _08899_, _07775_);
  not (_09014_, _09013_);
  and (_09015_, _07993_, _07858_);
  and (_09016_, _09015_, _07907_);
  and (_09017_, _09016_, _07746_);
  not (_09018_, _09017_);
  or (_09019_, _09018_, _08370_);
  and (_09020_, _08493_, _07841_);
  not (_09021_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_09022_, _08908_, _08496_);
  nor (_09023_, _09022_, _09021_);
  and (_09024_, _09022_, word_in[0]);
  or (_09025_, _09024_, _09023_);
  or (_09026_, _09025_, _09020_);
  not (_09027_, _09020_);
  or (_09028_, _09027_, word_in[8]);
  and (_09029_, _09028_, _09026_);
  or (_09030_, _09029_, _09017_);
  and (_09031_, _09030_, _09019_);
  and (_09032_, _09031_, _09014_);
  and (_09033_, _09013_, word_in[24]);
  or (_07991_, _09033_, _09032_);
  and (_09034_, _09022_, word_in[1]);
  not (_09035_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_09036_, _09022_, _09035_);
  nor (_09037_, _09036_, _09034_);
  nor (_09038_, _09037_, _09020_);
  and (_09039_, _09020_, word_in[9]);
  or (_09040_, _09039_, _09038_);
  and (_09041_, _09040_, _09018_);
  and (_09042_, _09017_, _08511_);
  or (_09043_, _09042_, _09013_);
  or (_09044_, _09043_, _09041_);
  or (_09045_, _09014_, word_in[25]);
  and (_07994_, _09045_, _09044_);
  and (_09046_, _09017_, _08525_);
  and (_09047_, _09022_, word_in[2]);
  not (_09048_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_09049_, _09022_, _09048_);
  nor (_09050_, _09049_, _09047_);
  nor (_09051_, _09050_, _09020_);
  and (_09052_, _09020_, word_in[10]);
  or (_09053_, _09052_, _09051_);
  and (_09054_, _09053_, _09018_);
  or (_09055_, _09054_, _09046_);
  and (_09056_, _09055_, _09014_);
  and (_09057_, _09013_, word_in[26]);
  or (_07997_, _09057_, _09056_);
  or (_09058_, _09018_, _08546_);
  not (_09059_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_09060_, _09022_, _09059_);
  and (_09061_, _09022_, word_in[3]);
  or (_09062_, _09061_, _09060_);
  or (_09063_, _09062_, _09020_);
  or (_09064_, _09027_, word_in[11]);
  and (_09065_, _09064_, _09063_);
  or (_09066_, _09065_, _09017_);
  and (_09067_, _09066_, _09058_);
  or (_09068_, _09067_, _09013_);
  or (_09069_, _09014_, word_in[27]);
  and (_08000_, _09069_, _09068_);
  and (_09070_, _09022_, word_in[4]);
  not (_09071_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_09072_, _09022_, _09071_);
  nor (_09073_, _09072_, _09070_);
  nor (_09074_, _09073_, _09020_);
  and (_09075_, _09020_, word_in[12]);
  or (_09076_, _09075_, _09074_);
  and (_09077_, _09076_, _09018_);
  and (_09078_, _09017_, _08564_);
  or (_09079_, _09078_, _09013_);
  or (_09080_, _09079_, _09077_);
  or (_09081_, _09014_, word_in[28]);
  and (_08003_, _09081_, _09080_);
  not (_09082_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_09083_, _09022_, _09082_);
  and (_09084_, _09022_, word_in[5]);
  nor (_09085_, _09084_, _09083_);
  nor (_09086_, _09085_, _09020_);
  and (_09087_, _09020_, word_in[13]);
  or (_09088_, _09087_, _09086_);
  and (_09089_, _09088_, _09018_);
  and (_09090_, _09017_, _08572_);
  or (_09091_, _09090_, _09013_);
  or (_09092_, _09091_, _09089_);
  or (_09093_, _09014_, word_in[29]);
  and (_08006_, _09093_, _09092_);
  and (_09094_, _09022_, word_in[6]);
  not (_09095_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_09096_, _09022_, _09095_);
  nor (_09097_, _09096_, _09094_);
  nor (_09098_, _09097_, _09020_);
  and (_09099_, _09020_, word_in[14]);
  or (_09100_, _09099_, _09098_);
  and (_09101_, _09100_, _09018_);
  and (_09102_, _09017_, _08593_);
  or (_09103_, _09102_, _09013_);
  or (_09104_, _09103_, _09101_);
  or (_09105_, _09014_, word_in[30]);
  and (_08009_, _09105_, _09104_);
  and (_09106_, _09017_, _08023_);
  and (_09107_, _09022_, word_in[7]);
  nor (_09108_, _09022_, _07727_);
  nor (_09109_, _09108_, _09107_);
  nor (_09110_, _09109_, _09020_);
  and (_09111_, _09020_, word_in[15]);
  or (_09112_, _09111_, _09110_);
  and (_09113_, _09112_, _09018_);
  or (_09114_, _09113_, _09106_);
  and (_09115_, _09114_, _09014_);
  and (_09116_, _09013_, word_in[31]);
  or (_08012_, _09116_, _09115_);
  and (_09117_, _08630_, _07841_);
  not (_09118_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_09119_, _08633_, _07754_);
  nor (_09120_, _09119_, _09118_);
  and (_09121_, _09119_, _08495_);
  or (_09122_, _09121_, _09120_);
  or (_09123_, _09122_, _09117_);
  and (_09124_, _09016_, _07783_);
  not (_09125_, _09124_);
  not (_09126_, _09117_);
  or (_09127_, _09126_, word_in[8]);
  and (_09128_, _09127_, _09125_);
  and (_09129_, _09128_, _09123_);
  and (_09130_, _08899_, _07746_);
  and (_09131_, _09124_, _08370_);
  or (_09132_, _09131_, _09130_);
  or (_09133_, _09132_, _09129_);
  not (_09134_, _09130_);
  or (_09135_, _09134_, word_in[24]);
  and (_08077_, _09135_, _09133_);
  not (_09136_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_09137_, _09119_, _09136_);
  and (_09138_, _09119_, _08513_);
  nor (_09139_, _09138_, _09137_);
  nor (_09140_, _09139_, _09117_);
  and (_09141_, _09117_, word_in[9]);
  or (_09142_, _09141_, _09140_);
  and (_09143_, _09142_, _09125_);
  and (_09144_, _09124_, _08511_);
  or (_09145_, _09144_, _09130_);
  or (_09146_, _09145_, _09143_);
  or (_09147_, _09134_, word_in[25]);
  and (_08080_, _09147_, _09146_);
  not (_09148_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_09149_, _09119_, _09148_);
  and (_09150_, _09119_, _08401_);
  or (_09151_, _09150_, _09149_);
  or (_09152_, _09151_, _09117_);
  or (_09153_, _09126_, word_in[10]);
  and (_09154_, _09153_, _09125_);
  and (_09155_, _09154_, _09152_);
  and (_09156_, _09124_, _08525_);
  or (_09157_, _09156_, _09130_);
  or (_09158_, _09157_, _09155_);
  or (_09159_, _09134_, word_in[26]);
  and (_08084_, _09159_, _09158_);
  not (_09160_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_09161_, _09119_, _09160_);
  and (_09162_, _09119_, _08415_);
  or (_09163_, _09162_, _09161_);
  or (_09164_, _09163_, _09117_);
  or (_09165_, _09126_, word_in[11]);
  and (_09166_, _09165_, _09125_);
  and (_09167_, _09166_, _09164_);
  and (_09168_, _09124_, _08546_);
  or (_09169_, _09168_, _09130_);
  or (_09170_, _09169_, _09167_);
  or (_09171_, _09134_, word_in[27]);
  and (_08089_, _09171_, _09170_);
  not (_09172_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_09173_, _09119_, _09172_);
  and (_09174_, _09119_, _08429_);
  or (_09175_, _09174_, _09173_);
  or (_09176_, _09175_, _09117_);
  or (_09177_, _09126_, word_in[12]);
  and (_09178_, _09177_, _09125_);
  and (_09179_, _09178_, _09176_);
  and (_09180_, _09124_, _08564_);
  or (_09181_, _09180_, _09130_);
  or (_09182_, _09181_, _09179_);
  or (_09183_, _09134_, word_in[28]);
  and (_08091_, _09183_, _09182_);
  not (_09184_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_09185_, _09119_, _09184_);
  and (_09186_, _09119_, _08443_);
  or (_09187_, _09186_, _09185_);
  or (_09188_, _09187_, _09117_);
  or (_09189_, _09126_, word_in[13]);
  and (_09190_, _09189_, _09125_);
  and (_09191_, _09190_, _09188_);
  and (_09192_, _09124_, _08572_);
  or (_09193_, _09192_, _09130_);
  or (_09194_, _09193_, _09191_);
  or (_09195_, _09134_, word_in[29]);
  and (_08094_, _09195_, _09194_);
  or (_09196_, _09125_, _08593_);
  not (_09197_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_09198_, _09119_, _09197_);
  and (_09199_, _09119_, _08457_);
  or (_09200_, _09199_, _09198_);
  or (_09201_, _09200_, _09117_);
  or (_09202_, _09126_, word_in[14]);
  and (_09203_, _09202_, _09201_);
  or (_09204_, _09203_, _09124_);
  and (_09205_, _09204_, _09196_);
  or (_09206_, _09205_, _09130_);
  or (_09207_, _09134_, word_in[30]);
  and (_08098_, _09207_, _09206_);
  or (_09208_, _09125_, _08023_);
  nor (_09209_, _09119_, _07847_);
  and (_09210_, _09119_, _08011_);
  or (_09211_, _09210_, _09209_);
  or (_09212_, _09211_, _09117_);
  or (_09213_, _09126_, word_in[15]);
  and (_09214_, _09213_, _09212_);
  or (_09215_, _09214_, _09124_);
  and (_09216_, _09215_, _09208_);
  or (_09217_, _09216_, _09130_);
  or (_09218_, _09134_, word_in[31]);
  and (_08103_, _09218_, _09217_);
  and (_09219_, _09016_, _07744_);
  not (_09220_, _09219_);
  and (_09221_, _08001_, _07841_);
  not (_09222_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_09223_, _08908_, _08005_);
  nor (_09224_, _09223_, _09222_);
  and (_09225_, _09223_, word_in[0]);
  nor (_09226_, _09225_, _09224_);
  nor (_09227_, _09226_, _09221_);
  and (_09228_, _09221_, word_in[8]);
  or (_09229_, _09228_, _09227_);
  and (_09230_, _09229_, _09220_);
  and (_09232_, _08021_, _08059_);
  and (_09233_, _09219_, _08370_);
  or (_09235_, _09233_, _09232_);
  or (_09236_, _09235_, _09230_);
  not (_09237_, _09232_);
  or (_09238_, _09237_, _08925_);
  and (_08171_, _09238_, _09236_);
  not (_09239_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_09240_, _09223_, _09239_);
  and (_09241_, _09223_, word_in[1]);
  nor (_09242_, _09241_, _09240_);
  nor (_09244_, _09242_, _09221_);
  and (_09245_, _09221_, word_in[9]);
  or (_09246_, _09245_, _09244_);
  and (_09247_, _09246_, _09220_);
  and (_09248_, _09219_, _08511_);
  or (_09249_, _09248_, _09232_);
  or (_09250_, _09249_, _09247_);
  or (_09251_, _09237_, _08395_);
  and (_08175_, _09251_, _09250_);
  not (_09252_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_09253_, _09223_, _09252_);
  and (_09254_, _09223_, word_in[2]);
  nor (_09255_, _09254_, _09253_);
  nor (_09256_, _09255_, _09221_);
  and (_09257_, _09221_, word_in[10]);
  or (_09258_, _09257_, _09256_);
  and (_09259_, _09258_, _09220_);
  and (_09260_, _09219_, _08525_);
  or (_09261_, _09260_, _09232_);
  or (_09262_, _09261_, _09259_);
  or (_09263_, _09237_, _08411_);
  and (_13444_, _09263_, _09262_);
  not (_09264_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_09265_, _09223_, _09264_);
  and (_09266_, _09223_, word_in[3]);
  nor (_09267_, _09266_, _09265_);
  nor (_09268_, _09267_, _09221_);
  and (_09269_, _09221_, word_in[11]);
  or (_09270_, _09269_, _09268_);
  and (_09271_, _09270_, _09220_);
  and (_09272_, _09219_, _08546_);
  or (_09273_, _09272_, _09232_);
  or (_09274_, _09273_, _09271_);
  or (_09275_, _09237_, _08425_);
  and (_13445_, _09275_, _09274_);
  not (_09276_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_09277_, _09223_, _09276_);
  and (_09278_, _09223_, word_in[4]);
  nor (_09279_, _09278_, _09277_);
  nor (_09280_, _09279_, _09221_);
  and (_09281_, _09221_, word_in[12]);
  or (_09282_, _09281_, _09280_);
  and (_09283_, _09282_, _09220_);
  and (_09284_, _09219_, _08564_);
  or (_09285_, _09284_, _09232_);
  or (_09286_, _09285_, _09283_);
  or (_09287_, _09237_, _08439_);
  and (_13446_, _09287_, _09286_);
  not (_09288_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_09289_, _09223_, _09288_);
  and (_09290_, _09223_, word_in[5]);
  nor (_09291_, _09290_, _09289_);
  nor (_09292_, _09291_, _09221_);
  and (_09293_, _09221_, word_in[13]);
  or (_09294_, _09293_, _09292_);
  and (_09295_, _09294_, _09220_);
  and (_09296_, _09219_, _08572_);
  or (_09297_, _09296_, _09232_);
  or (_09298_, _09297_, _09295_);
  or (_09299_, _09237_, _08453_);
  and (_13447_, _09299_, _09298_);
  not (_09300_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_09301_, _09223_, _09300_);
  and (_09302_, _09223_, word_in[6]);
  nor (_09303_, _09302_, _09301_);
  nor (_09304_, _09303_, _09221_);
  and (_09305_, _09221_, word_in[14]);
  or (_09306_, _09305_, _09304_);
  and (_09307_, _09306_, _09220_);
  and (_09308_, _09219_, _08593_);
  or (_09309_, _09308_, _09232_);
  or (_09310_, _09309_, _09307_);
  or (_09311_, _09237_, _08469_);
  and (_13448_, _09311_, _09310_);
  nor (_09312_, _09223_, _07721_);
  and (_09313_, _09223_, word_in[7]);
  nor (_09314_, _09313_, _09312_);
  nor (_09315_, _09314_, _09221_);
  and (_09316_, _09221_, word_in[15]);
  or (_09317_, _09316_, _09315_);
  and (_09318_, _09317_, _09220_);
  and (_09319_, _09219_, _08023_);
  or (_09320_, _09319_, _09232_);
  or (_09321_, _09320_, _09318_);
  or (_09322_, _09237_, _08028_);
  and (_08185_, _09322_, _09321_);
  nor (_09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_09324_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _05110_);
  and (_09326_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_08247_, _09326_, _09324_);
  nor (_09327_, _08342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_09328_, _08342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_09329_, _09328_, _09327_);
  nand (_09330_, _09329_, _05110_);
  nor (_08250_, _09330_, _08274_);
  and (_09331_, _07993_, _08096_);
  not (_09332_, _09331_);
  and (_09333_, _07999_, _07755_);
  not (_09334_, _09333_);
  not (_09335_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_09336_, _08354_, _07753_);
  and (_09337_, _09336_, _08352_);
  nor (_09338_, _09337_, _09335_);
  and (_09339_, _09337_, _08495_);
  or (_09340_, _09339_, _09338_);
  and (_09341_, _09340_, _09334_);
  and (_09342_, _09333_, word_in[8]);
  or (_09343_, _09342_, _09341_);
  and (_09344_, _09343_, _09332_);
  and (_09345_, _08021_, _08074_);
  and (_09346_, _09331_, word_in[16]);
  or (_09347_, _09346_, _09345_);
  or (_09348_, _09347_, _09344_);
  not (_09349_, _09345_);
  or (_09350_, _09349_, _08925_);
  and (_13449_, _09350_, _09348_);
  not (_09351_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_09352_, _09337_, _09351_);
  and (_09353_, _09337_, _08513_);
  or (_09354_, _09353_, _09352_);
  and (_09355_, _09354_, _09334_);
  and (_09356_, _09333_, word_in[9]);
  or (_09357_, _09356_, _09355_);
  and (_09358_, _09357_, _09332_);
  and (_09359_, _09331_, word_in[17]);
  or (_09360_, _09359_, _09358_);
  and (_09361_, _09360_, _09349_);
  and (_09362_, _09345_, word_in[25]);
  or (_08271_, _09362_, _09361_);
  not (_09363_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_09364_, _09337_, _09363_);
  and (_09365_, _09337_, _08401_);
  or (_09366_, _09365_, _09364_);
  and (_09367_, _09366_, _09334_);
  and (_09368_, _09333_, word_in[10]);
  or (_09369_, _09368_, _09367_);
  and (_09370_, _09369_, _09332_);
  and (_09371_, _09331_, word_in[18]);
  or (_09372_, _09371_, _09370_);
  and (_09373_, _09372_, _09349_);
  and (_09374_, _09345_, word_in[26]);
  or (_08275_, _09374_, _09373_);
  not (_09375_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_09376_, _09337_, _09375_);
  and (_09377_, _09337_, _08415_);
  or (_09378_, _09377_, _09376_);
  and (_09379_, _09378_, _09334_);
  and (_09380_, _09333_, word_in[11]);
  or (_09381_, _09380_, _09379_);
  and (_09382_, _09381_, _09332_);
  and (_09383_, _09331_, word_in[19]);
  or (_09384_, _09383_, _09345_);
  or (_09385_, _09384_, _09382_);
  or (_09386_, _09349_, _08425_);
  and (_08279_, _09386_, _09385_);
  not (_09387_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_09388_, _09337_, _09387_);
  and (_09389_, _09337_, _08429_);
  or (_09390_, _09389_, _09388_);
  and (_09391_, _09390_, _09334_);
  and (_09392_, _09333_, word_in[12]);
  or (_09393_, _09392_, _09391_);
  and (_09394_, _09393_, _09332_);
  and (_09395_, _09331_, word_in[20]);
  or (_09396_, _09395_, _09345_);
  or (_09397_, _09396_, _09394_);
  or (_09398_, _09349_, _08439_);
  and (_08284_, _09398_, _09397_);
  not (_09399_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_09400_, _09337_, _09399_);
  and (_09401_, _09337_, _08443_);
  or (_09402_, _09401_, _09400_);
  and (_09403_, _09402_, _09334_);
  and (_09404_, _09333_, word_in[13]);
  or (_09405_, _09404_, _09403_);
  and (_09406_, _09405_, _09332_);
  and (_09407_, _09331_, word_in[21]);
  or (_09408_, _09407_, _09406_);
  and (_09409_, _09408_, _09349_);
  and (_09410_, _09345_, word_in[29]);
  or (_08289_, _09410_, _09409_);
  not (_09411_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_09412_, _09337_, _09411_);
  and (_09413_, _09337_, _08457_);
  or (_09414_, _09413_, _09412_);
  and (_09415_, _09414_, _09334_);
  and (_09416_, _09333_, word_in[14]);
  or (_09417_, _09416_, _09415_);
  and (_09418_, _09417_, _09332_);
  and (_09419_, _09331_, word_in[22]);
  or (_09420_, _09419_, _09418_);
  and (_09421_, _09420_, _09349_);
  and (_09422_, _09345_, word_in[30]);
  or (_08295_, _09422_, _09421_);
  and (_09423_, _09331_, word_in[23]);
  nor (_09424_, _09337_, _07804_);
  and (_09425_, _09337_, _08011_);
  or (_09426_, _09425_, _09424_);
  and (_09427_, _09426_, _09334_);
  and (_09428_, _09333_, word_in[15]);
  or (_09429_, _09428_, _09427_);
  and (_09430_, _09429_, _09332_);
  or (_09431_, _09430_, _09423_);
  and (_09432_, _09431_, _09349_);
  and (_09433_, _09345_, word_in[31]);
  or (_08299_, _09433_, _09432_);
  and (_09434_, _08490_, _07865_);
  and (_09435_, _08493_, _07757_);
  not (_09436_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_09437_, _09336_, _08496_);
  nor (_09438_, _09437_, _09436_);
  and (_09439_, _09437_, _08495_);
  or (_09440_, _09439_, _09438_);
  or (_09441_, _09440_, _09435_);
  not (_09442_, _09435_);
  or (_09443_, _09442_, word_in[8]);
  and (_09444_, _09443_, _09441_);
  or (_09445_, _09444_, _09434_);
  and (_09446_, _08021_, _07938_);
  and (_09447_, _09446_, _07775_);
  not (_09448_, _09434_);
  nor (_09449_, _09448_, _08370_);
  nor (_09450_, _09449_, _09447_);
  and (_09451_, _09450_, _09445_);
  and (_09452_, _09447_, _08925_);
  or (_08374_, _09452_, _09451_);
  not (_09453_, _09447_);
  and (_09454_, _09434_, _08511_);
  and (_09455_, _09437_, _08513_);
  not (_09456_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_09457_, _09437_, _09456_);
  or (_09458_, _09457_, _09455_);
  or (_09459_, _09458_, _09435_);
  or (_09460_, _09442_, word_in[9]);
  and (_09461_, _09460_, _09448_);
  and (_09462_, _09461_, _09459_);
  or (_09463_, _09462_, _09454_);
  and (_09464_, _09463_, _09453_);
  and (_09465_, _09447_, word_in[25]);
  or (_08377_, _09465_, _09464_);
  or (_09466_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not (_09467_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_09468_, _06205_, _09467_);
  and (_09469_, _09468_, _05110_);
  and (_08380_, _09469_, _09466_);
  and (_09470_, _09437_, _08401_);
  not (_09471_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_09472_, _09437_, _09471_);
  or (_09473_, _09472_, _09470_);
  or (_09474_, _09473_, _09435_);
  or (_09475_, _09442_, word_in[10]);
  and (_09476_, _09475_, _09448_);
  and (_09477_, _09476_, _09474_);
  and (_09478_, _09434_, _08525_);
  or (_09479_, _09478_, _09447_);
  or (_09480_, _09479_, _09477_);
  or (_09481_, _09453_, _08411_);
  and (_08382_, _09481_, _09480_);
  not (_09482_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_09483_, _09437_, _09482_);
  and (_09484_, _09437_, _08415_);
  or (_09485_, _09484_, _09483_);
  or (_09486_, _09485_, _09435_);
  or (_09487_, _09442_, word_in[11]);
  and (_09488_, _09487_, _09486_);
  or (_09489_, _09488_, _09434_);
  nor (_09490_, _09448_, _08546_);
  nor (_09491_, _09490_, _09447_);
  and (_09492_, _09491_, _09489_);
  and (_09493_, _09447_, _08425_);
  or (_08386_, _09493_, _09492_);
  not (_09494_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_09495_, _09437_, _09494_);
  and (_09496_, _09437_, _08429_);
  or (_09497_, _09496_, _09495_);
  or (_09498_, _09497_, _09435_);
  or (_09499_, _09442_, word_in[12]);
  and (_09500_, _09499_, _09498_);
  or (_09501_, _09500_, _09434_);
  nor (_09502_, _09448_, _08564_);
  nor (_09503_, _09502_, _09447_);
  and (_09504_, _09503_, _09501_);
  and (_09505_, _09447_, _08439_);
  or (_08389_, _09505_, _09504_);
  not (_09506_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_09507_, _09437_, _09506_);
  and (_09508_, _09437_, _08443_);
  or (_09509_, _09508_, _09507_);
  or (_09510_, _09509_, _09435_);
  or (_09511_, _09442_, word_in[13]);
  and (_09512_, _09511_, _09510_);
  or (_09513_, _09512_, _09434_);
  nor (_09514_, _09448_, _08572_);
  nor (_09515_, _09514_, _09447_);
  and (_09516_, _09515_, _09513_);
  and (_09517_, _09447_, _08453_);
  or (_08392_, _09517_, _09516_);
  not (_09518_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_09519_, _09437_, _09518_);
  and (_09520_, _09437_, _08457_);
  or (_09521_, _09520_, _09519_);
  or (_09522_, _09521_, _09435_);
  or (_09523_, _09442_, word_in[14]);
  and (_09524_, _09523_, _09522_);
  or (_09525_, _09524_, _09434_);
  nor (_09526_, _09448_, _08593_);
  nor (_09527_, _09526_, _09447_);
  and (_09528_, _09527_, _09525_);
  and (_09529_, _09447_, _08469_);
  or (_08396_, _09529_, _09528_);
  nor (_09530_, _09437_, _07706_);
  and (_09531_, _09437_, _08011_);
  or (_09532_, _09531_, _09530_);
  or (_09533_, _09532_, _09435_);
  or (_09534_, _09442_, word_in[15]);
  and (_09535_, _09534_, _09533_);
  or (_09536_, _09535_, _09434_);
  nor (_09537_, _09448_, _08023_);
  nor (_09538_, _09537_, _09447_);
  and (_09539_, _09538_, _09536_);
  and (_09540_, _09447_, _08028_);
  or (_08399_, _09540_, _09539_);
  and (_09541_, _08642_, _07865_);
  and (_09542_, _08630_, _07757_);
  not (_09543_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_09544_, _09336_, _08633_);
  nor (_09545_, _09544_, _09543_);
  and (_09546_, _09544_, _08495_);
  or (_09547_, _09546_, _09545_);
  or (_09548_, _09547_, _09542_);
  not (_09549_, _09542_);
  or (_09550_, _09549_, word_in[8]);
  and (_09551_, _09550_, _09548_);
  or (_09552_, _09551_, _09541_);
  and (_09553_, _09446_, _07746_);
  not (_09554_, _09541_);
  nor (_09555_, _09554_, _08370_);
  nor (_09556_, _09555_, _09553_);
  and (_09557_, _09556_, _09552_);
  and (_09558_, _09553_, _08925_);
  or (_08465_, _09558_, _09557_);
  not (_09559_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_09560_, _09544_, _09559_);
  and (_09561_, _09544_, _08513_);
  or (_09562_, _09561_, _09560_);
  or (_09563_, _09562_, _09542_);
  or (_09564_, _09549_, word_in[9]);
  and (_09565_, _09564_, _09563_);
  or (_09566_, _09565_, _09541_);
  nor (_09567_, _09554_, _08511_);
  nor (_09568_, _09567_, _09553_);
  and (_09569_, _09568_, _09566_);
  and (_09570_, _09553_, _08395_);
  or (_08468_, _09570_, _09569_);
  and (_09571_, _09544_, _08401_);
  not (_09572_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_09573_, _09544_, _09572_);
  or (_09574_, _09573_, _09571_);
  or (_09575_, _09574_, _09542_);
  or (_09576_, _09549_, word_in[10]);
  and (_09577_, _09576_, _09554_);
  and (_09578_, _09577_, _09575_);
  and (_09579_, _09541_, _08525_);
  or (_09580_, _09579_, _09553_);
  or (_09581_, _09580_, _09578_);
  not (_09582_, _09553_);
  or (_09583_, _09582_, _08411_);
  and (_08472_, _09583_, _09581_);
  and (_09584_, _09544_, _08415_);
  not (_09585_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_09586_, _09544_, _09585_);
  or (_09587_, _09586_, _09584_);
  or (_09588_, _09587_, _09542_);
  or (_09589_, _09549_, word_in[11]);
  and (_09590_, _09589_, _09554_);
  and (_09591_, _09590_, _09588_);
  and (_09592_, _09541_, _08546_);
  or (_09593_, _09592_, _09553_);
  or (_09594_, _09593_, _09591_);
  or (_09595_, _09582_, _08425_);
  and (_08475_, _09595_, _09594_);
  and (_09596_, _09541_, _08564_);
  and (_09597_, _09544_, _08429_);
  not (_09598_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_09599_, _09544_, _09598_);
  or (_09600_, _09599_, _09597_);
  or (_09601_, _09600_, _09542_);
  or (_09602_, _09549_, word_in[12]);
  and (_09603_, _09602_, _09554_);
  and (_09604_, _09603_, _09601_);
  or (_09605_, _09604_, _09596_);
  and (_09606_, _09605_, _09582_);
  and (_09607_, _09553_, word_in[28]);
  or (_08477_, _09607_, _09606_);
  not (_09608_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_09609_, _09544_, _09608_);
  and (_09610_, _09544_, _08443_);
  or (_09611_, _09610_, _09609_);
  or (_09612_, _09611_, _09542_);
  or (_09613_, _09549_, word_in[13]);
  and (_09614_, _09613_, _09612_);
  or (_09615_, _09614_, _09541_);
  nor (_09616_, _09554_, _08572_);
  nor (_09617_, _09616_, _09553_);
  and (_09618_, _09617_, _09615_);
  and (_09619_, _09553_, _08453_);
  or (_08479_, _09619_, _09618_);
  and (_09620_, _09544_, _08457_);
  not (_09621_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_09622_, _09544_, _09621_);
  or (_09623_, _09622_, _09620_);
  or (_09624_, _09623_, _09542_);
  or (_09625_, _09549_, word_in[14]);
  and (_09626_, _09625_, _09554_);
  and (_09627_, _09626_, _09624_);
  and (_09628_, _09541_, _08593_);
  or (_09630_, _09628_, _09553_);
  or (_09631_, _09630_, _09627_);
  or (_09632_, _09582_, _08469_);
  and (_08482_, _09632_, _09631_);
  and (_09634_, _09541_, _08023_);
  and (_09635_, _09544_, _08011_);
  nor (_09637_, _09544_, _07797_);
  nor (_09638_, _09637_, _09635_);
  nor (_09640_, _09638_, _09542_);
  and (_09641_, _09542_, word_in[15]);
  or (_09642_, _09641_, _09640_);
  and (_09643_, _09642_, _09554_);
  or (_09644_, _09643_, _09634_);
  and (_09645_, _09644_, _09582_);
  and (_09646_, _09553_, word_in[31]);
  or (_08485_, _09646_, _09645_);
  and (_09647_, _07995_, _07865_);
  and (_09648_, _08001_, _07757_);
  not (_09649_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_09650_, _09336_, _08005_);
  nor (_09651_, _09650_, _09649_);
  and (_09652_, _09650_, _08495_);
  or (_09653_, _09652_, _09651_);
  or (_09654_, _09653_, _09648_);
  not (_09655_, _09648_);
  or (_09656_, _09655_, word_in[8]);
  and (_09657_, _09656_, _09654_);
  or (_09658_, _09657_, _09647_);
  and (_09659_, _08021_, _08156_);
  not (_09660_, _09659_);
  not (_09661_, _09647_);
  or (_09662_, _09661_, _08370_);
  and (_09663_, _09662_, _09660_);
  and (_09664_, _09663_, _09658_);
  and (_09665_, _09659_, word_in[24]);
  or (_08550_, _09665_, _09664_);
  and (_09666_, _09659_, word_in[25]);
  not (_09667_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_09668_, _09650_, _09667_);
  and (_09669_, _09650_, _08513_);
  or (_09670_, _09669_, _09668_);
  or (_09671_, _09670_, _09648_);
  or (_09672_, _09655_, word_in[9]);
  and (_09673_, _09672_, _09671_);
  or (_09674_, _09673_, _09647_);
  or (_09675_, _09661_, _08511_);
  and (_09676_, _09675_, _09660_);
  and (_09677_, _09676_, _09674_);
  or (_08552_, _09677_, _09666_);
  and (_09678_, _09647_, _08525_);
  and (_09679_, _09650_, _08401_);
  not (_09680_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_09681_, _09650_, _09680_);
  or (_09682_, _09681_, _09679_);
  or (_09683_, _09682_, _09648_);
  or (_09684_, _09655_, word_in[10]);
  and (_09685_, _09684_, _09661_);
  and (_09686_, _09685_, _09683_);
  or (_09687_, _09686_, _09678_);
  and (_09688_, _09687_, _09660_);
  and (_09689_, _09659_, word_in[26]);
  or (_08556_, _09689_, _09688_);
  and (_09690_, _09647_, _08546_);
  and (_09691_, _09650_, _08415_);
  not (_09692_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_09693_, _09650_, _09692_);
  or (_09694_, _09693_, _09691_);
  or (_09695_, _09694_, _09648_);
  or (_09696_, _09655_, word_in[11]);
  and (_09697_, _09696_, _09661_);
  and (_09698_, _09697_, _09695_);
  or (_09699_, _09698_, _09690_);
  and (_09700_, _09699_, _09660_);
  and (_09701_, _09659_, word_in[27]);
  or (_08559_, _09701_, _09700_);
  and (_09702_, _09659_, word_in[28]);
  not (_09703_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_09704_, _09650_, _09703_);
  and (_09705_, _09650_, _08429_);
  or (_09706_, _09705_, _09704_);
  or (_09707_, _09706_, _09648_);
  or (_09708_, _09655_, word_in[12]);
  and (_09709_, _09708_, _09707_);
  or (_09710_, _09709_, _09647_);
  or (_09711_, _09661_, _08564_);
  and (_09712_, _09711_, _09660_);
  and (_09713_, _09712_, _09710_);
  or (_08562_, _09713_, _09702_);
  and (_09714_, _09647_, _08572_);
  and (_09715_, _09650_, _08443_);
  not (_09716_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_09717_, _09650_, _09716_);
  or (_09718_, _09717_, _09715_);
  or (_09719_, _09718_, _09648_);
  or (_09720_, _09655_, word_in[13]);
  and (_09721_, _09720_, _09661_);
  and (_09722_, _09721_, _09719_);
  or (_09723_, _09722_, _09714_);
  and (_09724_, _09723_, _09660_);
  and (_09725_, _09659_, word_in[29]);
  or (_08566_, _09725_, _09724_);
  and (_09726_, _09647_, _08593_);
  and (_09727_, _09650_, _08457_);
  not (_09728_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_09729_, _09650_, _09728_);
  or (_09730_, _09729_, _09727_);
  or (_09731_, _09730_, _09648_);
  or (_09732_, _09655_, word_in[14]);
  and (_09733_, _09732_, _09661_);
  and (_09734_, _09733_, _09731_);
  or (_09735_, _09734_, _09726_);
  and (_09736_, _09735_, _09660_);
  and (_09738_, _09659_, word_in[30]);
  or (_08568_, _09738_, _09736_);
  and (_09739_, _09659_, word_in[31]);
  nor (_09740_, _09650_, _07691_);
  and (_09741_, _09650_, _08011_);
  or (_09742_, _09741_, _09740_);
  or (_09743_, _09742_, _09648_);
  or (_09744_, _09655_, word_in[15]);
  and (_09745_, _09744_, _09743_);
  or (_09746_, _09745_, _09647_);
  or (_09747_, _09661_, _08023_);
  and (_09748_, _09747_, _09660_);
  and (_09749_, _09748_, _09746_);
  or (_08571_, _09749_, _09739_);
  and (_09750_, _07993_, _08190_);
  not (_09751_, _09750_);
  and (_09752_, _07999_, _08211_);
  not (_09753_, _09752_);
  not (_09754_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_09755_, _08352_, _08008_);
  nor (_09756_, _09755_, _09754_);
  and (_09757_, _09755_, word_in[0]);
  or (_09758_, _09757_, _09756_);
  and (_09759_, _09758_, _09753_);
  and (_09760_, _09752_, word_in[8]);
  or (_09761_, _09760_, _09759_);
  and (_09762_, _09761_, _09751_);
  not (_09763_, _07937_);
  and (_09764_, _08898_, _09763_);
  and (_09765_, _09764_, _07744_);
  and (_09766_, _09750_, word_in[16]);
  or (_09767_, _09766_, _09765_);
  or (_09768_, _09767_, _09762_);
  not (_09769_, _09765_);
  or (_09770_, _09769_, _08925_);
  and (_08636_, _09770_, _09768_);
  not (_09771_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_09772_, _09755_, _09771_);
  and (_09773_, _09755_, word_in[1]);
  or (_09774_, _09773_, _09772_);
  and (_09775_, _09774_, _09753_);
  and (_09776_, _09752_, word_in[9]);
  or (_09777_, _09776_, _09775_);
  and (_09778_, _09777_, _09751_);
  and (_09779_, _09750_, word_in[17]);
  or (_09780_, _09779_, _09765_);
  or (_09781_, _09780_, _09778_);
  or (_09782_, _09769_, _08395_);
  and (_08640_, _09782_, _09781_);
  not (_09783_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_09784_, _09755_, _09783_);
  and (_09785_, _09755_, word_in[2]);
  or (_09786_, _09785_, _09784_);
  and (_09787_, _09786_, _09753_);
  and (_09788_, _09752_, word_in[10]);
  or (_09789_, _09788_, _09787_);
  and (_09790_, _09789_, _09751_);
  and (_09791_, _09750_, word_in[18]);
  or (_09792_, _09791_, _09765_);
  or (_09793_, _09792_, _09790_);
  or (_09794_, _09769_, _08411_);
  and (_08645_, _09794_, _09793_);
  not (_09795_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_09796_, _09755_, _09795_);
  and (_09797_, _09755_, word_in[3]);
  or (_09798_, _09797_, _09796_);
  and (_09799_, _09798_, _09753_);
  and (_09800_, _09752_, word_in[11]);
  or (_09801_, _09800_, _09799_);
  and (_09802_, _09801_, _09751_);
  and (_09803_, _09750_, word_in[19]);
  or (_09804_, _09803_, _09765_);
  or (_09805_, _09804_, _09802_);
  or (_09806_, _09769_, _08425_);
  and (_08650_, _09806_, _09805_);
  not (_09807_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_09808_, _09755_, _09807_);
  and (_09809_, _09755_, word_in[4]);
  or (_09810_, _09809_, _09808_);
  and (_09811_, _09810_, _09753_);
  and (_09812_, _09752_, word_in[12]);
  or (_09813_, _09812_, _09811_);
  and (_09814_, _09813_, _09751_);
  and (_09815_, _09750_, word_in[20]);
  or (_09816_, _09815_, _09765_);
  or (_09817_, _09816_, _09814_);
  or (_09818_, _09769_, _08439_);
  and (_13433_, _09818_, _09817_);
  not (_09819_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_09820_, _09755_, _09819_);
  and (_09821_, _09755_, word_in[5]);
  or (_09822_, _09821_, _09820_);
  and (_09823_, _09822_, _09753_);
  and (_09824_, _09752_, word_in[13]);
  or (_09825_, _09824_, _09823_);
  and (_09826_, _09825_, _09751_);
  and (_09827_, _09750_, word_in[21]);
  or (_09828_, _09827_, _09765_);
  or (_09829_, _09828_, _09826_);
  or (_09830_, _09769_, _08453_);
  and (_13434_, _09830_, _09829_);
  not (_09831_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_09832_, _09755_, _09831_);
  and (_09833_, _09755_, word_in[6]);
  or (_09834_, _09833_, _09832_);
  and (_09835_, _09834_, _09753_);
  and (_09836_, _09752_, word_in[14]);
  or (_09837_, _09836_, _09835_);
  and (_09838_, _09837_, _09751_);
  and (_09839_, _09750_, word_in[22]);
  or (_09840_, _09839_, _09765_);
  or (_09841_, _09840_, _09838_);
  or (_09842_, _09769_, _08469_);
  and (_13435_, _09842_, _09841_);
  nor (_09844_, _09755_, _07820_);
  and (_09845_, _09755_, word_in[7]);
  or (_09846_, _09845_, _09844_);
  and (_09847_, _09846_, _09753_);
  and (_09848_, _09752_, word_in[15]);
  or (_09849_, _09848_, _09847_);
  and (_09850_, _09849_, _09751_);
  and (_09851_, _09750_, _08023_);
  or (_09852_, _09851_, _09765_);
  or (_09853_, _09852_, _09850_);
  or (_09854_, _09769_, _08028_);
  and (_13436_, _09854_, _09853_);
  and (_09855_, _08493_, _07813_);
  not (_09856_, _09855_);
  or (_09857_, _09856_, word_in[8]);
  and (_09858_, _08490_, _07992_);
  not (_09859_, _09858_);
  not (_09860_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_09861_, _08496_, _08008_);
  nor (_09862_, _09861_, _09860_);
  and (_09863_, _09861_, word_in[0]);
  or (_09864_, _09863_, _09862_);
  or (_09865_, _09864_, _09855_);
  and (_09866_, _09865_, _09859_);
  and (_09867_, _09866_, _09857_);
  and (_09868_, _09764_, _07775_);
  and (_09869_, _09858_, _08370_);
  or (_09870_, _09869_, _09868_);
  or (_09871_, _09870_, _09867_);
  not (_09872_, _09868_);
  or (_09873_, _09872_, word_in[24]);
  and (_13437_, _09873_, _09871_);
  and (_09874_, _09861_, word_in[1]);
  not (_09875_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_09876_, _09861_, _09875_);
  nor (_09878_, _09876_, _09874_);
  nor (_09879_, _09878_, _09855_);
  and (_09880_, _09855_, word_in[9]);
  or (_09881_, _09880_, _09879_);
  and (_09882_, _09881_, _09859_);
  and (_09883_, _09858_, _08511_);
  or (_09884_, _09883_, _09868_);
  or (_09885_, _09884_, _09882_);
  or (_09886_, _09872_, word_in[25]);
  and (_13438_, _09886_, _09885_);
  not (_09887_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_09888_, _09861_, _09887_);
  and (_09889_, _09861_, word_in[2]);
  nor (_09890_, _09889_, _09888_);
  nor (_09891_, _09890_, _09855_);
  and (_09892_, _09855_, word_in[10]);
  or (_09893_, _09892_, _09891_);
  and (_09894_, _09893_, _09859_);
  and (_09895_, _09858_, _08525_);
  or (_09896_, _09895_, _09868_);
  or (_09898_, _09896_, _09894_);
  or (_09899_, _09872_, word_in[26]);
  and (_13439_, _09899_, _09898_);
  and (_09901_, _09861_, word_in[3]);
  not (_09903_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_09904_, _09861_, _09903_);
  nor (_09906_, _09904_, _09901_);
  nor (_09907_, _09906_, _09855_);
  and (_09908_, _09855_, word_in[11]);
  or (_09909_, _09908_, _09907_);
  and (_09910_, _09909_, _09859_);
  and (_09911_, _09858_, _08546_);
  or (_09912_, _09911_, _09868_);
  or (_09913_, _09912_, _09910_);
  or (_09914_, _09872_, word_in[27]);
  and (_08744_, _09914_, _09913_);
  or (_09915_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_09916_, _06205_, _07167_);
  and (_09917_, _09916_, _05110_);
  and (_08747_, _09917_, _09915_);
  not (_09918_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_09919_, _09861_, _09918_);
  and (_09920_, _09861_, word_in[4]);
  nor (_09921_, _09920_, _09919_);
  nor (_09922_, _09921_, _09855_);
  and (_09923_, _09855_, word_in[12]);
  or (_09924_, _09923_, _09922_);
  and (_09925_, _09924_, _09859_);
  and (_09926_, _09858_, _08564_);
  or (_09927_, _09926_, _09868_);
  or (_09928_, _09927_, _09925_);
  or (_09929_, _09872_, word_in[28]);
  and (_13440_, _09929_, _09928_);
  not (_09930_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_09931_, _09861_, _09930_);
  and (_09932_, _09861_, word_in[5]);
  or (_09933_, _09932_, _09931_);
  or (_09934_, _09933_, _09855_);
  or (_09935_, _09856_, word_in[13]);
  and (_09936_, _09935_, _09934_);
  or (_09937_, _09936_, _09858_);
  or (_09938_, _09859_, _08572_);
  and (_09939_, _09938_, _09937_);
  or (_09940_, _09939_, _09868_);
  or (_09941_, _09872_, word_in[29]);
  and (_13441_, _09941_, _09940_);
  not (_09942_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_09943_, _09861_, _09942_);
  and (_09944_, _09861_, word_in[6]);
  nor (_09945_, _09944_, _09943_);
  nor (_09946_, _09945_, _09855_);
  and (_09947_, _09855_, word_in[14]);
  or (_09948_, _09947_, _09946_);
  and (_09949_, _09948_, _09859_);
  and (_09950_, _09858_, _08593_);
  or (_09951_, _09950_, _09868_);
  or (_09952_, _09951_, _09949_);
  or (_09953_, _09872_, word_in[30]);
  and (_13442_, _09953_, _09952_);
  and (_09954_, _09861_, word_in[7]);
  nor (_09955_, _09861_, _07699_);
  nor (_09956_, _09955_, _09954_);
  nor (_09957_, _09956_, _09855_);
  and (_09958_, _09855_, word_in[15]);
  or (_09959_, _09958_, _09957_);
  and (_09960_, _09959_, _09859_);
  and (_09961_, _09858_, _08023_);
  or (_09962_, _09961_, _09868_);
  or (_09963_, _09962_, _09960_);
  or (_09964_, _09872_, word_in[31]);
  and (_13443_, _09964_, _09963_);
  and (_09965_, _08642_, _07992_);
  not (_09966_, _09965_);
  and (_09967_, _08630_, _07813_);
  not (_09968_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_09969_, _08633_, _07988_);
  nor (_09970_, _09969_, _09968_);
  and (_09971_, _09969_, _08495_);
  nor (_09972_, _09971_, _09970_);
  nor (_09973_, _09972_, _09967_);
  and (_09974_, _09967_, word_in[8]);
  or (_09975_, _09974_, _09973_);
  and (_09976_, _09975_, _09966_);
  and (_09977_, _09764_, _07746_);
  and (_09978_, _09965_, _08370_);
  or (_09979_, _09978_, _09977_);
  or (_09980_, _09979_, _09976_);
  not (_09981_, _09977_);
  or (_09982_, _09981_, word_in[24]);
  and (_08823_, _09982_, _09980_);
  not (_09983_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_09984_, _09969_, _09983_);
  and (_09985_, _09969_, _08513_);
  or (_09986_, _09985_, _09984_);
  or (_09987_, _09986_, _09967_);
  not (_09988_, _09967_);
  or (_09989_, _09988_, word_in[9]);
  and (_09990_, _09989_, _09987_);
  or (_09991_, _09990_, _09965_);
  or (_09992_, _09966_, _08511_);
  and (_09993_, _09992_, _09991_);
  or (_09994_, _09993_, _09977_);
  or (_09995_, _09981_, word_in[25]);
  and (_08826_, _09995_, _09994_);
  not (_09996_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_09997_, _09969_, _09996_);
  and (_09998_, _09969_, _08401_);
  nor (_09999_, _09998_, _09997_);
  nor (_10000_, _09999_, _09967_);
  and (_10001_, _09967_, word_in[10]);
  or (_10002_, _10001_, _10000_);
  and (_10003_, _10002_, _09966_);
  and (_10004_, _09965_, _08525_);
  or (_10005_, _10004_, _09977_);
  or (_10006_, _10005_, _10003_);
  or (_10007_, _09981_, word_in[26]);
  and (_08829_, _10007_, _10006_);
  not (_10008_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_10009_, _09969_, _10008_);
  and (_10010_, _09969_, _08415_);
  nor (_10011_, _10010_, _10009_);
  nor (_10012_, _10011_, _09967_);
  and (_10013_, _09967_, word_in[11]);
  or (_10014_, _10013_, _10012_);
  and (_10015_, _10014_, _09966_);
  and (_10016_, _09965_, _08546_);
  or (_10017_, _10016_, _09977_);
  or (_10018_, _10017_, _10015_);
  or (_10019_, _09981_, word_in[27]);
  and (_08832_, _10019_, _10018_);
  or (_10020_, _09966_, _08564_);
  not (_10021_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_10022_, _09969_, _10021_);
  and (_10023_, _09969_, _08429_);
  or (_10024_, _10023_, _10022_);
  or (_10025_, _10024_, _09967_);
  or (_10026_, _09988_, word_in[12]);
  and (_10027_, _10026_, _10025_);
  or (_10028_, _10027_, _09965_);
  and (_10029_, _10028_, _10020_);
  or (_10030_, _10029_, _09977_);
  or (_10031_, _09981_, word_in[28]);
  and (_08835_, _10031_, _10030_);
  or (_10032_, _09966_, _08572_);
  not (_10033_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_10034_, _09969_, _10033_);
  and (_10035_, _09969_, _08443_);
  or (_10036_, _10035_, _10034_);
  or (_10037_, _10036_, _09967_);
  or (_10038_, _09988_, word_in[13]);
  and (_10039_, _10038_, _10037_);
  or (_10040_, _10039_, _09965_);
  and (_10041_, _10040_, _10032_);
  or (_10042_, _10041_, _09977_);
  or (_10043_, _09981_, word_in[29]);
  and (_08839_, _10043_, _10042_);
  or (_10044_, _09988_, word_in[14]);
  not (_10045_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_10046_, _09969_, _10045_);
  and (_10047_, _09969_, _08457_);
  or (_10048_, _10047_, _10046_);
  or (_10049_, _10048_, _09967_);
  and (_10050_, _10049_, _09966_);
  and (_10051_, _10050_, _10044_);
  and (_10052_, _09965_, _08593_);
  or (_10053_, _10052_, _09977_);
  or (_10054_, _10053_, _10051_);
  or (_10055_, _09981_, word_in[30]);
  and (_08843_, _10055_, _10054_);
  nor (_10056_, _09969_, _07814_);
  and (_10057_, _09969_, _08011_);
  nor (_10058_, _10057_, _10056_);
  nor (_10059_, _10058_, _09967_);
  and (_10060_, _09967_, word_in[15]);
  or (_10061_, _10060_, _10059_);
  and (_10062_, _10061_, _09966_);
  and (_10063_, _09965_, _08023_);
  or (_10064_, _10063_, _09977_);
  or (_10065_, _10064_, _10062_);
  or (_10066_, _09981_, word_in[31]);
  and (_08846_, _10066_, _10065_);
  not (_10067_, _08002_);
  or (_10068_, _10067_, word_in[8]);
  not (_10069_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_10070_, _08010_, _10069_);
  and (_10071_, _08495_, _08010_);
  or (_10072_, _10071_, _10070_);
  or (_10073_, _10072_, _08002_);
  and (_10074_, _10073_, _07998_);
  and (_10075_, _10074_, _10068_);
  and (_10076_, _08370_, _07996_);
  or (_10077_, _10076_, _08022_);
  or (_10078_, _10077_, _10075_);
  or (_10079_, _08925_, _08027_);
  and (_08906_, _10079_, _10078_);
  or (_10080_, _10067_, word_in[9]);
  not (_10081_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_10082_, _08010_, _10081_);
  and (_10083_, _08513_, _08010_);
  or (_10084_, _10083_, _10082_);
  or (_10085_, _10084_, _08002_);
  and (_10086_, _10085_, _07998_);
  and (_10087_, _10086_, _10080_);
  and (_10088_, _08511_, _07996_);
  or (_10089_, _10088_, _08022_);
  or (_10090_, _10089_, _10087_);
  or (_10091_, _08395_, _08027_);
  and (_08909_, _10091_, _10090_);
  not (_10092_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_10093_, _08010_, _10092_);
  and (_10094_, _08401_, _08010_);
  or (_10095_, _10094_, _10093_);
  or (_10096_, _10095_, _08002_);
  or (_10097_, _10067_, word_in[10]);
  and (_10098_, _10097_, _10096_);
  or (_10099_, _10098_, _07996_);
  or (_10100_, _08525_, _07998_);
  and (_10101_, _10100_, _10099_);
  or (_10102_, _10101_, _08022_);
  or (_10103_, _08411_, _08027_);
  and (_08913_, _10103_, _10102_);
  not (_10105_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_10106_, _08010_, _10105_);
  and (_10107_, _08415_, _08010_);
  nor (_10108_, _10107_, _10106_);
  nor (_10109_, _10108_, _08002_);
  and (_10110_, _08002_, word_in[11]);
  or (_10111_, _10110_, _10109_);
  and (_10112_, _10111_, _07998_);
  and (_10113_, _08546_, _07996_);
  or (_10114_, _10113_, _08022_);
  or (_10115_, _10114_, _10112_);
  or (_10116_, _08425_, _08027_);
  and (_08916_, _10116_, _10115_);
  or (_10117_, _10067_, word_in[12]);
  not (_10118_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_10119_, _08010_, _10118_);
  and (_10120_, _08429_, _08010_);
  or (_10121_, _10120_, _10119_);
  or (_10122_, _10121_, _08002_);
  and (_10123_, _10122_, _07998_);
  and (_10124_, _10123_, _10117_);
  and (_10125_, _08564_, _07996_);
  or (_10126_, _10125_, _08022_);
  or (_10127_, _10126_, _10124_);
  or (_10128_, _08439_, _08027_);
  and (_08920_, _10128_, _10127_);
  and (_10129_, _08572_, _07996_);
  and (_10130_, _08443_, _08010_);
  not (_10131_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_10132_, _08010_, _10131_);
  nor (_10133_, _10132_, _10130_);
  nor (_10134_, _10133_, _08002_);
  and (_10135_, _08002_, word_in[13]);
  or (_10136_, _10135_, _10134_);
  and (_10137_, _10136_, _07998_);
  or (_10138_, _10137_, _10129_);
  and (_10139_, _10138_, _08027_);
  and (_10140_, _08453_, _08022_);
  or (_08923_, _10140_, _10139_);
  or (_10141_, _10067_, word_in[14]);
  not (_10142_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_10143_, _08010_, _10142_);
  and (_10145_, _08457_, _08010_);
  or (_10146_, _10145_, _10143_);
  or (_10147_, _10146_, _08002_);
  and (_10148_, _10147_, _07998_);
  and (_10149_, _10148_, _10141_);
  and (_10150_, _08593_, _07996_);
  or (_10151_, _10150_, _08022_);
  or (_10152_, _10151_, _10149_);
  or (_10153_, _08469_, _08027_);
  and (_08926_, _10153_, _10152_);
  nor (_09231_, _05845_, rst);
  and (_10154_, _06624_, _05419_);
  nor (_10155_, _05447_, _06121_);
  and (_10156_, _10155_, _05794_);
  and (_10157_, _10156_, _10154_);
  and (_10158_, _10157_, _08272_);
  or (_10159_, _10158_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_10160_, _05806_, _05992_);
  and (_10161_, _10160_, _06618_);
  and (_10162_, _10161_, _05434_);
  not (_10163_, _10162_);
  and (_10164_, _10163_, _10159_);
  nand (_10165_, _10158_, _05872_);
  and (_10166_, _10165_, _10164_);
  nor (_10167_, _10163_, _05938_);
  or (_10168_, _10167_, _10166_);
  and (_09234_, _10168_, _05110_);
  nor (_10169_, _06173_, _05785_);
  not (_10170_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_10171_, _05376_, _10170_);
  nor (_10172_, _10171_, _10169_);
  or (_10173_, _10172_, _06632_);
  and (_10174_, _10173_, _10157_);
  and (_10175_, _10160_, _05434_);
  and (_10176_, _10175_, _06618_);
  and (_10177_, _10176_, _06194_);
  nor (_10178_, _05376_, _05485_);
  nand (_10179_, _10178_, _10157_);
  nor (_10180_, _10176_, _10170_);
  and (_10181_, _10180_, _10179_);
  or (_10182_, _10181_, _10177_);
  or (_10183_, _10182_, _10174_);
  and (_09629_, _10183_, _05110_);
  and (_10184_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_10185_, _10184_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_10186_, _05711_, _05650_);
  and (_10187_, _05575_, _05489_);
  nand (_10188_, _05158_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_10189_, _10188_, _10184_);
  or (_10190_, _10189_, _10187_);
  or (_10191_, _10190_, _10186_);
  and (_10192_, _10191_, _10185_);
  or (_10193_, _10192_, _10157_);
  or (_10194_, _05488_, _06646_);
  nand (_10195_, _10194_, _10157_);
  or (_10196_, _10195_, _05784_);
  and (_10197_, _10196_, _10193_);
  or (_10198_, _10197_, _10162_);
  nand (_10199_, _10162_, _05841_);
  and (_10200_, _10199_, _05110_);
  and (_09633_, _10200_, _10198_);
  and (_10201_, _10157_, _08133_);
  or (_10202_, _10201_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_10203_, _10202_, _10163_);
  nand (_10204_, _10201_, _05872_);
  and (_10205_, _10204_, _10203_);
  nor (_10206_, _10163_, _06054_);
  or (_10207_, _10206_, _10205_);
  and (_09636_, _10207_, _05110_);
  and (_10208_, _05376_, _05485_);
  and (_10209_, _10208_, _05782_);
  and (_10210_, _10209_, _10157_);
  not (_10211_, _10157_);
  nor (_10212_, _10178_, _10208_);
  or (_10213_, _10212_, _10211_);
  and (_10214_, _10213_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  not (_10215_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_10216_, _10179_, _10215_);
  or (_10217_, _10216_, _10214_);
  or (_10218_, _10217_, _10210_);
  and (_10219_, _10218_, _10163_);
  nor (_10220_, _10163_, _05334_);
  or (_10221_, _10220_, _10219_);
  and (_09639_, _10221_, _05110_);
  or (_10222_, _06384_, _07153_);
  or (_10223_, _05473_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_10224_, _10223_, _05110_);
  and (_09737_, _10224_, _10222_);
  and (_10225_, _07742_, word_in[0]);
  nand (_10226_, _07603_, _09436_);
  or (_10227_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_10228_, _10227_, _10226_);
  and (_10229_, _10228_, _07624_);
  nand (_10230_, _07603_, _09649_);
  or (_10231_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_10232_, _10231_, _10230_);
  and (_10233_, _10232_, _07636_);
  nand (_10234_, _07603_, _09860_);
  or (_10235_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_10236_, _10235_, _10234_);
  and (_10237_, _10236_, _07633_);
  or (_10238_, _10237_, _10233_);
  or (_10239_, _10238_, _10229_);
  nand (_10240_, _07603_, _10069_);
  or (_10241_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_10242_, _10241_, _10240_);
  and (_10243_, _10242_, _07644_);
  or (_10244_, _10243_, _07659_);
  or (_10245_, _10244_, _10239_);
  nand (_10246_, _07603_, _08499_);
  or (_10247_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_10248_, _10247_, _10246_);
  and (_10249_, _10248_, _07624_);
  nand (_10250_, _07603_, _08765_);
  or (_10251_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_10252_, _10251_, _10250_);
  and (_10253_, _10252_, _07636_);
  nand (_10254_, _07603_, _09021_);
  or (_10255_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_10257_, _10255_, _10254_);
  and (_10258_, _10257_, _07633_);
  or (_10259_, _10258_, _10253_);
  or (_10260_, _10259_, _10249_);
  nand (_10261_, _07603_, _09222_);
  or (_10262_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_10263_, _10262_, _10261_);
  and (_10264_, _10263_, _07644_);
  or (_10265_, _10264_, _07612_);
  or (_10266_, _10265_, _10260_);
  and (_10267_, _10266_, _10245_);
  and (_10268_, _10267_, _07683_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _10268_, _10225_);
  nor (_10269_, _07683_, _08379_);
  nand (_10270_, _07603_, _09456_);
  or (_10271_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_10272_, _10271_, _10270_);
  and (_10273_, _10272_, _07624_);
  nand (_10274_, _07603_, _09875_);
  or (_10275_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_10276_, _10275_, _10274_);
  and (_10277_, _10276_, _07633_);
  nand (_10278_, _07603_, _09667_);
  or (_10279_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_10280_, _10279_, _10278_);
  and (_10281_, _10280_, _07636_);
  or (_10282_, _10281_, _10277_);
  or (_10283_, _10282_, _10273_);
  nand (_10284_, _07603_, _10081_);
  or (_10285_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_10286_, _10285_, _10284_);
  and (_10287_, _10286_, _07644_);
  or (_10288_, _10287_, _07659_);
  or (_10289_, _10288_, _10283_);
  nand (_10290_, _07603_, _08515_);
  or (_10291_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_10292_, _10291_, _10290_);
  and (_10293_, _10292_, _07624_);
  nand (_10294_, _07603_, _08779_);
  or (_10295_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_10296_, _10295_, _10294_);
  and (_10297_, _10296_, _07636_);
  nand (_10298_, _07603_, _09035_);
  or (_10299_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_10300_, _10299_, _10298_);
  and (_10301_, _10300_, _07633_);
  or (_10302_, _10301_, _10297_);
  or (_10303_, _10302_, _10293_);
  nand (_10304_, _07603_, _09239_);
  or (_10305_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_10307_, _10305_, _10304_);
  and (_10308_, _10307_, _07644_);
  or (_10309_, _10308_, _07612_);
  or (_10310_, _10309_, _10303_);
  and (_10311_, _10310_, _10289_);
  and (_10312_, _10311_, _07683_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _10312_, _10269_);
  and (_10313_, _07742_, word_in[2]);
  nand (_10314_, _07603_, _09471_);
  or (_10315_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_10316_, _10315_, _10314_);
  and (_10317_, _10316_, _07624_);
  nand (_10318_, _07603_, _09680_);
  or (_10319_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_10320_, _10319_, _10318_);
  and (_10321_, _10320_, _07636_);
  nand (_10322_, _07603_, _09887_);
  or (_10323_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_10324_, _10323_, _10322_);
  and (_10325_, _10324_, _07633_);
  or (_10326_, _10325_, _10321_);
  or (_10327_, _10326_, _10317_);
  nand (_10328_, _07603_, _10092_);
  or (_10329_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_10330_, _10329_, _10328_);
  and (_10331_, _10330_, _07644_);
  or (_10332_, _10331_, _07659_);
  or (_10333_, _10332_, _10327_);
  nand (_10334_, _07603_, _08528_);
  or (_10335_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_10336_, _10335_, _10334_);
  and (_10337_, _10336_, _07624_);
  nand (_10338_, _07603_, _08791_);
  or (_10339_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_10340_, _10339_, _10338_);
  and (_10341_, _10340_, _07636_);
  nand (_10342_, _07603_, _09048_);
  or (_10343_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_10344_, _10343_, _10342_);
  and (_10345_, _10344_, _07633_);
  or (_10346_, _10345_, _10341_);
  or (_10347_, _10346_, _10337_);
  nand (_10348_, _07603_, _09252_);
  or (_10349_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_10350_, _10349_, _10348_);
  and (_10351_, _10350_, _07644_);
  or (_10352_, _10351_, _07612_);
  or (_10353_, _10352_, _10347_);
  and (_10354_, _10353_, _10333_);
  and (_10355_, _10354_, _07683_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _10355_, _10313_);
  and (_10356_, _07742_, word_in[3]);
  nand (_10357_, _07603_, _09482_);
  or (_10358_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_10359_, _10358_, _10357_);
  and (_10360_, _10359_, _07624_);
  nand (_10361_, _07603_, _09692_);
  or (_10362_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_10363_, _10362_, _10361_);
  and (_10364_, _10363_, _07636_);
  nand (_10365_, _07603_, _09903_);
  or (_10366_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_10367_, _10366_, _10365_);
  and (_10368_, _10367_, _07633_);
  or (_10369_, _10368_, _10364_);
  or (_10370_, _10369_, _10360_);
  nand (_10371_, _07603_, _10105_);
  or (_10372_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_10373_, _10372_, _10371_);
  and (_10374_, _10373_, _07644_);
  or (_10375_, _10374_, _07659_);
  or (_10376_, _10375_, _10370_);
  nand (_10377_, _07603_, _08538_);
  or (_10378_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_10379_, _10378_, _10377_);
  and (_10380_, _10379_, _07624_);
  nand (_10381_, _07603_, _08803_);
  or (_10382_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_10383_, _10382_, _10381_);
  and (_10384_, _10383_, _07636_);
  nand (_10386_, _07603_, _09059_);
  or (_10387_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_10388_, _10387_, _10386_);
  and (_10389_, _10388_, _07633_);
  or (_10390_, _10389_, _10384_);
  or (_10391_, _10390_, _10380_);
  nand (_10392_, _07603_, _09264_);
  or (_10393_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_10394_, _10393_, _10392_);
  and (_10395_, _10394_, _07644_);
  or (_10396_, _10395_, _07612_);
  or (_10397_, _10396_, _10391_);
  and (_10398_, _10397_, _10376_);
  and (_10399_, _10398_, _07683_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _10399_, _10356_);
  and (_10401_, _07742_, word_in[4]);
  nand (_10402_, _07603_, _09494_);
  or (_10403_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_10404_, _10403_, _10402_);
  and (_10405_, _10404_, _07624_);
  nand (_10407_, _07603_, _09703_);
  or (_10408_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_10409_, _10408_, _10407_);
  and (_10410_, _10409_, _07636_);
  nand (_10411_, _07603_, _09918_);
  or (_10412_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_10413_, _10412_, _10411_);
  and (_10414_, _10413_, _07633_);
  or (_10415_, _10414_, _10410_);
  or (_10416_, _10415_, _10405_);
  nand (_10417_, _07603_, _10118_);
  or (_10418_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_10419_, _10418_, _10417_);
  and (_10420_, _10419_, _07644_);
  or (_10421_, _10420_, _07659_);
  or (_10422_, _10421_, _10416_);
  nand (_10423_, _07603_, _08553_);
  or (_10424_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_10425_, _10424_, _10423_);
  and (_10426_, _10425_, _07624_);
  nand (_10428_, _07603_, _08815_);
  or (_10429_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_10430_, _10429_, _10428_);
  and (_10431_, _10430_, _07636_);
  nand (_10432_, _07603_, _09071_);
  or (_10433_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_10434_, _10433_, _10432_);
  and (_10435_, _10434_, _07633_);
  or (_10436_, _10435_, _10431_);
  or (_10437_, _10436_, _10426_);
  nand (_10438_, _07603_, _09276_);
  or (_10439_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_10440_, _10439_, _10438_);
  and (_10441_, _10440_, _07644_);
  or (_10442_, _10441_, _07612_);
  or (_10443_, _10442_, _10437_);
  and (_10444_, _10443_, _10422_);
  and (_10445_, _10444_, _07683_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _10445_, _10401_);
  and (_10446_, _07742_, word_in[5]);
  nand (_10447_, _07603_, _09506_);
  or (_10448_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_10449_, _10448_, _10447_);
  and (_10450_, _10449_, _07624_);
  nand (_10451_, _07603_, _09930_);
  or (_10452_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_10453_, _10452_, _10451_);
  and (_10454_, _10453_, _07633_);
  nand (_10455_, _07603_, _09716_);
  or (_10456_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_10457_, _10456_, _10455_);
  and (_10458_, _10457_, _07636_);
  or (_10459_, _10458_, _10454_);
  or (_10461_, _10459_, _10450_);
  nand (_10462_, _07603_, _10131_);
  or (_10463_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_10464_, _10463_, _10462_);
  and (_10465_, _10464_, _07644_);
  or (_10466_, _10465_, _07659_);
  or (_10467_, _10466_, _10461_);
  nand (_10468_, _07603_, _08575_);
  or (_10469_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_10470_, _10469_, _10468_);
  and (_10471_, _10470_, _07624_);
  nand (_10473_, _07603_, _08830_);
  or (_10474_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_10475_, _10474_, _10473_);
  and (_10476_, _10475_, _07636_);
  nand (_10477_, _07603_, _09082_);
  or (_10478_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_10479_, _10478_, _10477_);
  and (_10480_, _10479_, _07633_);
  or (_10481_, _10480_, _10476_);
  or (_10482_, _10481_, _10471_);
  nand (_10483_, _07603_, _09288_);
  or (_10484_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_10485_, _10484_, _10483_);
  and (_10486_, _10485_, _07644_);
  or (_10487_, _10486_, _07612_);
  or (_10488_, _10487_, _10482_);
  and (_10489_, _10488_, _10467_);
  and (_10490_, _10489_, _07683_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _10490_, _10446_);
  and (_10491_, _07742_, word_in[6]);
  nand (_10492_, _07603_, _09518_);
  or (_10493_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_10494_, _10493_, _10492_);
  and (_10495_, _10494_, _07624_);
  nand (_10496_, _07603_, _09942_);
  or (_10497_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_10498_, _10497_, _10496_);
  and (_10499_, _10498_, _07633_);
  nand (_10500_, _07603_, _09728_);
  or (_10501_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_10502_, _10501_, _10500_);
  and (_10503_, _10502_, _07636_);
  or (_10504_, _10503_, _10499_);
  or (_10505_, _10504_, _10495_);
  nand (_10506_, _07603_, _10142_);
  or (_10507_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_10508_, _10507_, _10506_);
  and (_10509_, _10508_, _07644_);
  or (_10510_, _10509_, _07659_);
  or (_10511_, _10510_, _10505_);
  nand (_10512_, _07603_, _08585_);
  or (_10513_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_10514_, _10513_, _10512_);
  and (_10515_, _10514_, _07624_);
  nand (_10516_, _07603_, _08847_);
  or (_10518_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_10519_, _10518_, _10516_);
  and (_10520_, _10519_, _07636_);
  nand (_10521_, _07603_, _09095_);
  or (_10522_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_10523_, _10522_, _10521_);
  and (_10525_, _10523_, _07633_);
  or (_10526_, _10525_, _10520_);
  or (_10527_, _10526_, _10515_);
  nand (_10528_, _07603_, _09300_);
  or (_10529_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_10530_, _10529_, _10528_);
  and (_10531_, _10530_, _07644_);
  or (_10532_, _10531_, _07612_);
  or (_10533_, _10532_, _10527_);
  and (_10534_, _10533_, _10511_);
  and (_10535_, _10534_, _07683_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _10535_, _10491_);
  and (_10536_, _07793_, word_in[8]);
  nand (_10537_, _07603_, _09543_);
  or (_10538_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_10540_, _10538_, _10537_);
  and (_10541_, _10540_, _07796_);
  nand (_10542_, _07603_, _09335_);
  or (_10543_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_10544_, _10543_, _10542_);
  and (_10545_, _10544_, _07794_);
  or (_10546_, _10545_, _10541_);
  and (_10547_, _10546_, _07757_);
  nand (_10548_, _07603_, _08637_);
  or (_10549_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_10550_, _10549_, _10548_);
  and (_10551_, _10550_, _07796_);
  nand (_10552_, _07603_, _08350_);
  or (_10553_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_10554_, _10553_, _10552_);
  and (_10555_, _10554_, _07794_);
  or (_10556_, _10555_, _10551_);
  and (_10557_, _10556_, _07760_);
  nand (_10559_, _07603_, _09118_);
  or (_10560_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_10561_, _10560_, _10559_);
  and (_10563_, _10561_, _07796_);
  nand (_10564_, _07603_, _08907_);
  or (_10565_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_10566_, _10565_, _10564_);
  and (_10568_, _10566_, _07794_);
  or (_10569_, _10568_, _10563_);
  and (_10570_, _10569_, _07841_);
  or (_10571_, _10570_, _10557_);
  nand (_10572_, _07603_, _09968_);
  or (_10573_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_10574_, _10573_, _10572_);
  and (_10575_, _10574_, _07796_);
  nand (_10576_, _07603_, _09754_);
  or (_10577_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_10578_, _10577_, _10576_);
  and (_10579_, _10578_, _07794_);
  or (_10580_, _10579_, _10575_);
  and (_10581_, _10580_, _07813_);
  or (_10583_, _10581_, _10571_);
  nor (_10584_, _10583_, _10547_);
  nor (_10586_, _10584_, _07793_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _10586_, _10536_);
  and (_10588_, _07793_, word_in[9]);
  nand (_10589_, _07603_, _09559_);
  or (_10590_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_10591_, _10590_, _10589_);
  and (_10592_, _10591_, _07796_);
  nand (_10593_, _07603_, _09351_);
  or (_10594_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_10595_, _10594_, _10593_);
  and (_10596_, _10595_, _07794_);
  or (_10598_, _10596_, _10592_);
  and (_10599_, _10598_, _07757_);
  nand (_10601_, _07603_, _08659_);
  or (_10602_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_10603_, _10602_, _10601_);
  and (_10604_, _10603_, _07796_);
  and (_10605_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_10606_, _07603_, _08515_);
  or (_10607_, _10606_, _10605_);
  and (_10608_, _10607_, _07794_);
  or (_10609_, _10608_, _10604_);
  and (_10610_, _10609_, _07760_);
  nand (_10611_, _07603_, _09136_);
  or (_10612_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_10613_, _10612_, _10611_);
  and (_10614_, _10613_, _07796_);
  nand (_10615_, _07603_, _08929_);
  or (_10616_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_10617_, _10616_, _10615_);
  and (_10618_, _10617_, _07794_);
  or (_10619_, _10618_, _10614_);
  and (_10621_, _10619_, _07841_);
  or (_10622_, _10621_, _10610_);
  nand (_10623_, _07603_, _09983_);
  or (_10624_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_10625_, _10624_, _10623_);
  and (_10626_, _10625_, _07796_);
  nand (_10627_, _07603_, _09771_);
  or (_10628_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_10629_, _10628_, _10627_);
  and (_10630_, _10629_, _07794_);
  or (_10631_, _10630_, _10626_);
  and (_10632_, _10631_, _07813_);
  or (_10633_, _10632_, _10622_);
  nor (_10634_, _10633_, _10599_);
  nor (_10635_, _10634_, _07793_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _10635_, _10588_);
  and (_10636_, _07793_, word_in[10]);
  nand (_10637_, _07603_, _09572_);
  or (_10638_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_10639_, _10638_, _10637_);
  and (_10640_, _10639_, _07796_);
  nand (_10642_, _07603_, _09363_);
  or (_10643_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_10644_, _10643_, _10642_);
  and (_10646_, _10644_, _07794_);
  or (_10647_, _10646_, _10640_);
  and (_10648_, _10647_, _07757_);
  nand (_10650_, _07603_, _08671_);
  or (_10651_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_10652_, _10651_, _10650_);
  and (_10653_, _10652_, _07796_);
  nand (_10655_, _07603_, _08398_);
  or (_10656_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_10657_, _10656_, _10655_);
  and (_10658_, _10657_, _07794_);
  or (_10659_, _10658_, _10653_);
  and (_10661_, _10659_, _07760_);
  nand (_10662_, _07603_, _09148_);
  or (_10664_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_10665_, _10664_, _10662_);
  and (_10666_, _10665_, _07796_);
  nand (_10667_, _07603_, _08941_);
  or (_10668_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_10669_, _10668_, _10667_);
  and (_10670_, _10669_, _07794_);
  or (_10671_, _10670_, _10666_);
  and (_10672_, _10671_, _07841_);
  or (_10673_, _10672_, _10661_);
  nand (_10674_, _07603_, _09996_);
  or (_10675_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_10676_, _10675_, _10674_);
  and (_10677_, _10676_, _07796_);
  nand (_10678_, _07603_, _09783_);
  or (_10680_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_10681_, _10680_, _10678_);
  and (_10682_, _10681_, _07794_);
  or (_10683_, _10682_, _10677_);
  and (_10685_, _10683_, _07813_);
  or (_10686_, _10685_, _10673_);
  nor (_10687_, _10686_, _10648_);
  nor (_10688_, _10687_, _07793_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _10688_, _10636_);
  and (_10689_, _07793_, word_in[11]);
  nand (_10690_, _07603_, _09585_);
  or (_10691_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_10692_, _10691_, _10690_);
  and (_10693_, _10692_, _07796_);
  nand (_10694_, _07603_, _09375_);
  or (_10695_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_10696_, _10695_, _10694_);
  and (_10698_, _10696_, _07794_);
  or (_10699_, _10698_, _10693_);
  and (_10700_, _10699_, _07757_);
  nand (_10701_, _07603_, _10008_);
  or (_10702_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_10703_, _10702_, _10701_);
  and (_10704_, _10703_, _07796_);
  nand (_10706_, _07603_, _09795_);
  or (_10707_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_10708_, _10707_, _10706_);
  and (_10710_, _10708_, _07794_);
  or (_10711_, _10710_, _10704_);
  and (_10713_, _10711_, _07813_);
  nand (_10715_, _07603_, _09160_);
  or (_10716_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_10718_, _10716_, _10715_);
  and (_10719_, _10718_, _07796_);
  nand (_10721_, _07603_, _08953_);
  or (_10722_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_10723_, _10722_, _10721_);
  and (_10725_, _10723_, _07794_);
  or (_10726_, _10725_, _10719_);
  and (_10727_, _10726_, _07841_);
  nand (_10728_, _07603_, _08683_);
  or (_10729_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_10731_, _10729_, _10728_);
  and (_10732_, _10731_, _07796_);
  nand (_10733_, _07603_, _08413_);
  or (_10734_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_10735_, _10734_, _10733_);
  and (_10737_, _10735_, _07794_);
  or (_10738_, _10737_, _10732_);
  and (_10740_, _10738_, _07760_);
  or (_10741_, _10740_, _10727_);
  or (_10742_, _10741_, _10713_);
  nor (_10743_, _10742_, _10700_);
  nor (_10744_, _10743_, _07793_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _10744_, _10689_);
  and (_10745_, _07793_, word_in[12]);
  nand (_10747_, _07603_, _09598_);
  or (_10748_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_10749_, _10748_, _10747_);
  and (_10750_, _10749_, _07796_);
  nand (_10751_, _07603_, _09387_);
  or (_10752_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_10753_, _10752_, _10751_);
  and (_10754_, _10753_, _07794_);
  or (_10756_, _10754_, _10750_);
  and (_10757_, _10756_, _07757_);
  nand (_10758_, _07603_, _08696_);
  or (_10759_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_10760_, _10759_, _10758_);
  and (_10761_, _10760_, _07796_);
  nand (_10762_, _07603_, _08427_);
  or (_10763_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_10764_, _10763_, _10762_);
  and (_10765_, _10764_, _07794_);
  or (_10766_, _10765_, _10761_);
  and (_10767_, _10766_, _07760_);
  nand (_10768_, _07603_, _09172_);
  or (_10769_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_10770_, _10769_, _10768_);
  and (_10771_, _10770_, _07796_);
  nand (_10772_, _07603_, _08965_);
  or (_10773_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_10774_, _10773_, _10772_);
  and (_10775_, _10774_, _07794_);
  or (_10776_, _10775_, _10771_);
  and (_10777_, _10776_, _07841_);
  or (_10778_, _10777_, _10767_);
  nand (_10779_, _07603_, _10021_);
  or (_10780_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_10781_, _10780_, _10779_);
  and (_10782_, _10781_, _07796_);
  nand (_10783_, _07603_, _09807_);
  or (_10785_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_10786_, _10785_, _10783_);
  and (_10787_, _10786_, _07794_);
  or (_10788_, _10787_, _10782_);
  and (_10790_, _10788_, _07813_);
  or (_10791_, _10790_, _10778_);
  nor (_10792_, _10791_, _10757_);
  nor (_10793_, _10792_, _07793_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _10793_, _10745_);
  and (_10794_, _07793_, word_in[13]);
  nand (_10795_, _07603_, _09608_);
  or (_10796_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_10797_, _10796_, _10795_);
  and (_10798_, _10797_, _07796_);
  nand (_10799_, _07603_, _09399_);
  or (_10800_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_10801_, _10800_, _10799_);
  and (_10802_, _10801_, _07794_);
  or (_10804_, _10802_, _10798_);
  and (_10805_, _10804_, _07757_);
  nand (_10806_, _07603_, _08708_);
  or (_10807_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_10808_, _10807_, _10806_);
  and (_10809_, _10808_, _07796_);
  nand (_10810_, _07603_, _08441_);
  or (_10811_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_10812_, _10811_, _10810_);
  and (_10814_, _10812_, _07794_);
  or (_10815_, _10814_, _10809_);
  and (_10816_, _10815_, _07760_);
  nand (_10817_, _07603_, _09184_);
  or (_10818_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_10819_, _10818_, _10817_);
  and (_10820_, _10819_, _07796_);
  nand (_10821_, _07603_, _08977_);
  or (_10822_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_10823_, _10822_, _10821_);
  and (_10824_, _10823_, _07794_);
  or (_10825_, _10824_, _10820_);
  and (_10826_, _10825_, _07841_);
  or (_10827_, _10826_, _10816_);
  nand (_10828_, _07603_, _10033_);
  or (_10829_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_10830_, _10829_, _10828_);
  and (_10831_, _10830_, _07796_);
  nand (_10832_, _07603_, _09819_);
  or (_10833_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_10834_, _10833_, _10832_);
  and (_10835_, _10834_, _07794_);
  or (_10836_, _10835_, _10831_);
  and (_10837_, _10836_, _07813_);
  or (_10838_, _10837_, _10827_);
  nor (_10839_, _10838_, _10805_);
  nor (_10840_, _10839_, _07793_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _10840_, _10794_);
  and (_10841_, _07793_, word_in[14]);
  nand (_10842_, _07603_, _09621_);
  or (_10843_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_10844_, _10843_, _10842_);
  and (_10845_, _10844_, _07796_);
  nand (_10846_, _07603_, _09411_);
  or (_10847_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_10848_, _10847_, _10846_);
  and (_10849_, _10848_, _07794_);
  or (_10850_, _10849_, _10845_);
  and (_10851_, _10850_, _07757_);
  nand (_10852_, _07603_, _10045_);
  or (_10853_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_10854_, _10853_, _10852_);
  and (_10855_, _10854_, _07796_);
  nand (_10856_, _07603_, _09831_);
  or (_10857_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_10858_, _10857_, _10856_);
  and (_10859_, _10858_, _07794_);
  or (_10860_, _10859_, _10855_);
  and (_10861_, _10860_, _07813_);
  nand (_10863_, _07603_, _09197_);
  or (_10864_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_10865_, _10864_, _10863_);
  and (_10866_, _10865_, _07796_);
  nand (_10867_, _07603_, _08990_);
  or (_10868_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_10869_, _10868_, _10867_);
  and (_10870_, _10869_, _07794_);
  or (_10871_, _10870_, _10866_);
  and (_10872_, _10871_, _07841_);
  nand (_10873_, _07603_, _08718_);
  or (_10874_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_10875_, _10874_, _10873_);
  and (_10876_, _10875_, _07796_);
  nand (_10877_, _07603_, _08455_);
  or (_10878_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_10879_, _10878_, _10877_);
  and (_10881_, _10879_, _07794_);
  or (_10882_, _10881_, _10876_);
  and (_10884_, _10882_, _07760_);
  or (_10885_, _10884_, _10872_);
  or (_10886_, _10885_, _10861_);
  nor (_10887_, _10886_, _10851_);
  nor (_10888_, _10887_, _07793_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _10888_, _10841_);
  and (_10889_, _07896_, word_in[16]);
  and (_10890_, _10232_, _07624_);
  and (_10891_, _10236_, _07636_);
  or (_10892_, _10891_, _10890_);
  and (_10893_, _10242_, _07633_);
  and (_10894_, _10228_, _07644_);
  or (_10895_, _10894_, _10893_);
  or (_10896_, _10895_, _10892_);
  or (_10897_, _10896_, _07907_);
  and (_10898_, _10257_, _07636_);
  and (_10899_, _10248_, _07644_);
  or (_10900_, _10899_, _10898_);
  and (_10901_, _10263_, _07633_);
  and (_10902_, _10252_, _07624_);
  or (_10903_, _10902_, _10901_);
  or (_10904_, _10903_, _10900_);
  or (_10905_, _10904_, _07863_);
  nand (_10906_, _10905_, _10897_);
  nor (_10907_, _10906_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _10907_, _10889_);
  and (_10908_, _07896_, word_in[17]);
  and (_10909_, _10286_, _07633_);
  and (_10910_, _10280_, _07624_);
  or (_10911_, _10910_, _10909_);
  and (_10912_, _10276_, _07636_);
  and (_10913_, _10272_, _07644_);
  or (_10914_, _10913_, _10912_);
  or (_10915_, _10914_, _10911_);
  or (_10916_, _10915_, _07907_);
  and (_10917_, _10307_, _07633_);
  and (_10918_, _10300_, _07636_);
  or (_10919_, _10918_, _10917_);
  and (_10920_, _10296_, _07624_);
  and (_10921_, _10292_, _07644_);
  or (_10922_, _10921_, _10920_);
  or (_10923_, _10922_, _10919_);
  or (_10924_, _10923_, _07863_);
  nand (_10925_, _10924_, _10916_);
  nor (_10926_, _10925_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _10926_, _10908_);
  and (_10927_, _07896_, word_in[18]);
  and (_10928_, _10350_, _07633_);
  and (_10929_, _10340_, _07624_);
  or (_10930_, _10929_, _10928_);
  and (_10931_, _10344_, _07636_);
  and (_10932_, _10336_, _07644_);
  or (_10933_, _10932_, _10931_);
  or (_10934_, _10933_, _10930_);
  or (_10936_, _10934_, _07863_);
  and (_10937_, _10320_, _07624_);
  and (_10938_, _10324_, _07636_);
  or (_10939_, _10938_, _10937_);
  and (_10940_, _10330_, _07633_);
  and (_10941_, _10316_, _07644_);
  or (_10943_, _10941_, _10940_);
  or (_10944_, _10943_, _10939_);
  or (_10945_, _10944_, _07907_);
  nand (_10946_, _10945_, _10936_);
  nor (_10947_, _10946_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _10947_, _10927_);
  and (_10948_, _07896_, word_in[19]);
  and (_10949_, _10363_, _07624_);
  and (_10950_, _10367_, _07636_);
  or (_10951_, _10950_, _10949_);
  and (_10952_, _10373_, _07633_);
  and (_10953_, _10359_, _07644_);
  or (_10954_, _10953_, _10952_);
  or (_10955_, _10954_, _10951_);
  or (_10956_, _10955_, _07907_);
  and (_10957_, _10388_, _07636_);
  and (_10958_, _10379_, _07644_);
  or (_10959_, _10958_, _10957_);
  and (_10960_, _10394_, _07633_);
  and (_10961_, _10383_, _07624_);
  or (_10962_, _10961_, _10960_);
  or (_10963_, _10962_, _10959_);
  or (_10964_, _10963_, _07863_);
  nand (_10965_, _10964_, _10956_);
  nor (_10967_, _10965_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _10967_, _10948_);
  and (_10968_, _07896_, word_in[20]);
  and (_10969_, _10430_, _07624_);
  and (_10970_, _10425_, _07644_);
  or (_10971_, _10970_, _10969_);
  and (_10972_, _10440_, _07633_);
  and (_10973_, _10434_, _07636_);
  or (_10975_, _10973_, _10972_);
  or (_10976_, _10975_, _10971_);
  or (_10977_, _10976_, _07863_);
  and (_10978_, _10409_, _07624_);
  and (_10980_, _10404_, _07644_);
  or (_10981_, _10980_, _10978_);
  and (_10982_, _10419_, _07633_);
  and (_10983_, _10413_, _07636_);
  or (_10984_, _10983_, _10982_);
  or (_10986_, _10984_, _10981_);
  or (_10987_, _10986_, _07907_);
  nand (_10988_, _10987_, _10977_);
  nor (_10989_, _10988_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _10989_, _10968_);
  and (_10990_, _07896_, word_in[21]);
  and (_10991_, _10475_, _07624_);
  and (_10992_, _10470_, _07644_);
  or (_10993_, _10992_, _10991_);
  and (_10994_, _10485_, _07633_);
  and (_10995_, _10479_, _07636_);
  or (_10996_, _10995_, _10994_);
  or (_10997_, _10996_, _10993_);
  or (_10998_, _10997_, _07863_);
  and (_10999_, _10464_, _07633_);
  and (_11000_, _10457_, _07624_);
  or (_11001_, _11000_, _10999_);
  and (_11002_, _10453_, _07636_);
  and (_11003_, _10449_, _07644_);
  or (_11005_, _11003_, _11002_);
  or (_11007_, _11005_, _11001_);
  or (_11008_, _11007_, _07907_);
  nand (_11009_, _11008_, _10998_);
  nor (_11010_, _11009_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11010_, _10990_);
  and (_11011_, _07896_, word_in[22]);
  and (_11012_, _10508_, _07633_);
  and (_11013_, _10502_, _07624_);
  or (_11014_, _11013_, _11012_);
  and (_11015_, _10498_, _07636_);
  and (_11016_, _10494_, _07644_);
  or (_11017_, _11016_, _11015_);
  or (_11018_, _11017_, _11014_);
  or (_11019_, _11018_, _07907_);
  and (_11020_, _10523_, _07636_);
  and (_11021_, _10514_, _07644_);
  or (_11022_, _11021_, _11020_);
  and (_11023_, _10530_, _07633_);
  and (_11024_, _10519_, _07624_);
  or (_11025_, _11024_, _11023_);
  or (_11026_, _11025_, _11022_);
  or (_11027_, _11026_, _07863_);
  nand (_11028_, _11027_, _11019_);
  nor (_11029_, _11028_, _07896_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11029_, _11011_);
  and (_11030_, _07964_, word_in[24]);
  and (_11031_, _10544_, _07796_);
  and (_11032_, _10540_, _07794_);
  or (_11033_, _11032_, _11031_);
  and (_11034_, _11033_, _07938_);
  and (_11035_, _10554_, _07796_);
  and (_11036_, _10550_, _07794_);
  or (_11037_, _11036_, _11035_);
  and (_11038_, _11037_, _07944_);
  and (_11039_, _10566_, _07796_);
  and (_11040_, _10561_, _07794_);
  or (_11041_, _11040_, _11039_);
  and (_11042_, _11041_, _07973_);
  and (_11043_, _10578_, _07796_);
  and (_11044_, _10574_, _07794_);
  or (_11045_, _11044_, _11043_);
  and (_11046_, _11045_, _07981_);
  or (_11047_, _11046_, _11042_);
  or (_11048_, _11047_, _11038_);
  nor (_11049_, _11048_, _11034_);
  nor (_11050_, _11049_, _07964_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11050_, _11030_);
  and (_11051_, _07964_, word_in[25]);
  and (_11052_, _10595_, _07796_);
  and (_11053_, _10591_, _07794_);
  or (_11054_, _11053_, _11052_);
  and (_11055_, _11054_, _07938_);
  and (_11056_, _10607_, _07796_);
  and (_11057_, _10603_, _07794_);
  or (_11059_, _11057_, _11056_);
  and (_11060_, _11059_, _07944_);
  and (_11061_, _10617_, _07796_);
  and (_11062_, _10613_, _07794_);
  or (_11063_, _11062_, _11061_);
  and (_11064_, _11063_, _07973_);
  and (_11065_, _10629_, _07796_);
  and (_11066_, _10625_, _07794_);
  or (_11067_, _11066_, _11065_);
  and (_11068_, _11067_, _07981_);
  or (_11069_, _11068_, _11064_);
  or (_11070_, _11069_, _11060_);
  nor (_11071_, _11070_, _11055_);
  nor (_11072_, _11071_, _07964_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _11072_, _11051_);
  and (_11074_, _07964_, word_in[26]);
  and (_11075_, _10657_, _07796_);
  and (_11076_, _10652_, _07794_);
  or (_11077_, _11076_, _11075_);
  and (_11078_, _11077_, _07944_);
  and (_11079_, _10644_, _07796_);
  and (_11080_, _10639_, _07794_);
  or (_11081_, _11080_, _11079_);
  and (_11082_, _11081_, _07938_);
  and (_11083_, _10669_, _07796_);
  and (_11084_, _10665_, _07794_);
  or (_11085_, _11084_, _11083_);
  and (_11086_, _11085_, _07973_);
  and (_11087_, _10681_, _07796_);
  and (_11088_, _10676_, _07794_);
  or (_11089_, _11088_, _11087_);
  and (_11090_, _11089_, _07981_);
  or (_11091_, _11090_, _11086_);
  or (_11092_, _11091_, _11082_);
  nor (_11093_, _11092_, _11078_);
  nor (_11094_, _11093_, _07964_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _11094_, _11074_);
  and (_11096_, _07964_, word_in[27]);
  and (_11097_, _10696_, _07796_);
  and (_11098_, _10692_, _07794_);
  or (_11099_, _11098_, _11097_);
  and (_11100_, _11099_, _07938_);
  and (_11101_, _10735_, _07796_);
  and (_11102_, _10731_, _07794_);
  or (_11103_, _11102_, _11101_);
  and (_11104_, _11103_, _07944_);
  and (_11105_, _10723_, _07796_);
  and (_11106_, _10718_, _07794_);
  or (_11107_, _11106_, _11105_);
  and (_11108_, _11107_, _07973_);
  and (_11109_, _10708_, _07796_);
  and (_11110_, _10703_, _07794_);
  or (_11111_, _11110_, _11109_);
  and (_11113_, _11111_, _07981_);
  or (_11114_, _11113_, _11108_);
  or (_11116_, _11114_, _11104_);
  nor (_11117_, _11116_, _11100_);
  nor (_11118_, _11117_, _07964_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _11118_, _11096_);
  and (_11119_, _07964_, word_in[28]);
  and (_11120_, _10753_, _07796_);
  and (_11122_, _10749_, _07794_);
  or (_11123_, _11122_, _11120_);
  and (_11124_, _11123_, _07938_);
  and (_11125_, _10764_, _07796_);
  and (_11127_, _10760_, _07794_);
  or (_11128_, _11127_, _11125_);
  and (_11129_, _11128_, _07944_);
  and (_11130_, _10774_, _07796_);
  and (_11131_, _10770_, _07794_);
  or (_11132_, _11131_, _11130_);
  and (_11133_, _11132_, _07973_);
  and (_11134_, _10786_, _07796_);
  and (_11135_, _10781_, _07794_);
  or (_11136_, _11135_, _11134_);
  and (_11137_, _11136_, _07981_);
  or (_11139_, _11137_, _11133_);
  or (_11140_, _11139_, _11129_);
  nor (_11141_, _11140_, _11124_);
  nor (_11142_, _11141_, _07964_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _11142_, _11119_);
  and (_11143_, _07964_, word_in[29]);
  and (_11144_, _10801_, _07796_);
  and (_11145_, _10797_, _07794_);
  or (_11146_, _11145_, _11144_);
  and (_11147_, _11146_, _07938_);
  and (_11149_, _10812_, _07796_);
  and (_11151_, _10808_, _07794_);
  or (_11152_, _11151_, _11149_);
  and (_11153_, _11152_, _07944_);
  and (_11155_, _10823_, _07796_);
  and (_11156_, _10819_, _07794_);
  or (_11157_, _11156_, _11155_);
  and (_11158_, _11157_, _07973_);
  and (_11159_, _10834_, _07796_);
  and (_11160_, _10830_, _07794_);
  or (_11162_, _11160_, _11159_);
  and (_11163_, _11162_, _07981_);
  or (_11165_, _11163_, _11158_);
  or (_11166_, _11165_, _11153_);
  nor (_11167_, _11166_, _11147_);
  nor (_11168_, _11167_, _07964_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _11168_, _11143_);
  and (_11169_, _07964_, word_in[30]);
  and (_11170_, _10848_, _07796_);
  and (_11171_, _10844_, _07794_);
  or (_11172_, _11171_, _11170_);
  and (_11173_, _11172_, _07938_);
  and (_11174_, _10879_, _07796_);
  and (_11175_, _10875_, _07794_);
  or (_11176_, _11175_, _11174_);
  and (_11177_, _11176_, _07944_);
  and (_11178_, _10869_, _07796_);
  and (_11179_, _10865_, _07794_);
  or (_11180_, _11179_, _11178_);
  and (_11181_, _11180_, _07973_);
  and (_11182_, _10858_, _07796_);
  and (_11183_, _10854_, _07794_);
  or (_11184_, _11183_, _11182_);
  and (_11185_, _11184_, _07981_);
  or (_11186_, _11185_, _11181_);
  or (_11187_, _11186_, _11177_);
  nor (_11188_, _11187_, _11173_);
  nor (_11189_, _11188_, _07964_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _11189_, _11169_);
  not (_11190_, _06881_);
  not (_11191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_11192_, _06880_, _11191_);
  nor (_11193_, _11192_, _11190_);
  not (_11194_, _11193_);
  or (_11196_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_11197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_11199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _11197_);
  and (_11200_, _11199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_11202_, _11200_, _11196_);
  and (_11203_, _11202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_11204_, _11203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_11206_, _11205_, _11202_);
  and (_11207_, _11206_, _11204_);
  and (_11208_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_11209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_11211_, _11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_11212_, _11211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_11213_, _11212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_11214_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_11215_, _11214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_11216_, _11215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_11217_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_11218_, _11217_, _11216_);
  and (_11219_, _11218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_11220_, _11219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_11222_, _11220_, _11209_);
  and (_11223_, _11222_, _11208_);
  not (_11225_, _06882_);
  and (_11226_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_11227_, _11226_, _11202_);
  and (_11228_, _11227_, _11223_);
  or (_11230_, _11228_, _11207_);
  and (_11231_, _11230_, _11194_);
  and (_11232_, _11193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_11233_, _05807_, _10208_);
  and (_11234_, _11233_, _06888_);
  or (_11235_, _11234_, _11232_);
  or (_11236_, _11235_, _11231_);
  nand (_11237_, _11234_, _05938_);
  and (_11238_, _08133_, _05807_);
  and (_11239_, _11238_, _06888_);
  not (_11240_, _11239_);
  and (_11241_, _11240_, _11237_);
  and (_11242_, _11241_, _11236_);
  and (_11243_, _11239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_11245_, _11243_, _11242_);
  and (_09843_, _11245_, _05110_);
  or (_11246_, _06406_, _07153_);
  or (_11247_, _05473_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_11248_, _11247_, _05110_);
  and (_09877_, _11248_, _11246_);
  nand (_11249_, _06338_, _05473_);
  or (_11250_, _05473_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_11251_, _11250_, _05110_);
  and (_09897_, _11251_, _11249_);
  nand (_11252_, _06427_, _05473_);
  or (_11253_, _05473_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_11254_, _11253_, _05110_);
  and (_09900_, _11254_, _11252_);
  or (_11255_, _06271_, _07153_);
  or (_11256_, _05473_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_11257_, _11256_, _05110_);
  and (_09902_, _11257_, _11255_);
  nand (_11258_, _06315_, _05473_);
  or (_11259_, _05473_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_11260_, _11259_, _05110_);
  and (_09905_, _11260_, _11258_);
  and (_11261_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_11262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_11263_, _05846_, _11262_);
  not (_11264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_11265_, _11264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_11266_, _11265_, _11263_);
  nor (_11268_, _11266_, _11261_);
  or (_11269_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_11271_, _11269_, _05110_);
  nor (_10104_, _11271_, _11268_);
  not (_11272_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_11273_, _05464_, _11272_);
  nor (_11274_, _06054_, _05465_);
  or (_11275_, _11274_, _11273_);
  and (_10144_, _11275_, _05110_);
  not (_11276_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_11277_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _11276_);
  and (_10400_, _11277_, _05110_);
  nor (_11279_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_11280_, _11279_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_10460_, _11280_, _05110_);
  and (_11281_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11282_, _11281_);
  and (_11283_, _07070_, _06451_);
  and (_11284_, _11283_, _06873_);
  and (_11286_, _11284_, _06342_);
  or (_11287_, _07137_, _06823_);
  nor (_11288_, _11287_, _07074_);
  and (_11289_, _06811_, _06451_);
  and (_11290_, _07071_, _06276_);
  or (_11292_, _11290_, _07038_);
  and (_11293_, _11292_, _06460_);
  nor (_11294_, _11293_, _11289_);
  and (_11295_, _11294_, _11288_);
  or (_11296_, _07087_, _06452_);
  and (_11297_, _11296_, _06448_);
  nor (_11298_, _11297_, _06449_);
  nor (_11299_, _07041_, _06461_);
  nand (_11300_, _06852_, _07063_);
  and (_11301_, _07038_, _06864_);
  and (_11302_, _06825_, _06460_);
  nor (_11303_, _11302_, _11301_);
  and (_11304_, _11303_, _11300_);
  and (_11305_, _11304_, _11299_);
  and (_11306_, _11305_, _11298_);
  nand (_11307_, _11306_, _11295_);
  and (_11308_, _06872_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11309_, _11301_, _11308_);
  or (_11310_, _11309_, _06870_);
  and (_11311_, _11310_, _11307_);
  or (_11312_, _11311_, _11286_);
  nand (_11313_, _11312_, _05151_);
  and (_11314_, _11313_, _11282_);
  and (_11315_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2]);
  not (_11316_, _11315_);
  nand (_11317_, _11298_, _06440_);
  nand (_11319_, _11317_, _06870_);
  nor (_11320_, _11284_, _07056_);
  nand (_11321_, _11320_, _11319_);
  nand (_11322_, _11321_, _05151_);
  and (_11323_, _11322_, _11316_);
  nand (_11324_, _11323_, _05110_);
  nor (_10472_, _11324_, _11314_);
  nor (_11325_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_10517_, _11325_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_11326_, _10155_, _05797_);
  and (_11327_, _11326_, _05805_);
  or (_11328_, _11327_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_11329_, _06888_, _05808_);
  not (_11330_, _11329_);
  and (_11331_, _11330_, _11328_);
  nand (_11332_, _11327_, _05872_);
  and (_11333_, _11332_, _11331_);
  and (_11334_, _11329_, _06799_);
  or (_11335_, _11334_, _11333_);
  and (_10524_, _11335_, _05110_);
  nor (_11336_, _06205_, _06200_);
  and (_11337_, _06920_, _06909_);
  not (_11338_, _11337_);
  and (_11339_, _06909_, _06271_);
  not (_11340_, _06315_);
  and (_11341_, _11340_, _06294_);
  and (_11342_, _11341_, _11339_);
  and (_11343_, _06338_, _06271_);
  nor (_11344_, _06315_, _06294_);
  and (_11345_, _11344_, _11343_);
  nor (_11346_, _11345_, _11342_);
  and (_11347_, _11346_, _11338_);
  nor (_11348_, _11347_, _06427_);
  not (_11349_, _11348_);
  not (_11350_, _06922_);
  and (_11351_, _11341_, _11343_);
  and (_11353_, _06338_, _06928_);
  and (_11354_, _11341_, _11353_);
  nor (_11355_, _11354_, _11351_);
  nor (_11356_, _11355_, _11350_);
  and (_11357_, _06926_, _06362_);
  and (_11358_, _06920_, _11339_);
  and (_11359_, _11358_, _11357_);
  and (_11360_, _11343_, _06920_);
  nor (_11362_, _06924_, _06406_);
  nor (_11363_, _06384_, _06362_);
  and (_11365_, _11363_, _11362_);
  and (_11366_, _11365_, _11360_);
  nor (_11367_, _11366_, _11359_);
  not (_11368_, _11367_);
  nor (_11369_, _11368_, _11356_);
  and (_11370_, _11369_, _11349_);
  nor (_11371_, _06926_, _06916_);
  and (_11372_, _11344_, _11339_);
  and (_11373_, _11357_, _11372_);
  nor (_11374_, _11373_, _11354_);
  nor (_11376_, _11374_, _11371_);
  not (_11377_, _06916_);
  nor (_11378_, _11353_, _11339_);
  and (_11379_, _11378_, _06920_);
  not (_11380_, _11379_);
  and (_11381_, _11380_, _11346_);
  nor (_11382_, _11381_, _11377_);
  nor (_11383_, _11382_, _11376_);
  and (_11384_, _11383_, _11370_);
  not (_11385_, _11365_);
  nor (_11386_, _06338_, _06315_);
  and (_11387_, _11386_, _06294_);
  nor (_11388_, _11358_, _11387_);
  nor (_11389_, _11388_, _11385_);
  not (_11391_, _11389_);
  not (_11393_, _06384_);
  and (_11394_, _11393_, _06362_);
  and (_11395_, _11394_, _11362_);
  and (_11396_, _11353_, _06920_);
  and (_11397_, _11396_, _06924_);
  nor (_11398_, _11397_, _11395_);
  and (_11399_, _11398_, _11391_);
  and (_11400_, _11387_, _06928_);
  not (_11401_, _11400_);
  nor (_11402_, _06926_, _06915_);
  nor (_11403_, _11402_, _11401_);
  not (_11404_, _06927_);
  nor (_11405_, _11360_, _06911_);
  nor (_11406_, _11405_, _11404_);
  nor (_11407_, _11406_, _11403_);
  and (_11408_, _11407_, _11399_);
  not (_11409_, _11351_);
  nor (_11410_, _11371_, _11409_);
  not (_11411_, _11357_);
  and (_11412_, _11386_, _06918_);
  and (_11414_, _11412_, _06928_);
  nor (_11415_, _11414_, _06910_);
  nor (_11416_, _11415_, _11411_);
  nor (_11417_, _11416_, _11410_);
  and (_11418_, _11417_, _11408_);
  nor (_11419_, _11387_, _11337_);
  nor (_11420_, _11419_, _06928_);
  nor (_11421_, _11420_, _06929_);
  and (_11422_, _06914_, _06406_);
  not (_11423_, _11422_);
  nor (_11424_, _11423_, _11421_);
  not (_11425_, _11424_);
  nor (_11426_, _11351_, _11396_);
  nor (_11427_, _11426_, _11385_);
  not (_11428_, _11427_);
  and (_11429_, _11342_, _06927_);
  and (_11430_, _11396_, _06916_);
  nor (_11431_, _11430_, _11429_);
  and (_11432_, _11431_, _11428_);
  and (_11433_, _11432_, _11425_);
  and (_11434_, _11433_, _11418_);
  and (_11435_, _11378_, _06910_);
  nand (_11436_, _11435_, _11365_);
  and (_11437_, _11345_, _11357_);
  not (_11438_, _11437_);
  and (_11439_, _11438_, _11436_);
  and (_11440_, _06910_, _06338_);
  and (_11441_, _11440_, _06916_);
  not (_11442_, _11441_);
  and (_11443_, _11358_, _06927_);
  nor (_11444_, _11342_, _11396_);
  nor (_11445_, _11444_, _11411_);
  nor (_11446_, _11445_, _11443_);
  and (_11447_, _11446_, _11442_);
  and (_11448_, _11447_, _11439_);
  and (_11449_, _11344_, _11353_);
  nor (_11450_, _11449_, _11360_);
  nor (_11451_, _11450_, _11411_);
  nor (_11452_, _11449_, _11358_);
  nor (_11453_, _11452_, _11377_);
  nor (_11454_, _11453_, _11451_);
  and (_11455_, _11339_, _06910_);
  and (_11456_, _11365_, _11455_);
  and (_11457_, _11354_, _11365_);
  nor (_11458_, _11457_, _11456_);
  not (_11459_, _11458_);
  and (_11460_, _11337_, _06928_);
  and (_11461_, _06338_, _11340_);
  and (_11462_, _11461_, _06918_);
  nor (_11463_, _11462_, _11460_);
  nor (_11464_, _11463_, _11385_);
  nor (_11465_, _11464_, _11459_);
  and (_11466_, _11465_, _11454_);
  and (_11467_, _11466_, _11448_);
  and (_11468_, _11467_, _11434_);
  and (_11469_, _11468_, _11384_);
  nor (_11470_, _11469_, _06255_);
  not (_11471_, _11469_);
  and (_11472_, _11400_, _06922_);
  not (_11473_, _11472_);
  and (_11474_, _06406_, _06384_);
  or (_11475_, _11474_, _06924_);
  and (_11476_, _11475_, _11358_);
  nor (_11477_, _11476_, _11456_);
  and (_11478_, _11477_, _11473_);
  and (_11479_, _11478_, _11369_);
  and (_11480_, _11479_, _11448_);
  nand (_11481_, _11480_, _11471_);
  and (_11482_, _11481_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_11483_, _11469_, _06255_);
  nor (_11484_, _11483_, _11470_);
  and (_11485_, _11484_, _11482_);
  nor (_11486_, _11485_, _11470_);
  nor (_11487_, _11486_, _06200_);
  and (_11488_, _11487_, _06201_);
  nor (_11489_, _11487_, _06201_);
  nor (_11490_, _11489_, _11488_);
  nor (_11491_, _11490_, _11336_);
  and (_11492_, _06256_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_11493_, _11492_, _11336_);
  nor (_11494_, _11493_, _11480_);
  or (_11495_, _11494_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_11497_, _11495_, _11491_);
  and (_10539_, _11497_, _05110_);
  not (_11498_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  not (_11499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_11500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_11501_, _11500_, _11499_);
  nor (_11502_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_11503_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_11504_, _11503_, _11502_);
  and (_11505_, _11504_, _11501_);
  and (_11506_, _11505_, _11498_);
  and (_11507_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_11508_, _11507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_10558_, _11508_, _05110_);
  not (_11510_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand (_11511_, _05474_, _11510_);
  nand (_11512_, _11511_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_11513_, _11512_, _11506_);
  and (_10562_, _11513_, _05110_);
  and (_10567_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _05110_);
  not (_11515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_11516_, _06880_, _11515_);
  or (_11517_, _11516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_11518_, _11517_, _11326_);
  not (_11519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_11520_, _05488_, _11519_);
  nand (_11521_, _11520_, _11326_);
  or (_11523_, _11521_, _05784_);
  and (_11524_, _11523_, _11518_);
  or (_11525_, _11524_, _11329_);
  nand (_11526_, _11329_, _05841_);
  and (_11527_, _11526_, _05110_);
  and (_10582_, _11527_, _11525_);
  and (_11528_, _11326_, _08133_);
  nand (_11529_, _11528_, _05872_);
  or (_11530_, _11528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_11532_, _11530_, _11330_);
  and (_11533_, _11532_, _11529_);
  nor (_11535_, _11330_, _06054_);
  or (_11536_, _11535_, _11533_);
  and (_10585_, _11536_, _05110_);
  and (_11537_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_11538_, _11537_, _10209_);
  and (_11539_, _11538_, _11326_);
  not (_11540_, _11326_);
  or (_11541_, _11540_, _10212_);
  and (_11542_, _11541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_11543_, _11542_, _11329_);
  or (_11544_, _11543_, _11539_);
  nand (_11545_, _11329_, _05334_);
  and (_11546_, _11545_, _05110_);
  and (_10587_, _11546_, _11544_);
  and (_11547_, _11326_, _06632_);
  not (_11548_, _05866_);
  nand (_11549_, _11326_, _05401_);
  or (_11550_, _11549_, _11548_);
  and (_11551_, _11550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_11552_, _11551_, _11329_);
  or (_11553_, _11552_, _11547_);
  nand (_11554_, _11329_, _06088_);
  and (_11555_, _11554_, _05110_);
  and (_10597_, _11555_, _11553_);
  and (_11556_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_11557_, _11556_, _08245_);
  and (_11558_, _11557_, _11326_);
  not (_11559_, _10169_);
  nand (_11560_, _11326_, _11559_);
  and (_11561_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_11562_, _11561_, _11329_);
  or (_11563_, _11562_, _11558_);
  nand (_11564_, _11329_, _06229_);
  and (_11565_, _11564_, _05110_);
  and (_10600_, _11565_, _11563_);
  not (_11566_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_11567_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor (_11568_, _11567_, _11566_);
  and (_11569_, _11567_, _11566_);
  nor (_11570_, _11569_, _11568_);
  not (_11571_, _11570_);
  and (_11572_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_11573_, _11572_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_11574_, _11572_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_11575_, _11574_, _11573_);
  or (_11576_, _11575_, _11567_);
  and (_11577_, _11576_, _11571_);
  nor (_11578_, _11568_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_11579_, _11568_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_11580_, _11579_, _11578_);
  or (_11581_, _11573_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_03099_, _11581_, _05110_);
  and (_11582_, _03099_, _11580_);
  and (_10620_, _11582_, _11577_);
  and (_10641_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _05110_);
  nor (_11583_, _11240_, _06229_);
  nor (_11584_, _11239_, _11234_);
  and (_11585_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_11586_, _11585_, _11202_);
  and (_11587_, _11586_, _11223_);
  nand (_11588_, _11218_, _11202_);
  nor (_11589_, _11588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_11590_, _11588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_11591_, _11590_, _11193_);
  or (_11592_, _11591_, _11589_);
  or (_11593_, _11592_, _11587_);
  or (_11594_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_11595_, _11594_, _11593_);
  and (_11596_, _11595_, _11584_);
  and (_11597_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_11598_, _11597_, _11596_);
  or (_11599_, _11598_, _11583_);
  and (_10645_, _11599_, _05110_);
  not (_11600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_11601_, _11216_, _11202_);
  nor (_11602_, _11601_, _11600_);
  or (_11603_, _11602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_11604_, _11603_, _11588_);
  or (_11605_, _11604_, _11193_);
  and (_11606_, _11202_, _11225_);
  and (_11607_, _11606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_11608_, _11607_, _11223_);
  or (_11609_, _11608_, _11605_);
  or (_11610_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_11611_, _11610_, _11609_);
  and (_11612_, _11611_, _11584_);
  nor (_11613_, _11240_, _05938_);
  and (_11614_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_11615_, _11614_, _11613_);
  or (_11616_, _11615_, _11612_);
  and (_10649_, _11616_, _05110_);
  and (_11617_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07601_);
  and (_11618_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_11619_, _11618_, _11617_);
  and (_10654_, _11619_, _05110_);
  and (_11620_, _11239_, _06799_);
  and (_11621_, _11601_, _11600_);
  nor (_11622_, _11621_, _11602_);
  or (_11623_, _11622_, _11193_);
  and (_11625_, _11606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_11626_, _11625_, _11223_);
  or (_11627_, _11626_, _11623_);
  not (_11628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_11629_, _11193_, _11628_);
  and (_11630_, _11629_, _11627_);
  and (_11631_, _11630_, _11584_);
  and (_11632_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_11633_, _11632_, _11631_);
  or (_11634_, _11633_, _11620_);
  and (_10660_, _11634_, _05110_);
  and (_11635_, _06380_, _06311_);
  and (_11636_, _11635_, _06423_);
  and (_11637_, _11325_, _05475_);
  and (_11638_, _11637_, _06266_);
  and (_11639_, _06334_, _06289_);
  and (_11640_, _11639_, _11638_);
  and (_11641_, _06402_, _06357_);
  and (_11642_, _11641_, _11640_);
  and (_10663_, _11642_, _11636_);
  and (_11644_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_11645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_11646_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_11647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_11648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_11650_, _11648_, _11646_);
  and (_11651_, _11650_, _11647_);
  nor (_11652_, _11651_, _11646_);
  nor (_11653_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_11654_, _11653_, _11645_);
  not (_11655_, _11654_);
  nor (_11656_, _11655_, _11652_);
  nor (_11657_, _11656_, _11645_);
  not (_11658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_11660_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_11661_, _11660_, _11658_);
  and (_11662_, _11661_, _11657_);
  and (_11664_, _11657_, _11660_);
  nor (_11665_, _11664_, _11658_);
  nor (_11666_, _11665_, _11662_);
  not (_11667_, _11666_);
  not (_11669_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_11670_, _11657_, _11669_);
  nor (_11671_, _11657_, _11669_);
  nor (_11672_, _11671_, _11670_);
  not (_11673_, _11672_);
  nor (_11675_, _11650_, _11647_);
  nor (_11676_, _11675_, _11651_);
  nand (_11677_, _11676_, _11471_);
  not (_11678_, _11677_);
  nor (_11680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_11681_, _11680_, _11647_);
  and (_11682_, _11681_, _11481_);
  or (_11683_, _11676_, _11471_);
  and (_11684_, _11683_, _11677_);
  and (_11685_, _11684_, _11682_);
  or (_11686_, _11685_, _11678_);
  and (_11687_, _11655_, _11652_);
  nor (_11688_, _11687_, _11656_);
  and (_11689_, _11688_, _11686_);
  and (_11690_, _11689_, _11673_);
  not (_11691_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_11692_, _11670_, _11691_);
  or (_11693_, _11692_, _11664_);
  and (_11695_, _11693_, _11690_);
  and (_11696_, _11695_, _11667_);
  nor (_11698_, _11695_, _11667_);
  nor (_11699_, _11698_, _11696_);
  or (_11700_, _11699_, _07437_);
  or (_11701_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_11703_, _11701_, _11510_);
  and (_11705_, _11703_, _11700_);
  or (_11706_, _11705_, _11644_);
  and (_10679_, _11706_, _05110_);
  and (_11708_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_11709_, _11708_, _11202_);
  and (_11710_, _11709_, _11223_);
  and (_11711_, _11220_, _11202_);
  and (_11712_, _11711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_11713_, _11711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_11714_, _11713_, _11712_);
  or (_11715_, _11714_, _11193_);
  or (_11716_, _11715_, _11710_);
  nor (_11717_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_11719_, _11717_, _11234_);
  and (_11720_, _11719_, _11716_);
  and (_11721_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_11722_, _11721_, _11239_);
  or (_11723_, _11722_, _11720_);
  nand (_11724_, _11239_, _05334_);
  and (_11726_, _11724_, _05110_);
  and (_10684_, _11726_, _11723_);
  and (_11727_, _06824_, _06813_);
  and (_11728_, _11727_, _06451_);
  and (_11729_, _07038_, _06277_);
  and (_11730_, _11729_, _06451_);
  nor (_11731_, _11730_, _07147_);
  not (_11732_, _11731_);
  nor (_11734_, _11732_, _11728_);
  nor (_11735_, _11734_, _06239_);
  not (_11736_, _11314_);
  and (_11737_, _07077_, _06277_);
  or (_11738_, _11737_, _07088_);
  or (_11740_, _11738_, _07122_);
  nand (_11741_, _07115_, _06276_);
  and (_11742_, _07077_, _06276_);
  nor (_11743_, _11742_, _07081_);
  nand (_11744_, _11743_, _11741_);
  or (_11745_, _11744_, _07086_);
  nor (_11746_, _11745_, _11740_);
  not (_11747_, _07076_);
  nand (_11748_, _06825_, _06810_);
  and (_11749_, _06856_, _06810_);
  nor (_11750_, _11749_, _11301_);
  and (_11751_, _11750_, _11748_);
  and (_11752_, _11751_, _11747_);
  and (_11753_, _11752_, _11734_);
  and (_11754_, _06864_, _06438_);
  or (_11755_, _11754_, _07139_);
  and (_11756_, _11292_, _06810_);
  nor (_11757_, _11756_, _11755_);
  or (_11758_, _07069_, _06463_);
  nand (_11759_, _11758_, _06810_);
  not (_11760_, _11759_);
  and (_11761_, _06941_, _06277_);
  nor (_11762_, _11761_, _11760_);
  and (_11763_, _11762_, _11757_);
  nor (_11764_, _07116_, _07051_);
  nor (_11765_, _07132_, _07127_);
  and (_11766_, _11765_, _11764_);
  nor (_11767_, _06845_, _06817_);
  and (_11768_, _11767_, _07110_);
  and (_11769_, _11768_, _11766_);
  and (_11770_, _11769_, _11763_);
  and (_11771_, _11770_, _11753_);
  nand (_11772_, _11771_, _11746_);
  nand (_11773_, _11772_, _06870_);
  nor (_11774_, _11309_, _11284_);
  nand (_11775_, _11774_, _11773_);
  nand (_11776_, _11775_, _05151_);
  and (_11777_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11778_, _11777_);
  and (_11779_, _11778_, _11776_);
  and (_11780_, _11779_, _11736_);
  and (_11781_, _11780_, _11323_);
  nor (_11782_, _10176_, _10215_);
  nor (_11783_, _11782_, _10220_);
  or (_11784_, _11783_, _05419_);
  nand (_11785_, _11783_, _05419_);
  and (_11786_, _11785_, _11784_);
  nor (_11787_, _10180_, _10177_);
  nand (_11788_, _11787_, _05390_);
  and (_11789_, _05433_, _05337_);
  and (_11790_, _11789_, _06173_);
  and (_11791_, _11790_, _05461_);
  and (_11792_, _11791_, _11788_);
  or (_11793_, _11787_, _05390_);
  nor (_11794_, _06366_, _05375_);
  and (_11795_, _06366_, _05375_);
  nor (_11796_, _11795_, _11794_);
  and (_11797_, _11796_, _11793_);
  and (_11798_, _11797_, _11792_);
  and (_11799_, _11798_, _11786_);
  and (_11800_, _11799_, _06088_);
  not (_11801_, _11783_);
  not (_11802_, _06366_);
  and (_11803_, _11787_, _11802_);
  and (_11804_, _11803_, _11801_);
  nand (_11805_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_11806_, _11787_, _06366_);
  and (_11807_, _11806_, _11783_);
  nand (_11808_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_11809_, _11808_, _11805_);
  nor (_11810_, _11787_, _11802_);
  and (_11811_, _11810_, _11801_);
  nand (_11812_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_11813_, _11787_, _06366_);
  and (_11814_, _11813_, _11783_);
  nand (_11815_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_11816_, _11815_, _11812_);
  and (_11817_, _11816_, _11809_);
  not (_11818_, _11799_);
  and (_11819_, _11813_, _11801_);
  nand (_11820_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_11821_, _11803_, _11783_);
  nand (_11822_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_11823_, _11822_, _11820_);
  and (_11824_, _11806_, _11801_);
  nand (_11825_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_11826_, _11810_, _11783_);
  nand (_11827_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_11828_, _11827_, _11825_);
  and (_11829_, _11828_, _11823_);
  and (_11830_, _11829_, _11818_);
  and (_11831_, _11830_, _11817_);
  nor (_11832_, _11831_, _11800_);
  nand (_11833_, _11832_, _11781_);
  nand (_11834_, _11778_, _11776_);
  and (_11835_, _11323_, _11314_);
  nand (_11836_, _11835_, _11834_);
  or (_11837_, _11836_, _07470_);
  and (_11838_, _11837_, _11833_);
  and (_11839_, _11834_, _11736_);
  nand (_11840_, _11839_, _11323_);
  nand (_11841_, _07206_, _08272_);
  or (_11842_, _11841_, _06088_);
  and (_11843_, _07206_, _08272_);
  nand (_11844_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_11845_, _11844_, _11842_);
  nand (_11846_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or (_11847_, _11841_, _06229_);
  and (_11848_, _11847_, _11846_);
  nand (_11849_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or (_11850_, _11841_, _05938_);
  and (_11851_, _11850_, _11849_);
  not (_11852_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  or (_11853_, _11843_, _05369_);
  or (_11854_, _11841_, _06798_);
  nand (_11855_, _11854_, _11853_);
  nor (_11856_, _11855_, _11852_);
  and (_11857_, _11856_, _11851_);
  and (_11858_, _11857_, _11848_);
  and (_11859_, _11858_, _11845_);
  or (_11860_, _11858_, _11845_);
  not (_11861_, _11860_);
  nor (_11862_, _11861_, _11859_);
  or (_11863_, _11862_, _05341_);
  and (_11864_, _11863_, _05384_);
  or (_11865_, _11864_, _11843_);
  and (_11866_, _11865_, _11842_);
  or (_11867_, _11866_, _11840_);
  nand (_11868_, _11835_, _11779_);
  or (_11869_, _11868_, _11787_);
  and (_11870_, _11869_, _11867_);
  and (_11871_, _11870_, _11838_);
  or (_11872_, _11871_, _05390_);
  nand (_11873_, _11870_, _11838_);
  or (_11874_, _11873_, _05389_);
  and (_11875_, _11874_, _11872_);
  and (_11876_, _11839_, _11323_);
  nor (_11877_, _11841_, _06054_);
  or (_11878_, _11841_, _05334_);
  nand (_11879_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_11880_, _11879_, _11878_);
  and (_11881_, _11880_, _11859_);
  and (_11882_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_11883_, _11882_, _11877_);
  and (_11884_, _11883_, _11881_);
  nor (_11885_, _11883_, _11881_);
  or (_11886_, _11885_, _11884_);
  nand (_11887_, _11886_, _05790_);
  nand (_11888_, _11887_, _05423_);
  and (_11889_, _11888_, _11841_);
  or (_11890_, _11889_, _11877_);
  nand (_11891_, _11890_, _11876_);
  nand (_11892_, _11799_, _06054_);
  nand (_11893_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nand (_11894_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_11895_, _11894_, _11893_);
  nand (_11896_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nand (_11897_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_11898_, _11897_, _11896_);
  and (_11899_, _11898_, _11895_);
  nand (_11900_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nand (_11901_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_11902_, _11901_, _11900_);
  nand (_11903_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand (_11904_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_11905_, _11904_, _11903_);
  and (_11906_, _11905_, _11902_);
  and (_11907_, _11906_, _11818_);
  nand (_11908_, _11907_, _11899_);
  and (_11909_, _11908_, _11892_);
  nand (_11910_, _11909_, _11781_);
  or (_11911_, _11836_, _07507_);
  and (_11912_, _11911_, _11910_);
  or (_11914_, _11779_, _11736_);
  nor (_11915_, _11780_, _11323_);
  nand (_11916_, _11915_, _11914_);
  and (_11917_, _11916_, _11912_);
  and (_11918_, _11917_, _11891_);
  and (_11919_, _11918_, _06121_);
  nand (_11920_, _11917_, _11891_);
  and (_11921_, _11920_, _05433_);
  nor (_11922_, _11921_, _11919_);
  or (_11923_, _11868_, _11783_);
  or (_11924_, _11836_, _07490_);
  and (_11925_, _11924_, _11923_);
  and (_11926_, _11799_, _05334_);
  and (_11927_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_11928_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_11929_, _11928_, _11927_);
  and (_11930_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_11931_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_11932_, _11931_, _11930_);
  and (_11933_, _11932_, _11929_);
  nand (_11934_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nand (_11935_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_11936_, _11935_, _11934_);
  nand (_11937_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nand (_11938_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_11939_, _11938_, _11937_);
  and (_11941_, _11939_, _11936_);
  and (_11942_, _11941_, _11818_);
  and (_11943_, _11942_, _11933_);
  nor (_11944_, _11943_, _11926_);
  nand (_11945_, _11944_, _11781_);
  not (_11946_, _11323_);
  and (_11948_, _11946_, _11314_);
  nor (_11949_, _11880_, _11859_);
  or (_11950_, _11949_, _11881_);
  nand (_11951_, _11950_, _05790_);
  nand (_11952_, _11951_, _05408_);
  nand (_11953_, _11952_, _11841_);
  nand (_11954_, _11953_, _11878_);
  and (_11955_, _11954_, _11876_);
  nor (_11956_, _11955_, _11948_);
  and (_11957_, _11956_, _11945_);
  nand (_11958_, _11957_, _11925_);
  or (_11959_, _11958_, _05418_);
  and (_11960_, _11957_, _11925_);
  or (_11961_, _11960_, _05419_);
  and (_11962_, _11961_, _11959_);
  and (_11963_, _11843_, _05901_);
  nor (_11964_, _11841_, _05841_);
  and (_11965_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_11966_, _11965_, _11964_);
  nand (_11967_, _11966_, _11884_);
  not (_11968_, _11967_);
  and (_11969_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_11970_, _11969_, _11968_);
  or (_11971_, _11969_, _11968_);
  and (_11972_, _11971_, _05790_);
  nand (_11973_, _11972_, _11970_);
  and (_11974_, _11841_, _05452_);
  and (_11975_, _11974_, _11973_);
  nor (_11976_, _11975_, _11963_);
  nand (_11977_, _11976_, _11839_);
  nand (_11978_, _11799_, _05901_);
  nand (_11979_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand (_11981_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_11982_, _11981_, _11979_);
  nand (_11984_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand (_11985_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_11986_, _11985_, _11984_);
  and (_11987_, _11986_, _11982_);
  nand (_11988_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand (_11989_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_11990_, _11989_, _11988_);
  nand (_11992_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand (_11993_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_11994_, _11993_, _11992_);
  and (_11995_, _11994_, _11990_);
  and (_11996_, _11995_, _11818_);
  nand (_11997_, _11996_, _11987_);
  and (_11998_, _11997_, _11978_);
  nand (_11999_, _11998_, _11781_);
  nor (_12000_, _05474_, _05454_);
  and (_12001_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  not (_12002_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_12003_, _06251_, _12002_);
  nor (_12004_, _12003_, _12001_);
  and (_12005_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_12006_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_12007_, _12006_, _12005_);
  and (_12008_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_12009_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_12010_, _12009_, _12008_);
  and (_12011_, _12010_, _12007_);
  and (_12012_, _12011_, _12004_);
  nor (_12013_, _12012_, _07437_);
  nor (_12014_, _12013_, _12000_);
  or (_12016_, _12014_, _11914_);
  and (_12017_, _12016_, _11323_);
  and (_12018_, _12017_, _11999_);
  and (_12020_, _12018_, _11977_);
  and (_12021_, _12020_, _05460_);
  nor (_12022_, _12020_, _05460_);
  nor (_12023_, _12022_, _12021_);
  or (_12024_, _11966_, _11884_);
  nand (_12025_, _12024_, _11967_);
  nand (_12026_, _12025_, _05790_);
  nand (_12027_, _12026_, _05439_);
  and (_12028_, _12027_, _11841_);
  or (_12029_, _12028_, _11964_);
  nand (_12030_, _12029_, _11876_);
  nand (_12031_, _11799_, _05841_);
  nand (_12032_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nand (_12033_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_12034_, _12033_, _12032_);
  nand (_12035_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nand (_12036_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_12037_, _12036_, _12035_);
  and (_12038_, _12037_, _12034_);
  nand (_12039_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nand (_12040_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_12041_, _12040_, _12039_);
  nand (_12042_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nand (_12043_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_12044_, _12043_, _12042_);
  and (_12045_, _12044_, _12041_);
  and (_12046_, _12045_, _11818_);
  nand (_12048_, _12046_, _12038_);
  and (_12049_, _12048_, _12031_);
  nand (_12050_, _12049_, _11781_);
  and (_12051_, _12050_, _12030_);
  nor (_12052_, _05474_, _05441_);
  and (_12053_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not (_12054_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_12056_, _06251_, _12054_);
  nor (_12057_, _12056_, _12053_);
  and (_12058_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_12059_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_12060_, _12059_, _12058_);
  and (_12061_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_12062_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_12063_, _12062_, _12061_);
  and (_12064_, _12063_, _12060_);
  and (_12065_, _12064_, _12057_);
  nor (_12066_, _12065_, _07437_);
  nor (_12067_, _12066_, _12052_);
  nor (_12068_, _12067_, _11836_);
  nor (_12070_, _11915_, _12068_);
  nand (_12071_, _12070_, _12051_);
  or (_12072_, _12071_, _05447_);
  and (_12073_, _12070_, _12051_);
  or (_12074_, _12073_, _05448_);
  and (_12075_, _12074_, _12072_);
  and (_12077_, _12075_, _12023_);
  and (_12078_, _12077_, _11962_);
  and (_12080_, _12078_, _11922_);
  and (_12082_, _12080_, _11875_);
  not (_12083_, _05867_);
  and (_12084_, _12083_, _05806_);
  and (_12086_, _12084_, _12082_);
  and (_12087_, _12086_, _11735_);
  not (_12088_, _12087_);
  not (_12089_, _06870_);
  nor (_12090_, _07105_, _06866_);
  nor (_12091_, _12090_, _12089_);
  not (_12092_, _06997_);
  not (_12093_, _11284_);
  not (_12094_, _06873_);
  or (_12095_, _11728_, _07147_);
  nor (_12096_, _12095_, _11730_);
  nor (_12097_, _12096_, _12094_);
  nor (_12098_, _12096_, _12089_);
  nor (_12099_, _12098_, _12097_);
  and (_12100_, _12099_, _12093_);
  and (_12101_, _07396_, _05696_);
  and (_12102_, _07309_, _06640_);
  nand (_12103_, _12102_, _12101_);
  nor (_12104_, _12103_, _07211_);
  and (_12105_, _12104_, _06516_);
  and (_12106_, _12105_, _12100_);
  and (_12108_, _12106_, _06759_);
  and (_12109_, _12108_, _12092_);
  nor (_12111_, _11735_, _06436_);
  nor (_12112_, _12111_, _12093_);
  and (_12114_, _12112_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_12115_, _11735_, _05185_);
  nor (_12117_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_12118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_12119_, _12118_, _12117_);
  nor (_12120_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_12121_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_12123_, _12121_, _12120_);
  and (_12125_, _12123_, _12119_);
  and (_12126_, _12125_, _11286_);
  or (_12127_, _12126_, _12115_);
  or (_12128_, _12127_, _12114_);
  nor (_12130_, _12128_, _12109_);
  and (_12131_, _06811_, _06431_);
  not (_12132_, _12131_);
  and (_12134_, _06825_, _06464_);
  nor (_12135_, _12134_, _06812_);
  and (_12137_, _12135_, _12132_);
  and (_12138_, _07138_, _06451_);
  and (_12140_, _07087_, _06451_);
  or (_12141_, _12140_, _11728_);
  or (_12142_, _12141_, _12138_);
  nor (_12144_, _12142_, _06828_);
  and (_12145_, _12144_, _12137_);
  not (_12146_, _12145_);
  and (_12147_, _12146_, _12130_);
  not (_12148_, _12147_);
  not (_12149_, _07073_);
  and (_12150_, _12149_, _06451_);
  nor (_12151_, _12150_, _11732_);
  nor (_12153_, _12151_, _12130_);
  not (_12154_, _11301_);
  and (_12156_, _07087_, _06448_);
  and (_12158_, _06451_, _06438_);
  nor (_12159_, _12158_, _12156_);
  and (_12160_, _12159_, _12154_);
  not (_12162_, _12160_);
  nor (_12163_, _12162_, _12153_);
  and (_12165_, _12163_, _12148_);
  nor (_12166_, _11309_, _06873_);
  nor (_12168_, _12166_, _12165_);
  nor (_12169_, _12168_, _12091_);
  nor (_12171_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_12172_, _12171_);
  nor (_12173_, _12172_, _10176_);
  and (_12175_, _12173_, _10211_);
  not (_12176_, _12175_);
  and (_12177_, _12176_, _12112_);
  not (_12178_, _06628_);
  and (_12179_, _06638_, _12178_);
  not (_12180_, _12179_);
  and (_12181_, _12180_, _11286_);
  nor (_12182_, _12181_, _12177_);
  not (_12183_, _12182_);
  nor (_12184_, _12183_, _12169_);
  and (_12185_, _11780_, _11946_);
  nor (_12186_, _11856_, _11851_);
  nor (_12187_, _12186_, _11857_);
  nor (_12188_, _12187_, _05341_);
  nor (_12189_, _12188_, _05346_);
  nor (_12190_, _12189_, _11843_);
  not (_12192_, _12190_);
  and (_12193_, _12192_, _11850_);
  not (_12194_, _12193_);
  and (_12195_, _12194_, _11876_);
  nor (_12197_, _12195_, _12185_);
  or (_12198_, _11836_, _07439_);
  nand (_12200_, _11799_, _05938_);
  nand (_12201_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nand (_12203_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_12204_, _12203_, _12201_);
  nand (_12205_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nand (_12207_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_12208_, _12207_, _12205_);
  and (_12209_, _12208_, _12204_);
  nand (_12210_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nand (_12211_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_12212_, _12211_, _12210_);
  nand (_12213_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand (_12214_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_12215_, _12214_, _12213_);
  and (_12216_, _12215_, _12212_);
  and (_12217_, _12216_, _11818_);
  nand (_12219_, _12217_, _12209_);
  and (_12220_, _12219_, _12200_);
  nand (_12221_, _12220_, _11781_);
  or (_12222_, _11868_, _06445_);
  and (_12223_, _12222_, _12221_);
  and (_12224_, _12223_, _12198_);
  and (_12225_, _12224_, _12197_);
  or (_12227_, _12225_, _05365_);
  nand (_12228_, _12224_, _12197_);
  or (_12229_, _12228_, _05486_);
  nand (_12230_, _12229_, _12227_);
  nand (_12231_, _11799_, _06229_);
  nand (_12232_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nand (_12233_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_12234_, _12233_, _12232_);
  nand (_12235_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nand (_12236_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_12237_, _12236_, _12235_);
  and (_12239_, _12237_, _12234_);
  nand (_12240_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nand (_12241_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_12242_, _12241_, _12240_);
  nand (_12243_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nand (_12245_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_12246_, _12245_, _12243_);
  and (_12248_, _12246_, _12242_);
  and (_12249_, _12248_, _11818_);
  nand (_12250_, _12249_, _12239_);
  and (_12252_, _12250_, _12231_);
  nand (_12253_, _12252_, _11781_);
  or (_12254_, _11836_, _07454_);
  and (_12255_, _12254_, _12253_);
  nor (_12256_, _11857_, _11848_);
  or (_12257_, _12256_, _11858_);
  and (_12258_, _12257_, _05790_);
  or (_12259_, _12258_, _05393_);
  nand (_12260_, _12259_, _11841_);
  nand (_12262_, _12260_, _11847_);
  nand (_12263_, _12262_, _11876_);
  not (_12264_, _06411_);
  or (_12265_, _11868_, _12264_);
  and (_12266_, _12265_, _12263_);
  and (_12268_, _12266_, _12255_);
  or (_12269_, _12268_, _05401_);
  nand (_12270_, _12266_, _12255_);
  or (_12272_, _12270_, _05485_);
  nand (_12273_, _12272_, _12269_);
  and (_12274_, _11799_, _06798_);
  nand (_12275_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nand (_12276_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_12277_, _12276_, _12275_);
  nand (_12278_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand (_12279_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_12280_, _12279_, _12278_);
  and (_12281_, _12280_, _12277_);
  nand (_12282_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nand (_12283_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_12284_, _12283_, _12282_);
  nand (_12285_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nand (_12286_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_12287_, _12286_, _12285_);
  and (_12288_, _12287_, _12284_);
  and (_12289_, _12288_, _11818_);
  and (_12290_, _12289_, _12281_);
  nor (_12291_, _12290_, _12274_);
  nand (_12292_, _12291_, _11781_);
  nor (_12294_, _05474_, _05234_);
  and (_12295_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  not (_12297_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_12298_, _06251_, _12297_);
  nor (_12300_, _12298_, _12295_);
  and (_12301_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_12303_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_12304_, _12303_, _12301_);
  and (_12305_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_12307_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_12308_, _12307_, _12305_);
  and (_12310_, _12308_, _12304_);
  and (_12311_, _12310_, _12300_);
  nor (_12312_, _12311_, _07437_);
  nor (_12313_, _12312_, _12294_);
  or (_12314_, _12313_, _11836_);
  and (_12315_, _12314_, _12292_);
  and (_12316_, _11855_, _11852_);
  nor (_12318_, _12316_, _11856_);
  nor (_12319_, _12318_, _05341_);
  nor (_12321_, _12319_, _05370_);
  nor (_12322_, _12321_, _11843_);
  not (_12323_, _12322_);
  and (_12324_, _12323_, _11854_);
  or (_12325_, _12324_, _11840_);
  or (_12326_, _11868_, _11802_);
  and (_12327_, _12326_, _12325_);
  nand (_12328_, _12327_, _12315_);
  and (_12329_, _12328_, _05375_);
  and (_12330_, _12327_, _12315_);
  and (_12332_, _12330_, _05911_);
  nor (_12333_, _12332_, _12329_);
  and (_12334_, _12333_, _05793_);
  and (_12336_, _12334_, _12273_);
  and (_12337_, _12336_, _12230_);
  and (_12338_, _12337_, _12082_);
  and (_12339_, _05460_, _05335_);
  nand (_12340_, _12339_, _12338_);
  and (_12341_, _12340_, _12184_);
  and (_12343_, _12341_, _12088_);
  and (_12344_, _12156_, _06873_);
  and (_12345_, _12344_, _06610_);
  not (_12346_, _07470_);
  and (_12347_, _07105_, _06870_);
  and (_12349_, _12347_, _12346_);
  and (_12350_, _06870_, _06451_);
  nand (_12351_, _12350_, _07038_);
  nor (_12352_, _12347_, _11309_);
  and (_12353_, _12352_, _12351_);
  not (_12354_, _06828_);
  nand (_12355_, _12135_, _12354_);
  and (_12356_, _12355_, _06873_);
  nor (_12357_, _12356_, _12097_);
  and (_12358_, _12357_, _12353_);
  nor (_12360_, _11283_, _06828_);
  and (_12361_, _12360_, _12159_);
  and (_12362_, _12361_, _12096_);
  and (_12363_, _12362_, _12137_);
  nor (_12364_, _12363_, _12094_);
  nor (_12365_, _12344_, _12091_);
  not (_12367_, _12365_);
  nor (_12368_, _12367_, _12364_);
  and (_12369_, _12368_, _12358_);
  and (_12370_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_12371_, _12364_);
  and (_12373_, _12358_, _12367_);
  and (_12374_, _12373_, _12371_);
  and (_12376_, \oc8051_top_1.oc8051_memory_interface1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_12377_, _12376_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_12378_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12379_, _12378_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_12380_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_12381_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_12382_, _12381_, _12380_);
  and (_12384_, _12382_, _12379_);
  and (_12385_, _12384_, _12377_);
  and (_12386_, _12385_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_12387_, _12385_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_12389_, _12387_, _12386_);
  and (_12390_, _12389_, _12374_);
  not (_12392_, _11309_);
  nor (_12393_, _12392_, _06668_);
  or (_12394_, _12393_, _12390_);
  or (_12395_, _12394_, _12370_);
  or (_12396_, _12395_, _12349_);
  nor (_12397_, _12396_, _12345_);
  nand (_12399_, _12397_, _12343_);
  and (_12400_, _12358_, _12014_);
  nand (_12401_, _12357_, _12353_);
  and (_12402_, _12401_, _07176_);
  nor (_12403_, _12402_, _12400_);
  not (_12404_, _12403_);
  and (_12405_, _12403_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_12406_, _12358_, _12067_);
  and (_12407_, _12401_, _07582_);
  nor (_12408_, _12407_, _12406_);
  and (_12409_, _12408_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_12410_, _12403_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_12411_, _12410_, _12405_);
  and (_12412_, _12411_, _12409_);
  or (_12413_, _12412_, _12405_);
  nor (_12414_, _12408_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_12415_, _12414_, _12409_);
  and (_12416_, _12415_, _12411_);
  not (_12417_, _07507_);
  or (_12418_, _12401_, _12417_);
  nor (_12419_, _05474_, _05578_);
  and (_12420_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12421_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_12422_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_12423_, _12422_, _12421_);
  and (_12424_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_12425_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_12426_, _12425_, _12424_);
  and (_12427_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_12428_, _06251_, _06207_);
  nor (_12429_, _12428_, _12427_);
  and (_12430_, _12429_, _12426_);
  and (_12431_, _12430_, _12423_);
  nor (_12432_, _12431_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12433_, _12432_, _12420_);
  nor (_12434_, _12433_, _06200_);
  nor (_12435_, _12434_, _12419_);
  not (_12436_, _12435_);
  or (_12437_, _12436_, _12358_);
  nand (_12438_, _12437_, _12418_);
  or (_12439_, _12438_, _05583_);
  and (_12440_, _12358_, _07490_);
  nor (_12441_, _05474_, _05117_);
  and (_12442_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12443_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_12444_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_12445_, _12444_, _12443_);
  and (_12446_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_12447_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_12448_, _12447_, _12446_);
  and (_12449_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  not (_12450_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_12451_, _06251_, _12450_);
  nor (_12452_, _12451_, _12449_);
  and (_12453_, _12452_, _12448_);
  and (_12454_, _12453_, _12445_);
  nor (_12455_, _12454_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12456_, _12455_, _12442_);
  nor (_12457_, _12456_, _06200_);
  nor (_12458_, _12457_, _12441_);
  and (_12459_, _12458_, _12401_);
  nor (_12460_, _12459_, _12440_);
  and (_12461_, _12460_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_12462_, _12438_, _05583_);
  and (_12463_, _12462_, _12439_);
  nand (_12464_, _12463_, _12461_);
  nand (_12465_, _12464_, _12439_);
  and (_12466_, _12465_, _12416_);
  or (_12467_, _12466_, _12413_);
  and (_12468_, _12358_, _07470_);
  and (_12469_, _12401_, _07561_);
  nor (_12470_, _12469_, _12468_);
  nor (_12471_, _12470_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12472_, _12470_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_12473_, _07454_);
  or (_12474_, _12401_, _12473_);
  not (_12475_, _07543_);
  or (_12476_, _12358_, _12475_);
  nand (_12477_, _12476_, _12474_);
  or (_12478_, _12477_, _05220_);
  not (_12479_, _12478_);
  not (_12480_, _07439_);
  or (_12481_, _12401_, _12480_);
  not (_12482_, _07525_);
  or (_12483_, _12358_, _12482_);
  and (_12484_, _12483_, _12481_);
  nand (_12485_, _12484_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_12486_, _12313_);
  or (_12487_, _12401_, _12486_);
  nor (_12488_, _05474_, _05236_);
  and (_12489_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_12490_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_12491_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_12492_, _12491_, _12490_);
  and (_12493_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  not (_12494_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_12495_, _06251_, _12494_);
  nor (_12496_, _12495_, _12493_);
  and (_12497_, _12496_, _12492_);
  and (_12498_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_12499_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_12500_, _12499_, _12498_);
  and (_12501_, _12500_, _12497_);
  nor (_12502_, _12501_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12503_, _12502_, _12489_);
  nor (_12504_, _12503_, _06200_);
  nor (_12505_, _12504_, _12488_);
  not (_12507_, _12505_);
  or (_12508_, _12507_, _12358_);
  and (_12509_, _12508_, _12487_);
  and (_12510_, _12509_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_12512_, _12484_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_12513_, _12512_, _12485_);
  and (_12514_, _12513_, _12510_);
  not (_12515_, _12514_);
  nand (_12516_, _12515_, _12485_);
  nand (_12517_, _12477_, _05220_);
  and (_12518_, _12517_, _12478_);
  and (_12519_, _12518_, _12516_);
  or (_12520_, _12519_, _12479_);
  nor (_12521_, _12520_, _12472_);
  nor (_12522_, _12521_, _12471_);
  nor (_12523_, _12460_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_12524_, _12523_, _12461_);
  and (_12525_, _12463_, _12524_);
  and (_12526_, _12525_, _12416_);
  and (_12527_, _12526_, _12522_);
  or (_12528_, _12527_, _12467_);
  or (_12529_, _12528_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_12530_, _12529_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_12531_, _12530_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_12532_, _12531_, _12404_);
  and (_12533_, _12528_, _12377_);
  nor (_12534_, _12533_, _12403_);
  or (_12535_, _12534_, _12532_);
  nand (_12536_, _12535_, _05195_);
  or (_12537_, _12535_, _05195_);
  and (_12538_, _12537_, _12536_);
  and (_12539_, _12351_, _12371_);
  nor (_12540_, _12539_, _12373_);
  and (_12541_, _12540_, _12538_);
  or (_12542_, _12541_, _12399_);
  not (_12543_, _06205_);
  and (_12544_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_12545_, _12544_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_12546_, _12545_, _12543_);
  and (_12547_, _12546_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12548_, _12547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12549_, _12548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_12550_, _12549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12551_, _12550_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_12552_, _12551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_12553_, _12552_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_12554_, _12552_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_12555_, _12554_, _12553_);
  or (_12556_, _12555_, _12343_);
  and (_12557_, _12556_, _05110_);
  and (_10697_, _12557_, _12542_);
  nand (_12558_, _11239_, _05841_);
  and (_12559_, _11222_, _11202_);
  and (_12560_, _12559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_12561_, _12559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_12562_, _12561_, _12560_);
  and (_12563_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_12564_, _12563_, _11202_);
  and (_12565_, _12564_, _11223_);
  or (_12566_, _12565_, _11193_);
  or (_12567_, _12566_, _12562_);
  nor (_12568_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_12569_, _12568_, _11234_);
  and (_12570_, _12569_, _12567_);
  and (_12571_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_12572_, _12571_, _11239_);
  or (_12573_, _12572_, _12570_);
  and (_12574_, _12573_, _05110_);
  and (_10705_, _12574_, _12558_);
  nor (_12575_, _11712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_12576_, _12575_, _12559_);
  and (_12577_, _11606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_12578_, _12577_, _11223_);
  or (_12579_, _12578_, _11193_);
  or (_12580_, _12579_, _12576_);
  or (_12581_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_12583_, _12581_, _11584_);
  and (_12584_, _12583_, _12580_);
  and (_12585_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_12586_, _12585_, _12584_);
  nor (_12587_, _11240_, _06054_);
  or (_12588_, _12587_, _12586_);
  and (_10709_, _12588_, _05110_);
  and (_10712_, _11998_, _05110_);
  nor (_10714_, _11783_, rst);
  and (_12589_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_12590_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or (_12591_, _12590_, _12589_);
  and (_10717_, _12591_, _05110_);
  or (_12592_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not (_12594_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_12595_, _06205_, _12594_);
  and (_12596_, _12595_, _05110_);
  and (_10720_, _12596_, _12592_);
  or (_12597_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_12598_, _06205_, _12494_);
  and (_12599_, _12598_, _05110_);
  and (_10724_, _12599_, _12597_);
  and (_12601_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_12602_, _12601_, _11202_);
  and (_12603_, _12602_, _11223_);
  and (_12604_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_12605_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_12606_, _12605_, _11193_);
  or (_12607_, _12606_, _12604_);
  or (_12608_, _12607_, _12603_);
  nor (_12609_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor (_12610_, _12609_, _11234_);
  and (_12611_, _12610_, _12608_);
  not (_12612_, _11234_);
  nor (_12613_, _12612_, _06229_);
  or (_12615_, _12613_, _11239_);
  or (_12616_, _12615_, _12611_);
  or (_12617_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_12618_, _12617_, _05110_);
  and (_10730_, _12618_, _12616_);
  nor (_12619_, _12612_, _05841_);
  and (_12620_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_12621_, _12620_, _11202_);
  and (_12622_, _12621_, _11223_);
  nand (_12623_, _11214_, _11202_);
  nor (_12624_, _12623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_12625_, _12623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_12626_, _12625_, _11193_);
  or (_12627_, _12626_, _12624_);
  or (_12628_, _12627_, _12622_);
  nor (_12629_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_12630_, _12629_, _11234_);
  and (_12631_, _12630_, _12628_);
  or (_12632_, _12631_, _11239_);
  or (_12633_, _12632_, _12619_);
  or (_12634_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_12635_, _12634_, _05110_);
  and (_10736_, _12635_, _12633_);
  and (_12636_, _06024_, _05376_);
  and (_12637_, _12636_, _06888_);
  and (_12638_, _12637_, _05806_);
  not (_12639_, _12638_);
  or (_12640_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_12641_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_12642_, _12641_, _11202_);
  and (_12643_, _12642_, _11223_);
  and (_12645_, _11213_, _11202_);
  or (_12646_, _12645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_12647_, _12646_, _12623_);
  or (_12648_, _12647_, _11193_);
  or (_12649_, _12648_, _12643_);
  and (_12650_, _12649_, _12640_);
  and (_12651_, _12650_, _12639_);
  nor (_12652_, _12612_, _06054_);
  or (_12653_, _12652_, _12651_);
  or (_12654_, _12653_, _11239_);
  or (_12655_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_12656_, _12655_, _05110_);
  and (_10739_, _12656_, _12654_);
  or (_12657_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12658_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12659_, _12658_, _11202_);
  and (_12660_, _12659_, _11223_);
  and (_12661_, _11212_, _11202_);
  nor (_12662_, _12661_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_12663_, _12662_, _12645_);
  or (_12664_, _12663_, _11193_);
  or (_12665_, _12664_, _12660_);
  and (_12666_, _12665_, _12657_);
  and (_12667_, _12666_, _12639_);
  nor (_12668_, _12639_, _05334_);
  or (_12669_, _12668_, _12667_);
  or (_12670_, _12669_, _11239_);
  or (_12671_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_12672_, _12671_, _05110_);
  and (_10746_, _12672_, _12670_);
  and (_12673_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_12674_, _12673_, _11202_);
  and (_12675_, _12674_, _11223_);
  and (_12676_, _11211_, _11202_);
  nor (_12677_, _12676_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_12678_, _12677_, _12661_);
  or (_12679_, _12678_, _11193_);
  or (_12680_, _12679_, _12675_);
  nor (_12681_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor (_12682_, _12681_, _11234_);
  and (_12683_, _12682_, _12680_);
  nor (_12684_, _12612_, _06088_);
  or (_12686_, _12684_, _11239_);
  or (_12687_, _12686_, _12683_);
  or (_12688_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_12689_, _12688_, _05110_);
  and (_10755_, _12689_, _12687_);
  and (_12690_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _05110_);
  and (_12691_, _12690_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_12692_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_12693_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_12694_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_12695_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_12696_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_12697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_12698_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_12699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_12700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12701_, _11661_, _12700_);
  and (_12702_, _12701_, _12699_);
  and (_12703_, _12702_, _12698_);
  and (_12704_, _12703_, _11657_);
  and (_12705_, _12704_, _12697_);
  and (_12706_, _12705_, _12696_);
  and (_12707_, _12706_, _12695_);
  and (_12708_, _12707_, _12694_);
  and (_12709_, _12708_, _12693_);
  nor (_12710_, _12709_, _12692_);
  and (_12711_, _12709_, _12692_);
  nor (_12712_, _12711_, _12710_);
  not (_12713_, _12712_);
  nor (_12714_, _12708_, _12693_);
  nor (_12715_, _12714_, _12709_);
  nor (_12716_, _12707_, _12694_);
  or (_12717_, _12716_, _12708_);
  nor (_12718_, _12706_, _12695_);
  nor (_12719_, _12718_, _12707_);
  nor (_12720_, _12705_, _12696_);
  nor (_12722_, _12720_, _12706_);
  not (_12723_, _12722_);
  nor (_12724_, _12704_, _12697_);
  nor (_12725_, _12724_, _12705_);
  not (_12726_, _12725_);
  not (_12727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_12728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12729_, _12702_, _11657_);
  and (_12730_, _12729_, _12728_);
  nor (_12731_, _12730_, _12727_);
  or (_12732_, _12731_, _12704_);
  and (_12733_, _12701_, _11657_);
  nor (_12734_, _12733_, _12699_);
  nor (_12735_, _12734_, _12729_);
  not (_12736_, _12735_);
  nor (_12737_, _11662_, _12700_);
  or (_12738_, _12737_, _12733_);
  and (_12739_, _12738_, _11696_);
  and (_12740_, _12739_, _12736_);
  nor (_12741_, _12729_, _12728_);
  or (_12742_, _12741_, _12730_);
  and (_12743_, _12742_, _12740_);
  and (_12744_, _12743_, _12732_);
  and (_12745_, _12744_, _12726_);
  and (_12747_, _12745_, _12723_);
  not (_12748_, _12747_);
  nor (_12749_, _12748_, _12719_);
  nand (_12750_, _12749_, _12717_);
  or (_12751_, _12750_, _12715_);
  nor (_12752_, _12751_, _12713_);
  and (_12753_, _12751_, _12713_);
  or (_12754_, _12753_, _12752_);
  or (_12755_, _12754_, _07437_);
  or (_12756_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_12757_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_12758_, _12757_, _12756_);
  and (_12759_, _12758_, _12755_);
  or (_10784_, _12759_, _12691_);
  and (_12760_, _12344_, _06984_);
  nor (_12761_, _12392_, _07028_);
  not (_12762_, _12014_);
  and (_12763_, _12347_, _12762_);
  and (_12764_, _12386_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_12765_, _12764_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_12766_, _12765_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_12767_, _12766_, _05496_);
  or (_12768_, _12766_, _05496_);
  and (_12769_, _12768_, _12767_);
  and (_12770_, _12769_, _12374_);
  and (_12771_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_12772_, _12771_, _12770_);
  or (_12773_, _12772_, _12763_);
  or (_12775_, _12773_, _12761_);
  nor (_12776_, _12775_, _12760_);
  nand (_12777_, _12776_, _12343_);
  and (_12778_, _12531_, _05195_);
  nor (_12779_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_12780_, _12779_, _12778_);
  nand (_12782_, _12780_, _05613_);
  and (_12783_, _12782_, _12403_);
  and (_12784_, _12533_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_12785_, _12784_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_12786_, _12785_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_12787_, _12786_, _05613_);
  and (_12788_, _12787_, _12404_);
  or (_12789_, _12788_, _12783_);
  nand (_12790_, _12789_, _05496_);
  or (_12791_, _12789_, _05496_);
  and (_12792_, _12791_, _12790_);
  and (_12793_, _12792_, _12540_);
  or (_12794_, _12793_, _12777_);
  and (_12795_, _12545_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12796_, _12795_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12797_, _12796_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_12798_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_12799_, _12798_, _12797_);
  nand (_12800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_12801_, _12800_, _06205_);
  and (_12802_, _12801_, _12799_);
  and (_12803_, _12802_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_12804_, _12803_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_12805_, _12804_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_12806_, _12805_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_12807_, _12805_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_12808_, _12807_, _12806_);
  or (_12809_, _12808_, _12343_);
  and (_12810_, _12809_, _05110_);
  and (_10789_, _12810_, _12794_);
  and (_10803_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _05110_);
  nor (_12811_, _11309_, rst);
  and (_10813_, _12811_, _12343_);
  and (_12812_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_12813_, _06229_, _06000_);
  and (_12814_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_12815_, _12814_, _12813_);
  and (_12816_, _12815_, _05337_);
  or (_12817_, _12816_, _12812_);
  and (_10862_, _12817_, _05110_);
  and (_12818_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_12819_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or (_12820_, _12819_, _12818_);
  and (_10880_, _12820_, _05110_);
  or (_12821_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_12822_, _06205_, _07514_);
  and (_12823_, _12822_, _05110_);
  and (_10883_, _12823_, _12821_);
  and (_12824_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_12825_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or (_12826_, _12825_, _12824_);
  and (_10935_, _12826_, _05110_);
  and (_12827_, _08287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_12828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_12829_, _08280_, _12828_);
  nor (_12830_, _12829_, _08287_);
  or (_12831_, _12830_, _12827_);
  nor (_12832_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_12833_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_12834_, _12833_, _12832_);
  nor (_12835_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_12836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_12837_, _12836_, _12835_);
  and (_12838_, _12837_, _12834_);
  nor (_12839_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_12841_, _12839_, _12838_);
  and (_12843_, _12841_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_12844_, _12843_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_12845_, _12844_, _08280_);
  nor (_12847_, _12845_, _12831_);
  nor (_12848_, _12847_, _08274_);
  nor (_12849_, _08236_, _06798_);
  and (_12850_, _12849_, _08274_);
  or (_12851_, _12850_, _12848_);
  and (_10942_, _12851_, _05110_);
  and (_12853_, _08297_, _06194_);
  and (_12854_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_12855_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_12856_, _12855_, _12854_);
  nor (_12857_, _12856_, _08274_);
  and (_12858_, _08276_, _06230_);
  or (_12859_, _12858_, _12857_);
  or (_12860_, _12859_, _12853_);
  and (_10966_, _12860_, _05110_);
  and (_12861_, _08297_, _06230_);
  and (_12862_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_12863_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_12864_, _12863_, _12862_);
  nor (_12865_, _12864_, _08274_);
  and (_12866_, _08276_, _06559_);
  or (_12867_, _12866_, _12865_);
  or (_12868_, _12867_, _12861_);
  and (_10974_, _12868_, _05110_);
  nor (_10979_, _12313_, rst);
  and (_12869_, _08297_, _06183_);
  and (_12870_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_12871_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_12872_, _12871_, _12870_);
  nor (_12873_, _12872_, _08274_);
  not (_12874_, _05334_);
  and (_12875_, _08276_, _12874_);
  or (_12876_, _12875_, _12873_);
  or (_12877_, _12876_, _12869_);
  and (_10985_, _12877_, _05110_);
  and (_12878_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_12879_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_12880_, pc_log_change, _12879_);
  or (_12881_, _12880_, _12878_);
  and (_11004_, _12881_, _05110_);
  and (_12882_, _08297_, _12874_);
  and (_12883_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_12884_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_12885_, _12884_, _12883_);
  nor (_12887_, _12885_, _08274_);
  and (_12888_, _08276_, _06194_);
  or (_12889_, _12888_, _12887_);
  or (_12890_, _12889_, _12882_);
  and (_11006_, _12890_, _05110_);
  nand (_12891_, _11280_, _07418_);
  or (_12892_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_12893_, _12892_, _05110_);
  and (_11058_, _12893_, _12891_);
  not (_12894_, _05901_);
  and (_12895_, _08297_, _12894_);
  and (_12896_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_12897_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_12898_, _12897_, _12896_);
  nor (_12899_, _12898_, _08274_);
  and (_12900_, _08276_, _08224_);
  or (_12901_, _12900_, _12899_);
  or (_12902_, _12901_, _12895_);
  and (_11073_, _12902_, _05110_);
  and (_12903_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not (_12904_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_12905_, _06205_, _12904_);
  or (_12906_, _12905_, _12903_);
  and (_11095_, _12906_, _05110_);
  and (_12907_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not (_12908_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_12909_, _06205_, _12908_);
  or (_12910_, _12909_, _12907_);
  and (_11112_, _12910_, _05110_);
  and (_12911_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_12912_, _06205_, _07571_);
  or (_12913_, _12912_, _12911_);
  and (_11115_, _12913_, _05110_);
  and (_12914_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_12915_, _06205_, _07514_);
  or (_12916_, _12915_, _12914_);
  and (_11121_, _12916_, _05110_);
  and (_11126_, _11576_, _05110_);
  not (_12917_, _06895_);
  or (_12918_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  not (_12919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_12920_, _08884_, _12919_);
  and (_12921_, _12920_, _12918_);
  and (_12922_, _12921_, _12917_);
  nor (_12923_, _12917_, _06088_);
  or (_12924_, _12923_, _12922_);
  and (_11138_, _12924_, _05110_);
  or (_12925_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_12926_, _06205_, _12297_);
  and (_12927_, _12926_, _05110_);
  and (_11148_, _12927_, _12925_);
  or (_12928_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_12929_, _06205_, _06330_);
  and (_12930_, _12929_, _05110_);
  and (_11150_, _12930_, _12928_);
  or (_12931_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_12932_, _06205_, _07474_);
  and (_12933_, _12932_, _05110_);
  and (_11154_, _12933_, _12931_);
  and (_12934_, _08297_, _08224_);
  and (_12935_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_12936_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_12937_, _12936_, _12935_);
  nor (_12938_, _12937_, _08274_);
  and (_12939_, _08276_, _06183_);
  or (_12940_, _12939_, _12938_);
  or (_12942_, _12940_, _12934_);
  and (_11161_, _12942_, _05110_);
  and (_12943_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_12944_, _12738_, _11696_);
  nor (_12946_, _12944_, _12739_);
  or (_12947_, _12946_, _07437_);
  or (_12948_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_12949_, _12948_, _11510_);
  and (_12950_, _12949_, _12947_);
  or (_12952_, _12950_, _12943_);
  and (_11164_, _12952_, _05110_);
  and (_12953_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_12954_, _12743_, _12732_);
  nor (_12955_, _12954_, _12744_);
  or (_12956_, _12955_, _07437_);
  or (_12957_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_12958_, _12957_, _11510_);
  and (_12959_, _12958_, _12956_);
  or (_12960_, _12959_, _12953_);
  and (_11195_, _12960_, _05110_);
  or (_12961_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_12962_, _06205_, _07532_);
  and (_12963_, _12962_, _05110_);
  and (_11198_, _12963_, _12961_);
  nor (_12964_, _12742_, _12740_);
  nor (_12965_, _12964_, _12743_);
  or (_12966_, _12965_, _07437_);
  or (_12967_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_12968_, _12967_, _11510_);
  and (_12969_, _12968_, _12966_);
  and (_12970_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_12971_, _12970_, _12969_);
  and (_11201_, _12971_, _05110_);
  and (_12972_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_12973_, _12739_, _12736_);
  nor (_12974_, _12973_, _12740_);
  or (_12975_, _12974_, _07437_);
  or (_12976_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_12977_, _12976_, _11510_);
  and (_12978_, _12977_, _12975_);
  or (_12979_, _12978_, _12972_);
  and (_11210_, _12979_, _05110_);
  or (_12980_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_12981_, _06205_, _06352_);
  and (_12982_, _12981_, _05110_);
  and (_11221_, _12982_, _12980_);
  and (_12983_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not (_12984_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_12985_, _06205_, _12984_);
  or (_12986_, _12985_, _12983_);
  and (_11224_, _12986_, _05110_);
  and (_12987_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_12988_, _06205_, _07532_);
  or (_12989_, _12988_, _12987_);
  and (_11229_, _12989_, _05110_);
  or (_12990_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_12991_, _06205_, _07425_);
  and (_12992_, _12991_, _05110_);
  and (_11244_, _12992_, _12990_);
  or (_12993_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_12994_, _06205_, _06370_);
  and (_12995_, _12994_, _05110_);
  and (_11267_, _12995_, _12993_);
  and (_12996_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_12997_, _06205_, _07553_);
  or (_12998_, _12997_, _12996_);
  and (_11270_, _12998_, _05110_);
  or (_12999_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_13000_, _06205_, _07494_);
  and (_13001_, _13000_, _05110_);
  and (_11278_, _13001_, _12999_);
  nand (_13002_, _11280_, _06512_);
  or (_13003_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_13004_, _13003_, _05110_);
  and (_11285_, _13004_, _13002_);
  or (_13005_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_13006_, _06205_, _06397_);
  and (_13007_, _13006_, _05110_);
  and (_11291_, _13007_, _13005_);
  or (_13008_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_13009_, _06205_, _07457_);
  and (_13010_, _13009_, _05110_);
  and (_11318_, _13010_, _13008_);
  or (_13011_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_13012_, _06205_, _07442_);
  and (_13013_, _13012_, _05110_);
  and (_11352_, _13013_, _13011_);
  or (_13014_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_13015_, _06205_, _06248_);
  and (_13016_, _13015_, _05110_);
  and (_11361_, _13016_, _13014_);
  or (_13017_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_13018_, _06205_, _06413_);
  and (_13019_, _13018_, _05110_);
  and (_11364_, _13019_, _13017_);
  or (_13020_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_13021_, _06205_, _06285_);
  and (_13023_, _13021_, _05110_);
  and (_11375_, _13023_, _13020_);
  or (_13024_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_13025_, _06205_, _06307_);
  and (_13026_, _13025_, _05110_);
  and (_11390_, _13026_, _13024_);
  and (_13028_, _06177_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_13029_, _06184_, _12894_);
  or (_13030_, _13029_, _13028_);
  and (_11392_, _13030_, _05110_);
  or (_13031_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_13032_, _06205_, _12054_);
  and (_13033_, _13032_, _05110_);
  and (_11413_, _13033_, _13031_);
  and (_13034_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _07601_);
  and (_13035_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_13036_, _13035_, _13034_);
  and (_11496_, _13036_, _05110_);
  nor (_11509_, _11580_, rst);
  and (_11514_, _11570_, _05110_);
  and (_13037_, _07601_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_13038_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_13039_, _13038_, _13037_);
  and (_11522_, _13039_, _05110_);
  and (_13040_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07601_);
  and (_13041_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_13042_, _13041_, _13040_);
  and (_11531_, _13042_, _05110_);
  and (_13043_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07601_);
  and (_13044_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_13045_, _13044_, _13043_);
  and (_11534_, _13045_, _05110_);
  and (_13046_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_13047_, _06205_, _12494_);
  or (_13048_, _13047_, _13046_);
  and (_11624_, _13048_, _05110_);
  and (_13049_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_13050_, _06205_, _06207_);
  or (_13051_, _13050_, _13049_);
  and (_11643_, _13051_, _05110_);
  and (_13052_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_13053_, _06205_, _12450_);
  or (_13054_, _13053_, _13052_);
  and (_11649_, _13054_, _05110_);
  and (_13055_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_13056_, _06205_, _09467_);
  or (_13057_, _13056_, _13055_);
  and (_11659_, _13057_, _05110_);
  and (_13058_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_13059_, _06205_, _07167_);
  or (_13060_, _13059_, _13058_);
  and (_11663_, _13060_, _05110_);
  and (_13061_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_13062_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_13063_, _06205_, _13062_);
  or (_13064_, _13063_, _13061_);
  and (_11668_, _13064_, _05110_);
  and (_13065_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not (_13066_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_13067_, _06205_, _13066_);
  or (_13068_, _13067_, _13065_);
  and (_11674_, _13068_, _05110_);
  and (_13069_, _06807_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_13070_, _11728_, _07120_);
  or (_13071_, _13070_, _11732_);
  and (_13072_, _06463_, _06448_);
  and (_13073_, _11283_, _06342_);
  or (_13074_, _13073_, _13072_);
  or (_13075_, _13074_, _13071_);
  and (_13076_, _06849_, _06277_);
  or (_13077_, _12158_, _12138_);
  and (_13078_, _06856_, _06434_);
  and (_13079_, _07080_, _06451_);
  or (_13080_, _13079_, _13078_);
  or (_13081_, _13080_, _13077_);
  or (_13082_, _13081_, _13076_);
  or (_13083_, _13082_, _06940_);
  or (_13084_, _13083_, _13075_);
  and (_13085_, _13084_, _06842_);
  or (_11679_, _13085_, _13069_);
  and (_13086_, _06852_, _06276_);
  or (_13087_, _06451_, _06447_);
  nand (_13088_, _13087_, _13086_);
  and (_13089_, _13088_, _06858_);
  or (_13090_, _06849_, _06954_);
  or (_11694_, _13090_, _13089_);
  and (_13091_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not (_13092_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_13093_, _06205_, _13092_);
  or (_13094_, _13093_, _13091_);
  and (_11697_, _13094_, _05110_);
  and (_13095_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_13096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_13097_, pc_log_change, _13096_);
  or (_13098_, _13097_, _13095_);
  and (_11702_, _13098_, _05110_);
  and (_11704_, _11321_, _05110_);
  and (_13099_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_13100_, _06205_, _12594_);
  or (_13101_, _13100_, _13099_);
  and (_11707_, _13101_, _05110_);
  and (_13102_, _11412_, _06915_);
  and (_13103_, _11358_, _06926_);
  or (_13104_, _13103_, _11395_);
  nor (_13105_, _13104_, _13102_);
  nand (_13106_, _13105_, _11439_);
  or (_13107_, _13106_, _11459_);
  and (_13109_, _11387_, _11365_);
  and (_13110_, _11342_, _06922_);
  and (_13111_, _11345_, _06924_);
  or (_13112_, _13111_, _13110_);
  or (_13113_, _13112_, _13109_);
  or (_13114_, _11441_, _11427_);
  and (_13115_, _11412_, _11365_);
  or (_13116_, _13115_, _11476_);
  or (_13117_, _13116_, _13114_);
  or (_13118_, _13117_, _13113_);
  or (_13119_, _13118_, _13107_);
  or (_13120_, _13119_, _06933_);
  and (_13121_, _13120_, _05475_);
  nor (_13122_, _06908_, _06238_);
  or (_13123_, _13122_, rst);
  or (_11718_, _13123_, _13121_);
  and (_11725_, _11312_, _05110_);
  nor (_13124_, _11484_, _11482_);
  nor (_13125_, _13124_, _11485_);
  or (_13126_, _13125_, _06200_);
  or (_13127_, _05474_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_13128_, _13127_, _12757_);
  and (_11733_, _13128_, _13126_);
  and (_13129_, _11481_, _05474_);
  nand (_13130_, _13129_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_13131_, _13129_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_13132_, _13131_, _12757_);
  and (_11739_, _13132_, _13130_);
  nand (_13133_, _06673_, _06229_);
  or (_13134_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_13135_, _13134_, _05110_);
  and (_11913_, _13135_, _13133_);
  nand (_13136_, _11280_, _06668_);
  or (_13137_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_13138_, _13137_, _05110_);
  and (_11940_, _13138_, _13136_);
  nand (_13139_, _11280_, _07337_);
  or (_13140_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_13141_, _13140_, _05110_);
  and (_11947_, _13141_, _13139_);
  or (_13142_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand (_13143_, _06205_, _13062_);
  and (_13144_, _13143_, _05110_);
  and (_11980_, _13144_, _13142_);
  and (_13145_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_13146_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_13147_, _13146_, _13145_);
  nor (_13148_, _13147_, _08274_);
  or (_13149_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _11264_);
  and (_13150_, _13149_, _08236_);
  and (_13151_, _13150_, _08274_);
  or (_13152_, _13151_, _13148_);
  and (_11983_, _13152_, _05110_);
  or (_13153_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_13154_, _06205_, _07571_);
  and (_13156_, _13154_, _05110_);
  and (_11991_, _13156_, _13153_);
  and (_13157_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_13158_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_13159_, _13158_, _13157_);
  and (_12015_, _13159_, _05110_);
  and (_13160_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_13161_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or (_13162_, _13161_, _13160_);
  and (_12019_, _13162_, _05110_);
  and (_12047_, _11944_, _05110_);
  nor (_12055_, _12067_, rst);
  and (_13163_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_13164_, _13163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_12069_, _13164_, _05110_);
  and (_13165_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_13166_, _13165_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_12076_, _13166_, _05110_);
  and (_13167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _05110_);
  and (_13168_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05110_);
  and (_13170_, _13168_, _11505_);
  or (_12079_, _13170_, _13167_);
  nor (_12081_, _12435_, rst);
  and (_13171_, _08869_, _05804_);
  nand (_13172_, _13171_, _05841_);
  not (_13174_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_13175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13174_);
  not (_13176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_13177_, _13176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor (_13178_, _13177_, _13175_);
  and (_13179_, _11238_, _05804_);
  nor (_13180_, _13179_, _13178_);
  not (_13181_, _13180_);
  and (_13182_, _13181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  not (_13183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_13184_, t1_i);
  and (_13185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _13184_);
  nor (_13186_, _13185_, _13183_);
  not (_13187_, _13186_);
  not (_13188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_13189_, _13188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_13190_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_13191_, _13190_);
  and (_13192_, _13191_, _13189_);
  and (_13193_, _13192_, _13187_);
  and (_13194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_13195_, _13194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_13196_, _13195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_13197_, _13196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_13198_, _13197_, _13193_);
  and (_13199_, _13198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_13200_, _13199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_13201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_13202_, _13201_, _13198_);
  nor (_13203_, _13202_, _13200_);
  and (_13204_, _13180_, _13203_);
  and (_13205_, _13199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_13206_, _13205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_13207_, _13206_, _13175_);
  nand (_13208_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_13209_, _13208_, _13179_);
  or (_13210_, _13209_, _13204_);
  or (_13211_, _13210_, _13182_);
  or (_13212_, _13171_, _13211_);
  and (_13213_, _13212_, _05110_);
  and (_12085_, _13213_, _13172_);
  and (_13214_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_13215_, _13214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_12107_, _13215_, _05110_);
  and (_13216_, _13196_, _13193_);
  nor (_13217_, _13216_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_13218_, _13217_, _13198_);
  and (_13219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor (_13220_, _13219_, _13179_);
  and (_13221_, _13220_, _13218_);
  not (_13222_, _13220_);
  and (_13223_, _13222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_13224_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_13225_, _13224_, _13179_);
  or (_13226_, _13225_, _13223_);
  or (_13227_, _13226_, _13221_);
  or (_13228_, _13227_, _13171_);
  nand (_13229_, _13171_, _05334_);
  and (_13230_, _13229_, _05110_);
  and (_12110_, _13230_, _13228_);
  and (_13231_, _13195_, _13193_);
  nor (_13232_, _13231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_13233_, _13232_, _13216_);
  and (_13234_, _13233_, _13220_);
  and (_13235_, _13222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_13236_, _13235_, _13234_);
  nand (_13237_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_13238_, _13237_, _13179_);
  or (_13239_, _13238_, _13171_);
  or (_13240_, _13239_, _13236_);
  nand (_13241_, _13171_, _06088_);
  and (_13242_, _13241_, _05110_);
  and (_12113_, _13242_, _13240_);
  and (_13243_, _13193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_13244_, _13243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_13245_, _13244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_13246_, _13245_, _13231_);
  nand (_13247_, _13246_, _13220_);
  or (_13248_, _13220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_13249_, _13248_, _13247_);
  and (_13250_, _06894_, _05804_);
  and (_13251_, _13202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_13252_, _13251_, _13175_);
  nand (_13253_, _13252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_13254_, _13253_, _13179_);
  or (_13255_, _13254_, _13250_);
  or (_13256_, _13255_, _13249_);
  nand (_13257_, _13250_, _06229_);
  and (_13258_, _13257_, _05110_);
  and (_12116_, _13258_, _13256_);
  nand (_13259_, _13171_, _06054_);
  nand (_13260_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_13261_, _13260_, _13179_);
  nor (_13262_, _13198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_13263_, _13262_, _13199_);
  and (_13264_, _13263_, _13180_);
  and (_13265_, _13181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_13266_, _13265_, _13264_);
  or (_13267_, _13266_, _13261_);
  or (_13268_, _13267_, _13171_);
  and (_13269_, _13268_, _05110_);
  and (_12122_, _13269_, _13259_);
  or (_13270_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand (_13271_, _06205_, _12908_);
  and (_13272_, _13271_, _05110_);
  and (_12124_, _13272_, _13270_);
  and (_13273_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_13274_, _13273_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_12129_, _13274_, _05110_);
  not (_13275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_13276_, _13220_, _13275_);
  or (_13277_, _13193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_13278_, _13219_, _13243_);
  and (_13279_, _13175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_13280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_13281_, _13280_, _13201_);
  and (_13282_, _13281_, _13197_);
  and (_13283_, _13282_, _13279_);
  or (_13284_, _13283_, _13278_);
  nand (_13285_, _13284_, _13277_);
  nor (_13286_, _13285_, _13179_);
  or (_13287_, _13286_, _13250_);
  or (_13288_, _13287_, _13276_);
  nand (_13289_, _13250_, _06798_);
  and (_13290_, _13289_, _05110_);
  and (_12133_, _13290_, _13288_);
  nor (_13291_, _13243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_13292_, _13291_, _13244_);
  nand (_13294_, _13292_, _13220_);
  or (_13295_, _13220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_13296_, _13295_, _13294_);
  nand (_13297_, _13252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_13298_, _13297_, _13179_);
  or (_13299_, _13298_, _13250_);
  or (_13300_, _13299_, _13296_);
  nand (_13301_, _13250_, _05938_);
  and (_13302_, _13301_, _05110_);
  and (_12136_, _13302_, _13300_);
  and (_13303_, _12528_, _12376_);
  or (_13304_, _13303_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_13305_, _13304_, _12534_);
  and (_13306_, _12530_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_13308_, _13306_, _12531_);
  and (_13309_, _13308_, _12403_);
  or (_13310_, _13309_, _13305_);
  and (_13311_, _13310_, _12540_);
  and (_13312_, _12344_, _07305_);
  and (_13313_, _12374_, _06918_);
  and (_13314_, _12347_, _12473_);
  and (_13315_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_13316_, _12392_, _07337_);
  or (_13317_, _13316_, _13315_);
  or (_13318_, _13317_, _13314_);
  or (_13319_, _13318_, _13313_);
  nor (_13320_, _13319_, _13312_);
  nand (_13321_, _13320_, _12343_);
  or (_13322_, _13321_, _13311_);
  nor (_13323_, _12551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_13324_, _13323_, _12552_);
  or (_13325_, _13324_, _12343_);
  and (_13326_, _13325_, _05110_);
  and (_12139_, _13326_, _13322_);
  and (_13327_, _07038_, _06870_);
  and (_13328_, _13327_, _06451_);
  nor (_13329_, _13328_, _12364_);
  nor (_13330_, _13329_, _12373_);
  not (_13331_, _12461_);
  nand (_13332_, _12524_, _12522_);
  nand (_13333_, _13332_, _13331_);
  or (_13334_, _12463_, _13333_);
  nand (_13335_, _12463_, _13333_);
  and (_13336_, _13335_, _13334_);
  and (_13337_, _13336_, _13330_);
  and (_13338_, _12436_, _12347_);
  not (_13339_, _06548_);
  or (_13340_, _12369_, _12344_);
  and (_13341_, _13340_, _13339_);
  and (_13342_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_13343_, _12374_, _12417_);
  or (_13344_, _13343_, _13342_);
  or (_13345_, _13344_, _13341_);
  or (_13346_, _13345_, _13338_);
  or (_13348_, _13346_, _13337_);
  and (_13349_, _13348_, _12343_);
  nor (_13350_, _12546_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_13351_, _13350_, _12547_);
  nor (_13352_, _13351_, _12343_);
  or (_13353_, _13352_, _13349_);
  and (_12143_, _13353_, _05110_);
  nand (_13354_, _13179_, _06798_);
  not (_13355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_13356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_13358_, _13356_, _13198_);
  and (_13359_, _13251_, _13177_);
  nor (_13361_, _13359_, _13358_);
  nor (_13362_, _13361_, _13355_);
  and (_13363_, _13361_, _13355_);
  nor (_13364_, _13363_, _13362_);
  or (_13365_, _13364_, _13179_);
  and (_13366_, _13365_, _13354_);
  or (_13367_, _13366_, _13171_);
  nand (_13368_, _13171_, _13355_);
  and (_13369_, _13368_, _05110_);
  and (_12152_, _13369_, _13367_);
  nand (_13370_, _13179_, _05938_);
  not (_13371_, _13171_);
  nor (_13372_, _13362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_13373_, _13362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_13374_, _13373_, _13372_);
  or (_13375_, _13374_, _13179_);
  and (_13376_, _13375_, _13371_);
  and (_13377_, _13376_, _13370_);
  and (_13378_, _13250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_13379_, _13378_, _13377_);
  and (_12155_, _13379_, _05110_);
  nor (_13380_, _11693_, _11690_);
  nor (_13381_, _13380_, _11695_);
  or (_13382_, _13381_, _07437_);
  or (_13383_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_13384_, _13383_, _11510_);
  and (_13385_, _13384_, _13382_);
  and (_13386_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_13387_, _13386_, _13385_);
  and (_12157_, _13387_, _05110_);
  nand (_13388_, _13179_, _06088_);
  and (_13389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_13390_, _13389_, _13197_);
  and (_13391_, _13390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_13392_, _13391_, _13193_);
  and (_13393_, _13392_, _13356_);
  and (_13394_, _13282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_13395_, _13394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_13396_, _13395_, _13193_);
  and (_13397_, _13396_, _13177_);
  nor (_13398_, _13397_, _13393_);
  or (_13399_, _13398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_13400_, _13398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_13401_, _13400_, _13399_);
  nor (_13402_, _13401_, _13179_);
  nor (_13403_, _13402_, _13171_);
  and (_13404_, _13403_, _13388_);
  and (_13405_, _06062_, _05806_);
  and (_13406_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_13407_, _13406_, _13404_);
  and (_12161_, _13407_, _05110_);
  nand (_13408_, _13179_, _06054_);
  and (_13409_, _13197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_13410_, _13409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_13411_, _13410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_13412_, _13411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_13413_, _13412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_13414_, _13413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_13415_, _13414_, _13193_);
  and (_13416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_13417_, _13416_, _13415_);
  or (_13418_, _13417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_13419_, _13177_);
  and (_13420_, _13416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_13421_, _13420_, _13396_);
  nor (_13422_, _13421_, _13419_);
  and (_13423_, _13422_, _13418_);
  and (_13424_, _13416_, _13393_);
  or (_13425_, _13424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_13426_, _13420_, _13176_);
  nand (_13427_, _13426_, _13392_);
  and (_13428_, _13427_, _13419_);
  and (_13429_, _13428_, _13425_);
  or (_13430_, _13429_, _13423_);
  nor (_13431_, _13430_, _13179_);
  nor (_13432_, _13431_, _13171_);
  and (_00002_, _13432_, _13408_);
  and (_00003_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_00005_, _00003_, _00002_);
  and (_12164_, _00005_, _05110_);
  nand (_00006_, _13179_, _05334_);
  and (_00007_, _13415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00008_, _00007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_00009_, _00008_, _13177_);
  nor (_00010_, _00009_, _13417_);
  and (_00011_, _13392_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00012_, _00011_, _13176_);
  not (_00013_, _00012_);
  nor (_00014_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00015_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_00016_, _00015_, _00014_);
  and (_00017_, _00016_, _13419_);
  or (_00019_, _00017_, _00010_);
  or (_00020_, _00019_, _13179_);
  and (_00021_, _00020_, _13371_);
  and (_00022_, _00021_, _00006_);
  and (_00023_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_00024_, _00023_, _00022_);
  and (_12167_, _00024_, _05110_);
  or (_00025_, _13373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00026_, _00025_, _13398_);
  or (_00027_, _00026_, _13179_);
  nand (_00029_, _13179_, _06229_);
  nand (_00030_, _00029_, _00027_);
  or (_00032_, _00030_, _13405_);
  nand (_00033_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00034_, _00033_, _00032_);
  nor (_12170_, _00034_, rst);
  and (_00036_, _06473_, _05807_);
  not (_00037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_00039_, t0_i);
  and (_00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00039_);
  nor (_00041_, _00040_, _00037_);
  not (_00042_, _00041_);
  not (_00043_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_00044_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_00045_, _00044_, _00043_);
  and (_00046_, _00045_, _00042_);
  not (_00047_, _00046_);
  and (_00048_, _11233_, _05804_);
  nor (_00049_, _00048_, _00047_);
  or (_00050_, _00049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00051_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_00053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00054_, _00053_, _00052_);
  and (_00055_, _00054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_00056_, _00055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00057_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00058_, _00057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_00059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _00059_);
  and (_00061_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00062_, _00061_, _00058_);
  nand (_00063_, _00062_, _00051_);
  or (_00064_, _00063_, _00048_);
  and (_00065_, _00064_, _00050_);
  or (_00066_, _00065_, _00036_);
  nand (_00067_, _00036_, _06798_);
  and (_00068_, _00067_, _05110_);
  and (_12174_, _00068_, _00066_);
  not (_00069_, _00048_);
  or (_00070_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_00071_, _00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_00072_, _00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_00073_, _00072_, _00071_);
  and (_00074_, _00058_, _00046_);
  and (_00075_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00076_, _00075_, _00074_);
  or (_00077_, _00076_, _00073_);
  or (_00078_, _00077_, _00048_);
  and (_00079_, _00078_, _00070_);
  or (_00080_, _00079_, _00036_);
  nand (_00081_, _00036_, _05938_);
  and (_00082_, _00081_, _05110_);
  and (_12191_, _00082_, _00080_);
  nand (_00083_, _00036_, _06088_);
  and (_00084_, _00054_, _00046_);
  not (_00085_, _00084_);
  or (_00086_, _00085_, _00048_);
  and (_00087_, _00086_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_00088_, _00074_, _00060_);
  nand (_00089_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00090_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand (_00091_, _00090_, _00085_);
  and (_00092_, _00091_, _00089_);
  nor (_00093_, _00092_, _00048_);
  or (_00094_, _00093_, _00087_);
  or (_00095_, _00094_, _00036_);
  and (_00096_, _00095_, _05110_);
  and (_12196_, _00096_, _00083_);
  not (_00097_, _00036_);
  or (_00098_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00099_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_00100_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_00101_, _00100_, _00090_);
  or (_00102_, _00101_, _00099_);
  or (_00103_, _00102_, _00048_);
  and (_00104_, _00103_, _00098_);
  and (_00105_, _00104_, _00097_);
  nor (_00106_, _00097_, _06229_);
  or (_00107_, _00106_, _00105_);
  and (_12199_, _00107_, _05110_);
  nor (_00108_, _12744_, _12726_);
  nor (_00109_, _00108_, _12745_);
  or (_00110_, _00109_, _07437_);
  or (_00111_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00112_, _00111_, _12757_);
  and (_00113_, _00112_, _00110_);
  and (_00114_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _05110_);
  and (_00115_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_12202_, _00115_, _00113_);
  nand (_00116_, _08870_, _05334_);
  and (_00117_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_00118_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_00119_, _00118_, _00117_);
  or (_00120_, _00119_, _08870_);
  and (_00121_, _00120_, _05110_);
  and (_12206_, _00121_, _00116_);
  nand (_00122_, _08870_, _05841_);
  and (_00123_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_00124_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_00125_, _00124_, _00123_);
  or (_00126_, _00125_, _08870_);
  and (_00127_, _00126_, _05110_);
  and (_12218_, _00127_, _00122_);
  not (_00129_, _11219_);
  nor (_00130_, _11711_, _00129_);
  and (_00131_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_00132_, _00131_, _11223_);
  or (_00133_, _00132_, _00130_);
  and (_00134_, _00133_, _11202_);
  nor (_00135_, _11711_, _12919_);
  or (_00136_, _00135_, _11193_);
  or (_00137_, _00136_, _00134_);
  nor (_00138_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_00139_, _00138_, _11234_);
  and (_00140_, _00139_, _00137_);
  and (_00141_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_00142_, _00141_, _11239_);
  or (_00143_, _00142_, _00140_);
  nand (_00144_, _11239_, _06088_);
  and (_00145_, _00144_, _05110_);
  and (_12226_, _00145_, _00143_);
  nand (_00146_, _13179_, _05841_);
  not (_00147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00148_, _13428_, _00147_);
  not (_00149_, _00148_);
  nor (_00150_, _00149_, _13422_);
  nor (_00151_, _00150_, _00147_);
  and (_00152_, _13177_, _00147_);
  and (_00153_, _00152_, _13421_);
  nand (_00154_, _13420_, _13393_);
  nor (_00155_, _00154_, _00148_);
  or (_00156_, _00155_, _00153_);
  or (_00157_, _00156_, _00151_);
  or (_00158_, _00157_, _13179_);
  and (_00159_, _00158_, _13371_);
  and (_00160_, _00159_, _00146_);
  and (_00161_, _13250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_00162_, _00161_, _00160_);
  and (_12238_, _00162_, _05110_);
  nand (_00163_, _00036_, _06054_);
  and (_00164_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_00165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor (_00166_, _00165_, _00048_);
  and (_00167_, _00166_, _00164_);
  nand (_00168_, _00167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_00169_, _00167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00170_, _00169_, _00168_);
  nand (_00171_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_00172_, _00171_, _00048_);
  or (_00173_, _00172_, _00036_);
  or (_00174_, _00173_, _00170_);
  and (_00175_, _00174_, _05110_);
  and (_12244_, _00175_, _00163_);
  nand (_00176_, _00036_, _05841_);
  and (_00177_, _00164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_00178_, _00177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00179_, _00057_, _00046_);
  nor (_00180_, _00179_, _00165_);
  and (_00181_, _00180_, _00178_);
  and (_00182_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_00183_, _00182_, _00181_);
  nor (_00184_, _00183_, _00048_);
  not (_00185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_00186_, _00166_, _00185_);
  or (_00187_, _00186_, _00184_);
  or (_00188_, _00187_, _00036_);
  and (_00189_, _00188_, _05110_);
  and (_12247_, _00189_, _00176_);
  nand (_00190_, _00036_, _05334_);
  nor (_00191_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_00192_, _00191_, _00164_);
  and (_00193_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00194_, _00193_, _00192_);
  nor (_00195_, _00194_, _00048_);
  and (_00196_, _00048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_00197_, _00196_, _00195_);
  or (_00198_, _00197_, _00036_);
  and (_00199_, _00198_, _05110_);
  and (_12251_, _00199_, _00190_);
  and (_00200_, _11326_, _08272_);
  nand (_00201_, _00200_, _05872_);
  or (_00202_, _00200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_00203_, _00202_, _11330_);
  and (_00204_, _00203_, _00201_);
  nor (_00205_, _11330_, _05938_);
  or (_00206_, _00205_, _00204_);
  and (_12261_, _00206_, _05110_);
  or (_00207_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_00208_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_00209_, _00208_, _00207_);
  or (_00210_, _00209_, _06895_);
  nand (_00211_, _06895_, _05938_);
  and (_00212_, _00211_, _05110_);
  and (_12267_, _00212_, _00210_);
  or (_00213_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_00214_, _08884_, _11600_);
  and (_00215_, _00214_, _00213_);
  or (_00216_, _00215_, _06895_);
  nand (_00217_, _06895_, _06798_);
  and (_00218_, _00217_, _05110_);
  and (_12271_, _00218_, _00216_);
  nor (_00219_, _00069_, _05841_);
  and (_00220_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_00221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00222_, _00221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00223_, _00222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00224_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00225_, _00224_, _00220_);
  and (_00226_, _00225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00227_, _00226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_00228_, _00227_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00229_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00230_, _00226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00231_, _00230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00232_, _00231_, _00229_);
  and (_00233_, _00224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00234_, _00233_, _00055_);
  and (_00235_, _00234_, _00046_);
  or (_00236_, _00235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_00237_, _00165_);
  and (_00238_, _00235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_00239_, _00238_, _00237_);
  and (_00240_, _00239_, _00236_);
  and (_00241_, _00233_, _00074_);
  or (_00242_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_00243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00244_, _00243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00245_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_00246_, _00245_);
  and (_00247_, _00246_, _00244_);
  and (_00248_, _00247_, _00242_);
  or (_00249_, _00248_, _00240_);
  or (_00250_, _00249_, _00232_);
  and (_00251_, _00250_, _00069_);
  or (_00252_, _00251_, _00036_);
  or (_00254_, _00252_, _00219_);
  or (_00255_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00256_, _00255_, _05110_);
  and (_12293_, _00256_, _00254_);
  nand (_00257_, _00048_, _06054_);
  and (_00258_, _00074_, _00243_);
  and (_00259_, _00258_, _00224_);
  nand (_00260_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00261_, _00244_, _00060_);
  or (_00262_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00264_, _00262_, _00261_);
  and (_00265_, _00264_, _00260_);
  or (_00266_, _00225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00267_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_00268_, _00226_);
  and (_00269_, _00268_, _00267_);
  and (_00270_, _00269_, _00266_);
  and (_00271_, _00224_, _00164_);
  or (_00272_, _00271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00274_, _00233_, _00164_);
  nor (_00275_, _00274_, _00237_);
  and (_00276_, _00275_, _00272_);
  or (_00277_, _00276_, _00270_);
  or (_00278_, _00277_, _00265_);
  or (_00279_, _00278_, _00048_);
  and (_00280_, _00279_, _00257_);
  or (_00281_, _00280_, _00036_);
  or (_00282_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00283_, _00282_, _05110_);
  and (_12296_, _00283_, _00281_);
  nand (_00284_, _06890_, _05334_);
  and (_00285_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_00286_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_00287_, _00286_, _00285_);
  or (_00288_, _00287_, _06890_);
  and (_00289_, _00288_, _08871_);
  and (_00290_, _00289_, _00284_);
  and (_00291_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_00292_, _00291_, _00290_);
  and (_12299_, _00292_, _05110_);
  nand (_00293_, _06890_, _06088_);
  and (_00294_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_00295_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_00296_, _00295_, _00294_);
  or (_00297_, _00296_, _06890_);
  and (_00298_, _00297_, _08871_);
  and (_00299_, _00298_, _00293_);
  and (_00300_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_00301_, _00300_, _00299_);
  and (_12302_, _00301_, _05110_);
  nand (_00303_, _06890_, _06229_);
  and (_00304_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_00305_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_00307_, _00305_, _00304_);
  or (_00308_, _00307_, _06890_);
  and (_00309_, _00308_, _08871_);
  and (_00310_, _00309_, _00303_);
  and (_00311_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_00312_, _00311_, _00310_);
  and (_12306_, _00312_, _05110_);
  nand (_00313_, _06890_, _05938_);
  or (_00314_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_00315_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_00316_, _00315_, _00314_);
  or (_00317_, _00316_, _06890_);
  and (_00318_, _00317_, _08871_);
  and (_00319_, _00318_, _00313_);
  and (_00320_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_00321_, _00320_, _00319_);
  and (_12309_, _00321_, _05110_);
  not (_00322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_00323_, _00258_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00324_, _00323_, _00322_);
  nand (_00325_, _00258_, _00221_);
  and (_00326_, _00325_, _00261_);
  and (_00327_, _00326_, _00324_);
  and (_00328_, _00220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00329_, _00328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00330_, _00221_, _00220_);
  not (_00331_, _00330_);
  and (_00332_, _00331_, _00267_);
  and (_00333_, _00332_, _00329_);
  nand (_00334_, _00164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00335_, _00334_, _00322_);
  and (_00336_, _00221_, _00164_);
  nor (_00337_, _00336_, _00237_);
  and (_00338_, _00337_, _00335_);
  or (_00339_, _00338_, _00333_);
  or (_00340_, _00339_, _00327_);
  or (_00341_, _00340_, _00048_);
  nand (_00342_, _00048_, _05938_);
  and (_00343_, _00342_, _00341_);
  or (_00344_, _00343_, _00036_);
  nand (_00345_, _00036_, _00322_);
  and (_00346_, _00345_, _05110_);
  and (_12317_, _00346_, _00344_);
  nand (_00347_, _00048_, _06229_);
  or (_00348_, _00336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00349_, _00222_, _00164_);
  nor (_00350_, _00349_, _00237_);
  and (_00351_, _00350_, _00348_);
  and (_00352_, _00221_, _00074_);
  or (_00353_, _00352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_00354_, _00222_, _00074_);
  and (_00355_, _00354_, _00244_);
  and (_00356_, _00355_, _00353_);
  and (_00357_, _00222_, _00220_);
  nand (_00358_, _00357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00359_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_00360_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00361_, _00360_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00362_, _00361_, _00358_);
  or (_00363_, _00362_, _00356_);
  or (_00364_, _00363_, _00351_);
  or (_00365_, _00364_, _00048_);
  and (_00366_, _00365_, _00347_);
  or (_00367_, _00366_, _00036_);
  or (_00368_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00369_, _00368_, _05110_);
  and (_12320_, _00369_, _00367_);
  nand (_00370_, _00048_, _06088_);
  and (_00371_, _00258_, _00222_);
  or (_00372_, _00371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00373_, _00371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00374_, _00373_);
  and (_00375_, _00374_, _00261_);
  and (_00376_, _00375_, _00372_);
  and (_00378_, _00223_, _00220_);
  or (_00379_, _00357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_00380_, _00379_, _00267_);
  nor (_00381_, _00380_, _00378_);
  or (_00382_, _00349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00384_, _00223_, _00164_);
  nor (_00386_, _00384_, _00237_);
  and (_00388_, _00386_, _00382_);
  or (_00389_, _00388_, _00381_);
  or (_00390_, _00389_, _00376_);
  or (_00391_, _00390_, _00048_);
  and (_00392_, _00391_, _00370_);
  or (_00393_, _00392_, _00036_);
  or (_00394_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00396_, _00394_, _05110_);
  and (_12331_, _00396_, _00393_);
  nand (_00397_, _00048_, _05334_);
  or (_00398_, _00373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_00400_, _00259_);
  and (_00401_, _00400_, _00261_);
  and (_00402_, _00401_, _00398_);
  not (_00403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00404_, _00378_, _00403_);
  and (_00405_, _00378_, _00403_);
  or (_00406_, _00405_, _00404_);
  and (_00407_, _00406_, _00267_);
  or (_00408_, _00384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00409_, _00271_, _00237_);
  and (_00410_, _00409_, _00408_);
  or (_00412_, _00410_, _00407_);
  or (_00413_, _00412_, _00402_);
  or (_00414_, _00413_, _00048_);
  and (_00416_, _00414_, _00397_);
  or (_00418_, _00416_, _00036_);
  nand (_00420_, _00036_, _00403_);
  and (_00421_, _00420_, _05110_);
  and (_12335_, _00421_, _00418_);
  nand (_00423_, _06890_, _05841_);
  and (_00424_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_00425_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_00426_, _00425_, _00424_);
  or (_00427_, _00426_, _06890_);
  and (_00428_, _00427_, _08871_);
  and (_00429_, _00428_, _00423_);
  and (_00430_, _06895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_00431_, _00430_, _00429_);
  and (_12342_, _00431_, _05110_);
  or (_00432_, _00258_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00433_, _00323_, _00261_);
  and (_00434_, _00433_, _00432_);
  or (_00435_, _00220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not (_00436_, _00328_);
  and (_00437_, _00436_, _00267_);
  and (_00438_, _00437_, _00435_);
  or (_00439_, _00164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00440_, _00334_, _00165_);
  and (_00441_, _00440_, _00439_);
  or (_00442_, _00441_, _00438_);
  or (_00443_, _00442_, _00434_);
  or (_00444_, _00443_, _00048_);
  nand (_00445_, _00048_, _06798_);
  and (_00446_, _00445_, _00444_);
  or (_00447_, _00446_, _00036_);
  not (_00448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00449_, _00036_, _00448_);
  and (_00450_, _00449_, _05110_);
  and (_12348_, _00450_, _00447_);
  and (_00452_, _08273_, _05804_);
  nor (_00453_, _00452_, _00059_);
  and (_00454_, _00452_, _06799_);
  or (_00455_, _00454_, _00453_);
  and (_12359_, _00455_, _05110_);
  nand (_00456_, _00452_, _06229_);
  or (_00457_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00458_, _00457_, _05110_);
  and (_12366_, _00458_, _00456_);
  nand (_00459_, _00452_, _06088_);
  or (_00460_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_00461_, _00460_, _05110_);
  and (_12372_, _00461_, _00459_);
  nand (_00463_, _00452_, _05938_);
  or (_00464_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00465_, _00464_, _05110_);
  and (_12375_, _00465_, _00463_);
  nand (_00466_, _00452_, _06054_);
  or (_00468_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00469_, _00468_, _05110_);
  and (_12383_, _00469_, _00466_);
  nand (_00470_, _00452_, _05841_);
  or (_00471_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00473_, _00471_, _05110_);
  and (_12388_, _00473_, _00470_);
  nand (_00474_, _00452_, _05334_);
  or (_00475_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00476_, _00475_, _05110_);
  and (_12391_, _00476_, _00474_);
  nand (_00477_, _08276_, _05901_);
  or (_00478_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  or (_00479_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  and (_00480_, _00479_, _00478_);
  or (_00481_, _00480_, _08274_);
  and (_00482_, _00481_, _05110_);
  and (_12398_, _00482_, _00477_);
  and (_12506_, _11775_, _05110_);
  and (_00484_, _06856_, _06451_);
  not (_00485_, _00484_);
  and (_00486_, _06852_, _06446_);
  and (_00487_, _00486_, _07062_);
  nor (_00488_, _00487_, _06849_);
  and (_00489_, _00488_, _00485_);
  or (_12511_, _00489_, _06954_);
  and (_00490_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07601_);
  and (_00491_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00492_, _00491_, _00490_);
  and (_12582_, _00492_, _05110_);
  nor (_12593_, _12458_, rst);
  and (_00493_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07601_);
  and (_00494_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00495_, _00494_, _00493_);
  and (_12600_, _00495_, _05110_);
  and (_00496_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _05110_);
  and (_00497_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05110_);
  and (_00498_, _00497_, _11506_);
  or (_12644_, _00498_, _00496_);
  and (_00499_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_00500_, _00499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_12685_, _00500_, _05110_);
  and (_00501_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _07601_);
  and (_00502_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00503_, _00502_, _00501_);
  and (_12721_, _00503_, _05110_);
  nor (_12746_, _12505_, rst);
  and (_12774_, _12029_, _05110_);
  and (_12781_, _11890_, _05110_);
  nor (_12840_, _11866_, rst);
  or (_12842_, _12262_, rst);
  nand (_12846_, _12193_, _05110_);
  nand (_12852_, _12324_, _05110_);
  and (_00504_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_00505_, _06184_, _06559_);
  nand (_00506_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_00507_, _00506_, _06171_);
  or (_00508_, _00507_, _00505_);
  or (_00509_, _00508_, _00504_);
  and (_12941_, _00509_, _05110_);
  nand (_00510_, _08257_, _05938_);
  or (_00511_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_00512_, _00511_, _05110_);
  and (_12951_, _00512_, _00510_);
  and (_00513_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_00514_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_00515_, pc_log_change, _00514_);
  or (_00516_, _00515_, _00513_);
  and (_13022_, _00516_, _05110_);
  or (_00517_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_00518_, pc_log_change, _05496_);
  and (_00519_, _00518_, _05110_);
  and (_13027_, _00519_, _00517_);
  and (_13155_, _10472_, _11834_);
  and (_00520_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_00521_, _07034_, _06169_);
  or (_00522_, _00521_, _00520_);
  and (_13169_, _00522_, _05110_);
  and (_00523_, _10154_, _06626_);
  and (_00524_, _00523_, _05488_);
  nand (_00525_, _00524_, _05872_);
  or (_00526_, _00524_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00527_, _00526_, _05794_);
  and (_00528_, _00527_, _00525_);
  not (_00529_, _05793_);
  and (_00530_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00531_, _00523_, _05805_);
  nand (_00532_, _00531_, _06780_);
  or (_00533_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00534_, _00533_, _05806_);
  and (_00535_, _00534_, _00532_);
  or (_00536_, _00535_, _00530_);
  or (_00537_, _00536_, _00528_);
  and (_13293_, _00537_, _05110_);
  and (_00538_, _00523_, _08133_);
  nand (_00539_, _00538_, _05872_);
  or (_00540_, _00538_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_00541_, _00540_, _05794_);
  and (_00542_, _00541_, _00539_);
  and (_00543_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_00544_, _00531_, _06548_);
  or (_00545_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_00546_, _00545_, _05806_);
  and (_00547_, _00546_, _00544_);
  or (_00548_, _00547_, _00543_);
  or (_00549_, _00548_, _00542_);
  and (_13307_, _00549_, _05110_);
  not (_00550_, _00531_);
  or (_00551_, _00550_, _05782_);
  or (_00552_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00553_, _00552_, _05794_);
  and (_00554_, _00553_, _00551_);
  and (_00555_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_00556_, _00531_, _07418_);
  and (_00557_, _00556_, _05806_);
  and (_00558_, _00557_, _00552_);
  or (_00559_, _00558_, _00555_);
  or (_00560_, _00559_, _00554_);
  and (_13347_, _00560_, _05110_);
  and (_00561_, _00523_, _06632_);
  nand (_00562_, _00523_, _05401_);
  or (_00563_, _00562_, _11548_);
  and (_00564_, _00563_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00565_, _00564_, _00561_);
  and (_00566_, _00565_, _05794_);
  and (_00567_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_00568_, _00531_, _06668_);
  or (_00569_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00570_, _00569_, _05806_);
  and (_00571_, _00570_, _00568_);
  or (_00572_, _00571_, _00567_);
  or (_00573_, _00572_, _00566_);
  and (_13357_, _00573_, _05110_);
  nand (_00574_, _00523_, _11559_);
  and (_00575_, _00574_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00576_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00577_, _00576_, _08245_);
  and (_00578_, _00577_, _00523_);
  or (_00579_, _00578_, _00575_);
  and (_00580_, _00579_, _05794_);
  and (_00581_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00582_, _00550_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor (_00583_, _00550_, _07337_);
  or (_00584_, _00583_, _00582_);
  and (_00585_, _00584_, _05806_);
  or (_00586_, _00585_, _00581_);
  or (_00587_, _00586_, _00580_);
  and (_13360_, _00587_, _05110_);
  or (_00588_, _12745_, _12723_);
  nor (_00589_, _12747_, _07437_);
  and (_00591_, _00589_, _00588_);
  nor (_00592_, _07436_, _05195_);
  or (_00593_, _00592_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00594_, _00593_, _00591_);
  or (_00595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _11510_);
  and (_00596_, _00595_, _05110_);
  and (_00004_, _00596_, _00594_);
  and (_00597_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_00598_, _06088_, _06000_);
  and (_00599_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_00600_, _00599_, _00598_);
  and (_00601_, _00600_, _05337_);
  or (_00602_, _00601_, _00597_);
  and (_00018_, _00602_, _05110_);
  nand (_00603_, _12750_, _12715_);
  and (_00604_, _00603_, _12751_);
  or (_00605_, _00604_, _07437_);
  or (_00606_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00607_, _00606_, _12757_);
  and (_00608_, _00607_, _00605_);
  and (_00609_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_00028_, _00609_, _00608_);
  nand (_00610_, _08257_, _06798_);
  or (_00611_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_00612_, _00611_, _05110_);
  and (_00031_, _00612_, _00610_);
  or (_00613_, _12749_, _12717_);
  and (_00614_, _00613_, _12750_);
  or (_00615_, _00614_, _07437_);
  or (_00616_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00617_, _00616_, _12757_);
  and (_00618_, _00617_, _00615_);
  and (_00619_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00035_, _00619_, _00618_);
  and (_00620_, _12748_, _12719_);
  nor (_00621_, _00620_, _12749_);
  or (_00622_, _00621_, _07437_);
  or (_00623_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00624_, _00623_, _12757_);
  and (_00625_, _00624_, _00622_);
  and (_00626_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_00038_, _00626_, _00625_);
  or (_00627_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_00628_, _00627_, _05110_);
  nand (_00629_, _08257_, _06088_);
  and (_00128_, _00629_, _00628_);
  nor (_00630_, _11681_, _11481_);
  nor (_00631_, _00630_, _11682_);
  or (_00632_, _00631_, _07437_);
  or (_00633_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00634_, _00633_, _12757_);
  and (_00635_, _00634_, _00632_);
  and (_00636_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00253_, _00636_, _00635_);
  nand (_00637_, _08257_, _06229_);
  or (_00638_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_00639_, _00638_, _05110_);
  and (_00263_, _00639_, _00637_);
  nor (_00640_, _11689_, _11673_);
  nor (_00641_, _00640_, _11690_);
  or (_00642_, _00641_, _07437_);
  or (_00643_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00644_, _00643_, _12757_);
  and (_00645_, _00644_, _00642_);
  and (_00646_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_00273_, _00646_, _00645_);
  or (_00647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _11510_);
  and (_00649_, _00647_, _05110_);
  or (_00650_, _11688_, _11686_);
  nor (_00651_, _11689_, _07437_);
  and (_00652_, _00651_, _00650_);
  nor (_00653_, _07436_, _05220_);
  or (_00654_, _00653_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00655_, _00654_, _00652_);
  and (_00302_, _00655_, _00649_);
  nor (_00656_, _11684_, _11682_);
  nor (_00657_, _00656_, _11685_);
  or (_00658_, _00657_, _07437_);
  or (_00659_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00660_, _00659_, _12757_);
  and (_00661_, _00660_, _00658_);
  and (_00662_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00306_, _00662_, _00661_);
  and (_00663_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_00664_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_00665_, pc_log_change, _00664_);
  or (_00666_, _00665_, _00663_);
  and (_00377_, _00666_, _05110_);
  and (_00667_, _00047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_00668_, _00245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_00669_, _00668_, _00667_);
  and (_00670_, _00669_, _00244_);
  and (_00671_, _00238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_00672_, _00671_, _00667_);
  and (_00673_, _00672_, _00165_);
  or (_00674_, _00667_, _00074_);
  and (_00675_, _00674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_00676_, _00675_, _00673_);
  or (_00677_, _00676_, _00670_);
  nor (_00678_, _00036_, rst);
  and (_00679_, _00678_, _00069_);
  and (_00383_, _00679_, _00677_);
  nand (_00680_, _00048_, _05901_);
  and (_00681_, _00245_, _00243_);
  or (_00682_, _00681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_00683_, _00681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_00684_, _00683_, _00682_);
  and (_00685_, _00684_, _00261_);
  nand (_00686_, _00230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_00687_, _00230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_00688_, _00687_, _00686_);
  and (_00689_, _00688_, _00267_);
  or (_00690_, _00238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_00691_, _00671_, _00237_);
  and (_00692_, _00691_, _00690_);
  or (_00693_, _00692_, _00689_);
  or (_00694_, _00693_, _00685_);
  or (_00695_, _00694_, _00048_);
  and (_00696_, _00695_, _00680_);
  or (_00697_, _00696_, _00036_);
  or (_00698_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_00699_, _00698_, _05110_);
  and (_00385_, _00699_, _00697_);
  and (_00700_, _00166_, _00179_);
  or (_00701_, _00700_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_00702_, _00243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_00703_, _00702_, _00059_);
  nand (_00704_, _00703_, _00074_);
  or (_00705_, _00704_, _00048_);
  and (_00706_, _00705_, _00678_);
  and (_00707_, _00706_, _00701_);
  nand (_00708_, _00036_, _05110_);
  nor (_00709_, _00708_, _05901_);
  or (_00387_, _00709_, _00707_);
  nand (_00710_, _00452_, _05901_);
  or (_00711_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_00712_, _00711_, _05110_);
  and (_00395_, _00712_, _00710_);
  not (_00713_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_00714_, _00220_, _00713_);
  and (_00715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00716_, _00715_, _00226_);
  or (_00717_, _00716_, _00714_);
  and (_00718_, _00717_, _00267_);
  and (_00399_, _00718_, _00679_);
  and (_00411_, t0_i, _05110_);
  nand (_00719_, _13171_, _05901_);
  nor (_00720_, _13202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_00721_, _00720_, _13251_);
  and (_00722_, _00721_, _13180_);
  and (_00723_, _13181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand (_00724_, _13252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_00725_, _00724_, _13179_);
  or (_00726_, _00725_, _00723_);
  or (_00727_, _00726_, _00722_);
  or (_00728_, _00727_, _13171_);
  and (_00729_, _00728_, _05110_);
  and (_00415_, _00729_, _00719_);
  not (_00730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_00731_, _13193_, _00730_);
  and (_00732_, _13193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_00733_, _00732_, _13420_);
  and (_00734_, _00733_, _13414_);
  and (_00735_, _00734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_00736_, _00735_, _00731_);
  and (_00737_, _00736_, _13177_);
  and (_00738_, _13420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00739_, _00738_, _13391_);
  and (_00740_, _00739_, _00732_);
  or (_00741_, _00740_, _00731_);
  and (_00742_, _00741_, _13356_);
  nand (_00743_, _13193_, _13174_);
  and (_00744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00745_, _00744_, _00743_);
  or (_00746_, _00745_, _13252_);
  or (_00747_, _00746_, _00742_);
  or (_00748_, _00747_, _00737_);
  nor (_00749_, _13171_, _13179_);
  and (_00750_, _00749_, _05110_);
  and (_00417_, _00750_, _00748_);
  nand (_00751_, _13179_, _05901_);
  not (_00752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_00753_, _00150_, _00752_);
  and (_00754_, _00150_, _00752_);
  or (_00755_, _00754_, _00753_);
  or (_00756_, _00755_, _13179_);
  and (_00757_, _00756_, _13371_);
  and (_00758_, _00757_, _00751_);
  and (_00759_, _13250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_00760_, _00759_, _00758_);
  and (_00419_, _00760_, _05110_);
  and (_00422_, t1_i, _05110_);
  or (_00761_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_00762_, _00761_, _05110_);
  nand (_00763_, _08257_, _05841_);
  and (_00451_, _00763_, _00762_);
  and (_00764_, _12344_, _06745_);
  nor (_00765_, _12392_, _06780_);
  not (_00766_, _12067_);
  and (_00768_, _12347_, _00766_);
  or (_00770_, _12765_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00771_, _00770_, _12766_);
  and (_00772_, _00771_, _12374_);
  and (_00773_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_00774_, _00773_, _00772_);
  or (_00775_, _00774_, _00768_);
  or (_00776_, _00775_, _00765_);
  nor (_00777_, _00776_, _00764_);
  nand (_00778_, _00777_, _12343_);
  nand (_00779_, _12786_, _12404_);
  or (_00780_, _12780_, _12404_);
  and (_00781_, _00780_, _00779_);
  nor (_00782_, _00781_, _05613_);
  and (_00783_, _00781_, _05613_);
  or (_00784_, _00783_, _00782_);
  and (_00786_, _00784_, _13330_);
  or (_00787_, _00786_, _00778_);
  nor (_00788_, _12804_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_00789_, _00788_, _12805_);
  or (_00790_, _00789_, _12343_);
  and (_00791_, _00790_, _05110_);
  and (_00462_, _00791_, _00787_);
  nor (_00793_, _12785_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00794_, _00793_, _00779_);
  nand (_00795_, _12778_, _05123_);
  and (_00797_, _00795_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_00798_, _00797_, _12780_);
  and (_00799_, _00798_, _12403_);
  or (_00800_, _00799_, _00794_);
  and (_00801_, _00800_, _13330_);
  and (_00802_, _12344_, _07277_);
  and (_00803_, _12347_, _12417_);
  nor (_00804_, _12392_, _06548_);
  nor (_00805_, _12764_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00806_, _00805_, _12765_);
  and (_00807_, _00806_, _12374_);
  and (_00808_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00809_, _00808_, _00807_);
  or (_00810_, _00809_, _00804_);
  or (_00811_, _00810_, _00803_);
  nor (_00812_, _00811_, _00802_);
  nand (_00813_, _00812_, _12343_);
  or (_00814_, _00813_, _00801_);
  nor (_00815_, _12803_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_00816_, _00815_, _12804_);
  or (_00817_, _00816_, _12343_);
  and (_00818_, _00817_, _05110_);
  and (_00467_, _00818_, _00814_);
  or (_00819_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_00820_, _00819_, _05110_);
  nand (_00821_, _08257_, _06054_);
  and (_00472_, _00821_, _00820_);
  and (_00822_, _12344_, _07204_);
  not (_00823_, _07490_);
  and (_00825_, _12347_, _00823_);
  and (_00826_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00827_, _12386_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00828_, _00827_, _12764_);
  and (_00829_, _00828_, _12374_);
  nor (_00830_, _12392_, _07235_);
  or (_00831_, _00830_, _00829_);
  or (_00832_, _00831_, _00826_);
  or (_00833_, _00832_, _00825_);
  nor (_00834_, _00833_, _00822_);
  nand (_00835_, _00834_, _12343_);
  and (_00836_, _12784_, _12404_);
  and (_00837_, _12778_, _12403_);
  nor (_00838_, _00837_, _00836_);
  nand (_00839_, _00838_, _05123_);
  or (_00840_, _00838_, _05123_);
  and (_00841_, _00840_, _00839_);
  and (_00842_, _00841_, _12540_);
  or (_00843_, _00842_, _00835_);
  nor (_00844_, _12802_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00845_, _00844_, _12803_);
  or (_00846_, _00845_, _12343_);
  and (_00847_, _00846_, _05110_);
  and (_00483_, _00847_, _00843_);
  nor (_00590_, _11787_, rst);
  and (_00848_, _08614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_00849_, _08617_, _06230_);
  nand (_00850_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_00851_, _00850_, _06004_);
  or (_00852_, _00851_, _00849_);
  or (_00853_, _00852_, _00848_);
  and (_00648_, _00853_, _05110_);
  or (_00854_, _12524_, _12522_);
  and (_00855_, _13330_, _13332_);
  and (_00856_, _00855_, _00854_);
  not (_00857_, _12458_);
  and (_00858_, _00857_, _12347_);
  not (_00859_, _07235_);
  and (_00860_, _13340_, _00859_);
  and (_00861_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_00862_, _12374_, _00823_);
  or (_00863_, _00862_, _00861_);
  or (_00864_, _00863_, _00860_);
  or (_00865_, _00864_, _00858_);
  or (_00866_, _00865_, _00856_);
  and (_00867_, _00866_, _12343_);
  nor (_00868_, _07607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00869_, _00868_, _12546_);
  nor (_00870_, _00869_, _12343_);
  or (_00872_, _00870_, _00867_);
  and (_00767_, _00872_, _05110_);
  not (_00873_, _12343_);
  or (_00874_, _12471_, _12472_);
  not (_00875_, _00874_);
  nand (_00876_, _00875_, _12520_);
  or (_00877_, _00875_, _12520_);
  and (_00878_, _00877_, _13330_);
  and (_00879_, _00878_, _00876_);
  not (_00880_, _06668_);
  and (_00881_, _13340_, _00880_);
  not (_00882_, _07561_);
  and (_00883_, _12347_, _00882_);
  and (_00885_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_00886_, _12374_, _12346_);
  or (_00887_, _00886_, _00885_);
  or (_00888_, _00887_, _00883_);
  or (_00889_, _00888_, _00881_);
  or (_00890_, _00889_, _00879_);
  or (_00891_, _00890_, _00873_);
  or (_00892_, _12343_, _07609_);
  and (_00893_, _00892_, _05110_);
  and (_00769_, _00893_, _00891_);
  nand (_00894_, _12374_, _12473_);
  or (_00895_, _12518_, _12516_);
  nand (_00896_, _00895_, _12540_);
  or (_00897_, _00896_, _12519_);
  and (_00898_, _12347_, _12475_);
  not (_00899_, _07337_);
  and (_00900_, _13340_, _00899_);
  and (_00901_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_00902_, _00901_, _00900_);
  nor (_00903_, _00902_, _00898_);
  and (_00904_, _00903_, _00897_);
  nand (_00905_, _00904_, _00894_);
  and (_00906_, _00905_, _12343_);
  and (_00907_, _00873_, _07620_);
  or (_00908_, _00907_, _00906_);
  and (_00785_, _00908_, _05110_);
  and (_00909_, _12347_, _12482_);
  and (_00910_, _12374_, _12480_);
  or (_00911_, _00910_, _00909_);
  not (_00912_, _06512_);
  and (_00913_, _13340_, _00912_);
  and (_00914_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00916_, _00914_, _00913_);
  nor (_00917_, _12513_, _12510_);
  nor (_00918_, _00917_, _12514_);
  and (_00919_, _00918_, _12540_);
  or (_00920_, _00919_, _00916_);
  or (_00922_, _00920_, _00911_);
  or (_00923_, _00922_, _00873_);
  or (_00924_, _12343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00925_, _00924_, _05110_);
  and (_00792_, _00925_, _00923_);
  not (_00926_, _07418_);
  and (_00927_, _13340_, _00926_);
  and (_00928_, _12507_, _12347_);
  and (_00930_, _12374_, _12486_);
  and (_00932_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00934_, _00932_, _00930_);
  or (_00935_, _00934_, _00928_);
  or (_00936_, _00935_, _00927_);
  nor (_00937_, _12509_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00938_, _00937_, _12510_);
  and (_00939_, _00938_, _12540_);
  or (_00940_, _00939_, _00936_);
  or (_00941_, _00940_, _00873_);
  or (_00942_, _12343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00943_, _00942_, _05110_);
  and (_00796_, _00943_, _00941_);
  and (_00824_, _06411_, _05110_);
  and (_00944_, _12344_, _07364_);
  and (_00945_, _12374_, _11340_);
  and (_00946_, _12347_, _12480_);
  and (_00947_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00948_, _12392_, _06512_);
  or (_00949_, _00948_, _00947_);
  or (_00950_, _00949_, _00946_);
  or (_00951_, _00950_, _00945_);
  or (_00952_, _00951_, _00944_);
  and (_00953_, _12528_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00954_, _00953_, _12403_);
  and (_00955_, _12529_, _12403_);
  nor (_00956_, _00955_, _00954_);
  or (_00957_, _00956_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_00958_, _00956_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00959_, _00958_, _00957_);
  and (_00960_, _00959_, _12540_);
  nor (_00961_, _00960_, _00952_);
  nand (_00962_, _00961_, _12343_);
  nor (_00963_, _12550_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00964_, _00963_, _12551_);
  or (_00965_, _00964_, _12343_);
  and (_00966_, _00965_, _05110_);
  and (_00871_, _00966_, _00962_);
  and (_00967_, _12344_, _07391_);
  and (_00968_, _12374_, _06909_);
  and (_00969_, _12347_, _12486_);
  and (_00970_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00971_, _11309_, _00926_);
  or (_00972_, _00971_, _00970_);
  or (_00973_, _00972_, _00969_);
  or (_00974_, _00973_, _00968_);
  or (_00975_, _00974_, _00967_);
  nand (_00976_, _12528_, _05240_);
  or (_00977_, _12528_, _05240_);
  and (_00978_, _00977_, _00976_);
  and (_00979_, _00978_, _12403_);
  and (_00980_, _00954_, _12529_);
  or (_00981_, _00980_, _00979_);
  and (_00982_, _00981_, _13330_);
  or (_00983_, _00982_, _00975_);
  and (_00984_, _00983_, _12343_);
  nor (_00985_, _12549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00986_, _00985_, _12550_);
  nor (_00987_, _00986_, _12343_);
  or (_00988_, _00987_, _00984_);
  and (_00884_, _00988_, _05110_);
  and (_00989_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_00990_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_00991_, pc_log_change, _00990_);
  or (_00992_, _00991_, _00989_);
  and (_00915_, _00992_, _05110_);
  and (_00993_, _06904_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_00994_, _06901_, _12874_);
  or (_00995_, _00994_, _00993_);
  and (_00921_, _00995_, _05110_);
  or (_00996_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_00997_, _00996_, _08243_);
  and (_00998_, _05782_, _08272_);
  not (_00999_, _08272_);
  nand (_01000_, _00999_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_01002_, _01000_, _08243_);
  or (_01003_, _01002_, _00998_);
  and (_01004_, _01003_, _00997_);
  or (_01005_, _01004_, _08253_);
  nand (_01006_, _08253_, _05938_);
  and (_01007_, _01006_, _05110_);
  and (_00929_, _01007_, _01005_);
  and (_01008_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01009_, _07028_);
  and (_01010_, _13340_, _01009_);
  not (_01011_, _07176_);
  and (_01012_, _12347_, _01011_);
  and (_01013_, _12374_, _12762_);
  or (_01014_, _01013_, _01012_);
  or (_01015_, _01014_, _01010_);
  and (_01016_, _12525_, _12522_);
  or (_01017_, _01016_, _12465_);
  and (_01018_, _01017_, _12415_);
  nor (_01019_, _01018_, _12409_);
  nor (_01020_, _01019_, _12411_);
  and (_01021_, _01019_, _12411_);
  or (_01022_, _01021_, _01020_);
  and (_01023_, _01022_, _12540_);
  or (_01024_, _01023_, _01015_);
  nor (_01025_, _01024_, _01008_);
  nand (_01026_, _01025_, _12343_);
  nor (_01027_, _12548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_01028_, _01027_, _12549_);
  or (_01029_, _01028_, _12343_);
  and (_01030_, _01029_, _05110_);
  and (_00931_, _01030_, _01026_);
  not (_01031_, _07582_);
  and (_01032_, _12347_, _01031_);
  and (_01033_, _12374_, _00766_);
  or (_01034_, _01033_, _01032_);
  not (_01035_, _06780_);
  and (_01036_, _13340_, _01035_);
  and (_01037_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_01038_, _01037_, _01036_);
  nor (_01039_, _01017_, _12415_);
  nor (_01040_, _01039_, _01018_);
  and (_01041_, _01040_, _12540_);
  or (_01042_, _01041_, _01038_);
  or (_01044_, _01042_, _01034_);
  and (_01045_, _01044_, _12343_);
  nor (_01046_, _12547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_01047_, _01046_, _12548_);
  nor (_01048_, _01047_, _12343_);
  or (_01049_, _01048_, _01045_);
  and (_00933_, _01049_, _05110_);
  not (_01050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand (_01051_, _01050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_01052_, _01051_, _08235_);
  and (_01053_, _01052_, _08237_);
  or (_01054_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_01055_, _01054_, _08243_);
  and (_01056_, _05782_, _05805_);
  not (_01057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_01058_, _05805_, _01057_);
  nand (_01059_, _01058_, _08243_);
  or (_01060_, _01059_, _01056_);
  and (_01061_, _01060_, _01055_);
  or (_01062_, _01061_, _08253_);
  nand (_01063_, _08253_, _06798_);
  and (_01064_, _01063_, _05110_);
  and (_01043_, _01064_, _01062_);
  and (_01065_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_01066_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01447_, _01066_, _01065_);
  not (_01067_, _08243_);
  or (_01068_, _10212_, _01067_);
  and (_01069_, _01068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_01070_, _01069_, _08253_);
  and (_01071_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_01072_, _01071_, _10209_);
  and (_01073_, _01072_, _08243_);
  or (_01074_, _01073_, _01070_);
  nand (_01075_, _08253_, _05334_);
  and (_01076_, _01075_, _05110_);
  and (_01453_, _01076_, _01074_);
  and (_01077_, _05795_, _05419_);
  and (_01078_, _01077_, _05460_);
  and (_01079_, _01078_, _06122_);
  not (_01080_, _01079_);
  or (_01081_, _10212_, _01080_);
  and (_01082_, _01081_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01083_, _01082_, _06148_);
  and (_01084_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01085_, _01084_, _10209_);
  and (_01086_, _01085_, _06153_);
  or (_01087_, _01086_, _01083_);
  nand (_01088_, _06148_, _05334_);
  and (_01089_, _01088_, _05110_);
  and (_01459_, _01089_, _01087_);
  and (_01090_, _06153_, _08272_);
  or (_01091_, _01090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_01092_, _01091_, _06149_);
  nand (_01093_, _01090_, _05872_);
  and (_01094_, _01093_, _01092_);
  nor (_01095_, _06149_, _05938_);
  or (_01096_, _01095_, _01094_);
  and (_01460_, _01096_, _05110_);
  and (_01097_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01098_, _01097_, _10209_);
  and (_01099_, _01098_, _06123_);
  not (_01100_, _06123_);
  or (_01101_, _10212_, _01100_);
  and (_01102_, _01101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01103_, _01102_, _06129_);
  or (_01104_, _01103_, _01099_);
  nand (_01105_, _06129_, _05334_);
  and (_01106_, _01105_, _05110_);
  and (_01463_, _01106_, _01104_);
  and (_01107_, _06123_, _08272_);
  nand (_01108_, _01107_, _05872_);
  or (_01109_, _01107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_01110_, _01109_, _06130_);
  and (_01111_, _01110_, _01108_);
  nor (_01112_, _06130_, _05938_);
  or (_01113_, _01112_, _01111_);
  and (_01465_, _01113_, _05110_);
  nand (_01114_, _08243_, _05401_);
  and (_01115_, _01114_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_01116_, _01115_, _08253_);
  and (_01117_, _11559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_01118_, _01117_, _06632_);
  and (_01119_, _01118_, _08243_);
  or (_01120_, _01119_, _01116_);
  nand (_01121_, _08253_, _06088_);
  and (_01122_, _01121_, _05110_);
  and (_01468_, _01122_, _01120_);
  nor (_01123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01124_, _01123_, _05976_);
  nor (_01125_, _01124_, _06105_);
  nand (_01126_, _05980_, _05860_);
  not (_01127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nand (_01128_, _05973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_01129_, _01128_, _01127_);
  nor (_01130_, _05972_, _05850_);
  or (_01131_, _01130_, _05980_);
  or (_01132_, _01131_, _01129_);
  and (_01133_, _01132_, _06104_);
  and (_01134_, _01133_, _01126_);
  or (_01135_, _01134_, _01125_);
  nand (_01136_, _05976_, _05860_);
  and (_01137_, _01136_, _01135_);
  nand (_01138_, _01137_, _06099_);
  not (_01139_, _05971_);
  nor (_01140_, _06099_, _01139_);
  nand (_01141_, _01140_, _01127_);
  nor (_01142_, _01123_, _05967_);
  and (_01143_, _05946_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01144_, _01143_, _05955_);
  and (_01145_, _05951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01146_, _01145_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01147_, _01146_, _05967_);
  and (_01148_, _01147_, _01144_);
  or (_01149_, _01148_, _01142_);
  and (_01150_, _01149_, _05960_);
  and (_01151_, _05967_, _05955_);
  or (_01152_, _01151_, _05959_);
  nand (_01153_, _01152_, _05860_);
  nand (_01154_, _01153_, _06100_);
  or (_01155_, _01154_, _01150_);
  and (_01156_, _01155_, _01141_);
  and (_01157_, _01156_, _01138_);
  or (_01158_, _01157_, _05986_);
  nand (_01159_, _05986_, _01127_);
  and (_01160_, _01159_, _05110_);
  and (_01471_, _01160_, _01158_);
  nand (_01161_, _01140_, _06092_);
  nor (_01162_, _05986_, _06099_);
  or (_01163_, _01162_, _05850_);
  and (_01164_, _01163_, _05110_);
  and (_01475_, _01164_, _01161_);
  nand (_01165_, _05969_, _06110_);
  nor (_01166_, _01165_, _06099_);
  and (_01167_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  not (_01168_, _05982_);
  or (_01169_, _06098_, _01168_);
  nor (_01170_, _01169_, _05975_);
  and (_01171_, _01170_, _06137_);
  or (_01172_, _01171_, _01167_);
  or (_01173_, _01172_, _01166_);
  and (_01478_, _01173_, _05110_);
  and (_01479_, _13167_, _05986_);
  and (_01174_, _06625_, _05789_);
  and (_01175_, _01174_, _05867_);
  nand (_01176_, _01175_, _05872_);
  or (_01177_, _01175_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_01178_, _01177_, _05794_);
  and (_01179_, _01178_, _01176_);
  and (_01180_, _05804_, _05992_);
  nand (_01181_, _01180_, _05901_);
  or (_01182_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_01183_, _01182_, _05806_);
  and (_01184_, _01183_, _01181_);
  and (_01185_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_01186_, _01185_, rst);
  or (_01187_, _01186_, _01184_);
  or (_01488_, _01187_, _01179_);
  and (_01188_, _06153_, _08133_);
  or (_01189_, _01188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01190_, _01189_, _06149_);
  nand (_01191_, _01188_, _05872_);
  and (_01192_, _01191_, _01190_);
  nor (_01193_, _06149_, _06054_);
  or (_01194_, _01193_, _01192_);
  and (_01494_, _01194_, _05110_);
  and (_01195_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_01196_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_01498_, _01196_, _01195_);
  and (_01197_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_01198_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_01500_, _01198_, _01197_);
  and (_01199_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_01200_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_01513_, _01200_, _01199_);
  and (_01201_, _06123_, _08133_);
  nand (_01202_, _01201_, _05872_);
  or (_01203_, _01201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_01204_, _01203_, _06130_);
  and (_01205_, _01204_, _01202_);
  nor (_01206_, _06130_, _06054_);
  or (_01207_, _01206_, _01205_);
  and (_01516_, _01207_, _05110_);
  and (_01520_, _00496_, _05986_);
  and (_01208_, _05798_, _05805_);
  or (_01209_, _01208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01210_, _01209_, _05844_);
  nand (_01211_, _01208_, _05872_);
  and (_01212_, _01211_, _01210_);
  and (_01213_, _06799_, _05809_);
  or (_01214_, _01213_, _01212_);
  and (_01522_, _01214_, _05110_);
  nor (_01215_, _01140_, _05986_);
  not (_01216_, _01215_);
  and (_01217_, _01216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_01218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_01219_, _05973_, _05850_);
  or (_01220_, _01219_, _01218_);
  nor (_01221_, _05972_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01222_, _01221_, _05980_);
  nand (_01223_, _01222_, _01220_);
  or (_01224_, _06114_, _05849_);
  and (_01225_, _01224_, _01223_);
  or (_01226_, _01225_, _05979_);
  not (_01227_, _05977_);
  not (_01228_, _05979_);
  or (_01229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _05850_);
  or (_01230_, _01229_, _01228_);
  and (_01231_, _01230_, _01227_);
  and (_01232_, _01231_, _01226_);
  and (_01233_, _05977_, _05849_);
  or (_01234_, _01233_, _05976_);
  or (_01235_, _01234_, _01232_);
  or (_01236_, _01229_, _06103_);
  and (_01237_, _01236_, _06099_);
  and (_01238_, _01237_, _01235_);
  and (_01239_, _05951_, _05850_);
  or (_01240_, _01239_, _01218_);
  and (_01241_, _05946_, _05850_);
  nor (_01242_, _01241_, _05955_);
  nand (_01243_, _01242_, _01240_);
  or (_01244_, _05956_, _05849_);
  and (_01245_, _01244_, _01243_);
  or (_01246_, _01245_, _05966_);
  not (_01247_, _05963_);
  not (_01248_, _05966_);
  or (_01249_, _01229_, _01248_);
  and (_01250_, _01249_, _01247_);
  and (_01251_, _01250_, _01246_);
  and (_01252_, _05963_, _05849_);
  or (_01253_, _01252_, _05959_);
  or (_01254_, _01253_, _01251_);
  and (_01255_, _06100_, _05960_);
  and (_01256_, _01229_, _06100_);
  or (_01257_, _01256_, _01255_);
  and (_01258_, _01257_, _01254_);
  or (_01259_, _01258_, _01238_);
  and (_01260_, _01259_, _06137_);
  or (_01261_, _01260_, _01217_);
  and (_01527_, _01261_, _05110_);
  and (_01531_, _06388_, _05110_);
  nor (_01262_, _05841_, _05465_);
  and (_01263_, _05465_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_01264_, _01263_, _01262_);
  and (_01540_, _01264_, _05110_);
  and (_01561_, _06366_, _05110_);
  and (_01265_, _05798_, _10208_);
  or (_01266_, _01265_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01267_, _01266_, _05844_);
  nand (_01268_, _01265_, _05872_);
  and (_01269_, _01268_, _01267_);
  nor (_01270_, _05844_, _05334_);
  or (_01271_, _01270_, _01269_);
  and (_01565_, _01271_, _05110_);
  and (_01272_, _05798_, _06472_);
  nand (_01273_, _01272_, _05872_);
  or (_01274_, _01272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_01275_, _01274_, _05844_);
  and (_01276_, _01275_, _01273_);
  nor (_01277_, _06229_, _05844_);
  or (_01278_, _01277_, _01276_);
  and (_01567_, _01278_, _05110_);
  and (_01279_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_01280_, _01279_, _01215_);
  and (_01571_, _01280_, _05110_);
  and (_01281_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_01282_, _01281_, _01215_);
  and (_01574_, _01282_, _05110_);
  and (_01283_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_01284_, _08617_, _12894_);
  or (_01285_, _01284_, _01283_);
  and (_01577_, _01285_, _05110_);
  or (_01286_, _05966_, _05955_);
  and (_01287_, _05952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01288_, _01287_, _01286_);
  and (_01289_, _01288_, _01247_);
  and (_01290_, _01289_, _01255_);
  nand (_01291_, _05975_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nand (_01292_, _01291_, _05981_);
  and (_01293_, _01292_, _05978_);
  and (_01294_, _01293_, _06099_);
  or (_01295_, _01294_, _05986_);
  or (_01296_, _01295_, _01290_);
  nand (_01297_, _05986_, _11499_);
  and (_01298_, _01297_, _05110_);
  and (_01581_, _01298_, _01296_);
  nor (_01299_, _05951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01300_, _01299_, _05946_);
  or (_01301_, _01300_, _05955_);
  and (_01302_, _01301_, _01248_);
  or (_01303_, _01302_, _05963_);
  and (_01304_, _01303_, _01255_);
  and (_01305_, _06099_, _06103_);
  or (_01306_, _05973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01307_, _01306_, _05972_);
  or (_01308_, _01307_, _05980_);
  and (_01309_, _01308_, _01228_);
  or (_01310_, _01309_, _05977_);
  and (_01311_, _01310_, _01305_);
  or (_01312_, _01311_, _05986_);
  or (_01313_, _01312_, _01304_);
  or (_01314_, _06137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01315_, _01314_, _05110_);
  and (_01590_, _01315_, _01313_);
  nor (_01316_, _11268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_01317_, _01316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_01318_, _01316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_01319_, _01318_, _05110_);
  and (_01600_, _01319_, _01317_);
  not (_01320_, _06560_);
  nor (_01321_, _01320_, _05901_);
  and (_01322_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_01323_, _01322_, _01321_);
  and (_01604_, _01323_, _05110_);
  and (_01324_, _08750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not (_01325_, _08745_);
  and (_01326_, _08754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_01327_, _01326_, _01325_);
  or (_01328_, _01327_, _01324_);
  and (_01329_, _08754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_01330_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_01331_, _01330_, _05110_);
  and (_01619_, _01331_, _01328_);
  or (_01332_, _06984_, _07177_);
  nor (_01333_, _07208_, _07028_);
  and (_01334_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01335_, _01334_, _06471_);
  or (_01336_, _01335_, _01333_);
  and (_01337_, _01336_, _05110_);
  and (_01636_, _01337_, _01332_);
  and (_01338_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_01339_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_01340_, pc_log_change, _01339_);
  or (_01341_, _01340_, _01338_);
  and (_01646_, _01341_, _05110_);
  nand (_01342_, _07028_, _06477_);
  or (_01343_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01344_, _01343_, _05110_);
  and (_01669_, _01344_, _01342_);
  or (_01345_, _05718_, _05716_);
  not (_01346_, _05653_);
  nand (_01347_, _05716_, _01346_);
  and (_01348_, _01347_, _05650_);
  and (_01349_, _01348_, _01345_);
  nand (_01350_, _05646_, _05519_);
  and (_01351_, _05647_, _05489_);
  and (_01352_, _01351_, _01350_);
  and (_01353_, _06485_, ABINPUT000000[0]);
  and (_01354_, _06487_, ABINPUT000[0]);
  nor (_01355_, _01354_, _01353_);
  nand (_01356_, _01355_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_01357_, _01356_, _01352_);
  or (_01358_, _01357_, _01349_);
  or (_01359_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_01360_, _01359_, _01358_);
  and (_01361_, _01360_, _10211_);
  not (_01362_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_01363_, _06472_, _01362_);
  or (_01364_, _01363_, _08245_);
  and (_01365_, _01364_, _10157_);
  nor (_01366_, _01365_, _01361_);
  nand (_01367_, _01366_, _10163_);
  nand (_01368_, _10162_, _06229_);
  and (_01369_, _01368_, _05110_);
  and (_01741_, _01369_, _01367_);
  nor (_01370_, _06054_, _06010_);
  and (_01371_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_01372_, _01371_, _05995_);
  or (_01373_, _01372_, _01370_);
  or (_01374_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_01375_, _01374_, _05110_);
  and (_01746_, _01375_, _01373_);
  or (_01376_, _11202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_01377_, _06882_, _06897_);
  nand (_01378_, _01377_, _11223_);
  nand (_01379_, _01378_, _11203_);
  and (_01380_, _01379_, _01376_);
  or (_01381_, _01380_, _11193_);
  and (_01382_, _11193_, _06897_);
  nor (_01383_, _01382_, _11234_);
  and (_01384_, _01383_, _01381_);
  and (_01385_, _11234_, _06799_);
  or (_01386_, _01385_, _11239_);
  or (_01387_, _01386_, _01384_);
  nand (_01388_, _11239_, _06885_);
  and (_01389_, _01388_, _05110_);
  and (_01752_, _01389_, _01387_);
  or (_01390_, _06137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01391_, _01390_, _05110_);
  or (_01392_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _05850_);
  and (_01393_, _01392_, _06103_);
  or (_01394_, _01393_, _06105_);
  and (_01395_, _05980_, _05859_);
  or (_01396_, _01219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand (_01397_, _01396_, _01222_);
  nand (_01398_, _01397_, _06104_);
  or (_01399_, _01398_, _01395_);
  and (_01400_, _01399_, _01394_);
  and (_01401_, _05976_, _05859_);
  or (_01402_, _01401_, _01400_);
  and (_01403_, _01402_, _06099_);
  and (_01404_, _05971_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01405_, _01152_, _05859_);
  or (_01406_, _01239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01407_, _01242_, _05967_);
  and (_01408_, _01407_, _01406_);
  not (_01409_, _05967_);
  and (_01410_, _01392_, _01409_);
  or (_01411_, _01410_, _01408_);
  and (_01412_, _01411_, _05960_);
  or (_01413_, _01412_, _01405_);
  and (_01414_, _01413_, _01139_);
  nor (_01415_, _01414_, _01404_);
  nor (_01416_, _01415_, _06099_);
  or (_01417_, _01416_, _01403_);
  or (_01418_, _01417_, _05986_);
  and (_01756_, _01418_, _01391_);
  and (_01419_, _01216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_01420_, _01128_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_01421_, _01420_, _01131_);
  or (_01422_, _06114_, _05851_);
  and (_01423_, _01422_, _01421_);
  or (_01424_, _01423_, _05979_);
  or (_01425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_01426_, _01425_, _01228_);
  and (_01427_, _01426_, _01227_);
  and (_01428_, _01427_, _01424_);
  and (_01429_, _05977_, _05851_);
  or (_01430_, _01429_, _05976_);
  or (_01431_, _01430_, _01428_);
  or (_01432_, _01425_, _06103_);
  and (_01433_, _01432_, _06099_);
  and (_01434_, _01433_, _01431_);
  not (_01435_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_01436_, _01145_, _01435_);
  nand (_01437_, _01436_, _01144_);
  or (_01438_, _05956_, _05851_);
  and (_01439_, _01438_, _01437_);
  or (_01440_, _01439_, _05966_);
  or (_01441_, _01425_, _01248_);
  and (_01442_, _01441_, _01247_);
  and (_01443_, _01442_, _01440_);
  and (_01444_, _05963_, _05851_);
  or (_01445_, _01444_, _05959_);
  or (_01446_, _01445_, _01443_);
  and (_01448_, _01425_, _06100_);
  or (_01449_, _01448_, _01255_);
  and (_01450_, _01449_, _01446_);
  or (_01451_, _01450_, _01434_);
  and (_01452_, _01451_, _06137_);
  or (_01454_, _01452_, _01419_);
  and (_01759_, _01454_, _05110_);
  nand (_01455_, _06100_, _06092_);
  and (_01456_, _06092_, _06099_);
  or (_01457_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_01458_, _01457_, _05110_);
  and (_01763_, _01458_, _01455_);
  nor (_01461_, _05986_, _05850_);
  and (_01462_, _01461_, _06099_);
  or (_01464_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  nand (_01466_, _01461_, _06100_);
  and (_01467_, _01466_, _05110_);
  and (_01767_, _01467_, _01464_);
  and (_01469_, _06123_, _05805_);
  or (_01470_, _01469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01472_, _01470_, _06130_);
  nand (_01473_, _01469_, _05872_);
  and (_01474_, _01473_, _01472_);
  and (_01476_, _06799_, _06129_);
  or (_01477_, _01476_, _01474_);
  and (_01795_, _01477_, _05110_);
  and (_01480_, _06632_, _06123_);
  nand (_01481_, _06123_, _05401_);
  or (_01482_, _01481_, _11548_);
  and (_01483_, _01482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_01484_, _01483_, _06129_);
  or (_01485_, _01484_, _01480_);
  nand (_01486_, _06129_, _06088_);
  and (_01487_, _01486_, _05110_);
  and (_01799_, _01487_, _01485_);
  and (_01489_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01490_, _01489_, _08245_);
  and (_01491_, _01490_, _06123_);
  nand (_01492_, _06123_, _11559_);
  and (_01493_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_01495_, _01493_, _06129_);
  or (_01496_, _01495_, _01491_);
  nand (_01497_, _06229_, _06129_);
  and (_01499_, _01497_, _05110_);
  and (_01801_, _01499_, _01496_);
  and (_01501_, _06123_, _05488_);
  nand (_01502_, _01501_, _05872_);
  or (_01503_, _01501_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_01504_, _01503_, _06130_);
  and (_01505_, _01504_, _01502_);
  nor (_01506_, _06130_, _05841_);
  or (_01507_, _01506_, _01505_);
  and (_01804_, _01507_, _05110_);
  and (_01508_, _06153_, _05805_);
  or (_01509_, _01508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01510_, _01509_, _06149_);
  nand (_01511_, _01508_, _05872_);
  and (_01512_, _01511_, _01510_);
  and (_01514_, _06799_, _06148_);
  or (_01515_, _01514_, _01512_);
  and (_01812_, _01515_, _05110_);
  and (_01517_, _06632_, _01079_);
  nand (_01518_, _01079_, _05401_);
  or (_01519_, _01518_, _11548_);
  and (_01521_, _01519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_01523_, _01521_, _06148_);
  or (_01524_, _01523_, _01517_);
  nand (_01525_, _06148_, _06088_);
  and (_01526_, _01525_, _05110_);
  and (_01822_, _01526_, _01524_);
  or (_01528_, _01518_, _05866_);
  and (_01529_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01530_, _01529_, _06148_);
  and (_01532_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01533_, _01532_, _08245_);
  and (_01534_, _01533_, _06153_);
  or (_01535_, _01534_, _01530_);
  nand (_01536_, _06229_, _06148_);
  and (_01537_, _01536_, _05110_);
  and (_01826_, _01537_, _01535_);
  and (_01538_, _06153_, _05488_);
  or (_01539_, _01538_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_01541_, _01539_, _06149_);
  nand (_01542_, _01538_, _05872_);
  and (_01543_, _01542_, _01541_);
  nor (_01544_, _06149_, _05841_);
  or (_01545_, _01544_, _01543_);
  and (_01845_, _01545_, _05110_);
  or (_01546_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_01547_, _01546_, _11326_);
  and (_01548_, _05867_, _05782_);
  nand (_01549_, _12083_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_01550_, _01549_, _11326_);
  or (_01551_, _01550_, _01548_);
  and (_01552_, _01551_, _01547_);
  or (_01553_, _01552_, _11329_);
  nand (_01554_, _11329_, _05901_);
  and (_01555_, _01554_, _05110_);
  and (_01851_, _01555_, _01553_);
  nand (_01556_, _06890_, _05901_);
  and (_01557_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01558_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_01559_, _01558_, _01557_);
  or (_01560_, _01559_, _06890_);
  and (_01562_, _01560_, _08871_);
  and (_01563_, _01562_, _01556_);
  and (_01564_, _06895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_01566_, _01564_, _01563_);
  and (_01860_, _01566_, _05110_);
  and (_01568_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_01569_, pc_log_change, _05478_);
  or (_01570_, _01569_, _01568_);
  and (_01869_, _01570_, _05110_);
  nor (_01572_, _05841_, _06010_);
  and (_01573_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_01575_, _01573_, _05995_);
  or (_01576_, _01575_, _01572_);
  or (_01578_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_01579_, _01578_, _05110_);
  and (_01905_, _01579_, _01576_);
  nor (_01580_, _11584_, _11515_);
  and (_01582_, _11192_, _06881_);
  and (_01583_, _01582_, _11202_);
  and (_01584_, _01583_, _11223_);
  and (_01585_, _01584_, _11584_);
  or (_01586_, _01585_, _01580_);
  and (_01908_, _01586_, _05110_);
  nand (_01587_, _11239_, _05901_);
  or (_01588_, _12560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_01589_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_01591_, _01589_, _11202_);
  nand (_01592_, _01591_, _11223_);
  and (_01594_, _01592_, _01588_);
  or (_01595_, _01594_, _11193_);
  nor (_01596_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_01597_, _01596_, _11234_);
  and (_01598_, _01597_, _01595_);
  and (_01599_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_01601_, _01599_, _11239_);
  or (_01602_, _01601_, _01598_);
  and (_01603_, _01602_, _05110_);
  and (_01911_, _01603_, _01587_);
  nor (_01605_, _12612_, _05901_);
  and (_01606_, _11601_, _11215_);
  and (_01607_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01608_, _01607_, _11223_);
  or (_01609_, _01608_, _01606_);
  and (_01610_, _01609_, _11202_);
  and (_01611_, _11601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_01612_, _01611_, _11193_);
  or (_01613_, _01612_, _01610_);
  nor (_01614_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_01616_, _01614_, _11234_);
  and (_01617_, _01616_, _01613_);
  or (_01618_, _01617_, _11239_);
  or (_01620_, _01618_, _01605_);
  or (_01621_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_01622_, _01621_, _05110_);
  and (_01914_, _01622_, _01620_);
  and (_01623_, _11202_, _11190_);
  and (_01624_, _01623_, _11584_);
  or (_01625_, _01624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_01626_, _11223_);
  nand (_01627_, _01624_, _01626_);
  and (_01628_, _01627_, _05110_);
  and (_01917_, _01628_, _01625_);
  nand (_01629_, _08870_, _05901_);
  and (_01630_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_01631_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_01632_, _01631_, _01630_);
  or (_01633_, _01632_, _08870_);
  and (_01634_, _01633_, _05110_);
  and (_01920_, _01634_, _01629_);
  and (_01931_, t2ex_i, _05110_);
  nor (_01635_, t2ex_i, rst);
  and (_01934_, _01635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor (_01637_, t2_i, rst);
  and (_01937_, _01637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and (_01940_, t2_i, _05110_);
  or (_01638_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_01640_, pc_log_change, _01639_);
  and (_01641_, _01640_, _05110_);
  and (_02010_, _01641_, _01638_);
  or (_01642_, _06860_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_01643_, _06861_, _05110_);
  and (_01644_, _01643_, _01642_);
  and (_01645_, _06811_, _06434_);
  or (_01647_, _01645_, _06947_);
  or (_01648_, _01647_, _06816_);
  and (_01649_, _07079_, _07040_);
  or (_01650_, _01649_, _07046_);
  or (_01651_, _07081_, _06453_);
  or (_01652_, _01651_, _07089_);
  or (_01653_, _01652_, _01650_);
  or (_01654_, _01653_, _01648_);
  or (_01655_, _07093_, _07052_);
  or (_01656_, _01655_, _07074_);
  and (_01657_, _06457_, _07067_);
  and (_01658_, _06852_, _06455_);
  or (_01659_, _01658_, _01657_);
  or (_01660_, _01659_, _07078_);
  or (_01661_, _01660_, _06449_);
  or (_01662_, _07048_, _07041_);
  or (_01663_, _01662_, _01661_);
  and (_01664_, _13086_, _06434_);
  and (_01665_, _07138_, _06464_);
  or (_01666_, _01665_, _01664_);
  and (_01667_, _07079_, _06830_);
  or (_01668_, _01667_, _07039_);
  and (_01670_, _07087_, _06434_);
  or (_01671_, _01670_, _01668_);
  or (_01672_, _01671_, _01666_);
  or (_01673_, _13078_, _11749_);
  not (_01674_, _07095_);
  nand (_01675_, _11300_, _01674_);
  or (_01676_, _01675_, _01673_);
  or (_01677_, _01676_, _01672_);
  or (_01678_, _01677_, _01663_);
  or (_01679_, _01678_, _01656_);
  or (_01680_, _01679_, _01654_);
  and (_01681_, _01680_, _06842_);
  or (_02048_, _01681_, _01644_);
  nand (_01682_, _06294_, _05473_);
  or (_01683_, _05473_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_01684_, _01683_, _05110_);
  and (_02086_, _01684_, _01682_);
  and (_01685_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_01686_, _05938_, _06010_);
  or (_01687_, _01686_, _01685_);
  or (_01688_, _01687_, _05995_);
  or (_01689_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_01690_, _01689_, _05110_);
  and (_02207_, _01690_, _01688_);
  nand (_01691_, _06673_, _05938_);
  or (_01692_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_01693_, _01692_, _05110_);
  and (_02218_, _01693_, _01691_);
  nor (_01694_, _06088_, _06010_);
  and (_01695_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_01696_, _01695_, _05995_);
  or (_01697_, _01696_, _01694_);
  or (_01698_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_01699_, _01698_, _05110_);
  and (_02222_, _01699_, _01697_);
  or (_01700_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand (_01701_, _06205_, _12450_);
  and (_01702_, _01701_, _05110_);
  and (_02255_, _01702_, _01700_);
  and (_01703_, _06807_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_01704_, _07075_, _13076_);
  or (_01705_, _01704_, _01652_);
  or (_01706_, _11760_, _07096_);
  and (_01707_, _12149_, _06864_);
  and (_01708_, _01665_, _11802_);
  or (_01709_, _01708_, _01707_);
  or (_01710_, _01709_, _01706_);
  or (_01711_, _06838_, _06828_);
  and (_01712_, _07069_, _06434_);
  and (_01713_, _07038_, _06434_);
  or (_01714_, _01713_, _13078_);
  or (_01715_, _01714_, _01712_);
  or (_01716_, _01715_, _01711_);
  or (_01717_, _01716_, _01710_);
  or (_01718_, _01717_, _01705_);
  and (_01719_, _01718_, _06842_);
  or (_02391_, _01719_, _01703_);
  not (_01720_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_01721_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_01722_, _01721_, _01720_);
  and (_01723_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _05110_);
  and (_02407_, _01723_, _01722_);
  and (_01724_, _12330_, _12228_);
  nand (_01725_, _12018_, _11977_);
  and (_01726_, _12073_, _01725_);
  and (_01727_, _01726_, _11918_);
  and (_01728_, _01727_, _11960_);
  and (_01729_, _12268_, _11871_);
  and (_01730_, _01729_, _01728_);
  and (_01731_, _01730_, _01724_);
  and (_01732_, _01731_, _06471_);
  and (_01733_, _12071_, _01725_);
  and (_01734_, _01733_, _11918_);
  and (_01735_, _01734_, _11960_);
  and (_01736_, _12268_, _11873_);
  and (_01737_, _12330_, _12225_);
  and (_01738_, _01737_, _01736_);
  and (_01739_, _01738_, _01735_);
  and (_01740_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_01742_, _12270_, _11873_);
  and (_01743_, _01737_, _01742_);
  and (_01744_, _01743_, _01735_);
  and (_01745_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_01747_, _01745_, _01740_);
  and (_01748_, _12328_, _12225_);
  and (_01749_, _01748_, _01742_);
  and (_01750_, _01749_, _01735_);
  and (_01751_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_01753_, _01724_, _01736_);
  and (_01754_, _01753_, _01735_);
  and (_01755_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_01757_, _01755_, _01751_);
  or (_01758_, _01757_, _01747_);
  and (_01760_, _01738_, _01728_);
  and (_01761_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_01762_, _12328_, _12228_);
  and (_01764_, _01762_, _01736_);
  and (_01765_, _01764_, _01735_);
  and (_01766_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_01768_, _01766_, _01761_);
  and (_01769_, _01726_, _11920_);
  and (_01770_, _01769_, _11958_);
  or (_01771_, _12330_, _12225_);
  or (_01772_, _01771_, _12268_);
  nor (_01773_, _01772_, _11873_);
  and (_01774_, _01773_, _01770_);
  and (_01775_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_01776_, _01769_, _11960_);
  and (_01777_, _01776_, _01738_);
  and (_01778_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_01779_, _01778_, _01775_);
  or (_01780_, _01779_, _01768_);
  or (_01781_, _01780_, _01758_);
  and (_01782_, _01736_, _01748_);
  and (_01783_, _01728_, _01782_);
  and (_01784_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_01785_, _01764_, _01728_);
  and (_01786_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_01787_, _01786_, _01784_);
  and (_01788_, _01753_, _01728_);
  and (_01789_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01790_, _01728_, _01749_);
  and (_01791_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01792_, _01791_, _01789_);
  or (_01793_, _01792_, _01787_);
  and (_01794_, _01727_, _11958_);
  and (_01796_, _01794_, _01782_);
  and (_01797_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_01798_, _01738_, _01794_);
  and (_01800_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_01802_, _01800_, _01797_);
  and (_01803_, _01743_, _01728_);
  and (_01805_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01806_, _01773_, _01728_);
  and (_01807_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_01808_, _01807_, _01805_);
  or (_01809_, _01808_, _01802_);
  or (_01810_, _01809_, _01793_);
  or (_01811_, _01810_, _01781_);
  and (_01813_, _01737_, _01729_);
  and (_01814_, _01813_, _11958_);
  and (_01815_, _01733_, _11920_);
  and (_01816_, _01815_, _01814_);
  and (_01817_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01818_, _01729_, _01748_);
  and (_01819_, _01818_, _01728_);
  and (_01820_, _01819_, _11976_);
  or (_01821_, _01820_, _01817_);
  and (_01823_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01824_, _01762_, _01729_);
  and (_01825_, _01824_, _01728_);
  and (_01827_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_01828_, _01827_, _01823_);
  or (_01829_, _01828_, _01821_);
  and (_01830_, _01770_, _01813_);
  and (_01831_, _07079_, _06431_);
  nor (_01832_, _01831_, _06817_);
  and (_01833_, _01832_, _06834_);
  nor (_01834_, _01649_, _07074_);
  and (_01835_, _01834_, _01833_);
  nor (_01836_, _01665_, _11755_);
  nor (_01837_, _06938_, _06823_);
  and (_01838_, _07069_, _06810_);
  nor (_01839_, _01838_, _07095_);
  and (_01840_, _01839_, _01837_);
  and (_01841_, _01840_, _11747_);
  and (_01842_, _01841_, _01836_);
  and (_01843_, _01842_, _01835_);
  and (_01844_, _01843_, _11746_);
  nor (_01846_, _01844_, _12089_);
  or (_01847_, _01846_, p3_in[7]);
  not (_01848_, _01846_);
  or (_01849_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_01850_, _01849_, _01847_);
  and (_01852_, _01850_, _01830_);
  and (_01853_, _01776_, _01813_);
  or (_01854_, _01846_, p2_in[7]);
  or (_01855_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_01856_, _01855_, _01854_);
  and (_01857_, _01856_, _01853_);
  or (_01858_, _01857_, _01852_);
  and (_01859_, _01813_, _01728_);
  or (_01861_, _01846_, p0_in[7]);
  or (_01862_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_01863_, _01862_, _01861_);
  and (_01864_, _01863_, _01859_);
  and (_01865_, _01813_, _01794_);
  or (_01866_, _01846_, p1_in[7]);
  or (_01867_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_01868_, _01867_, _01866_);
  and (_01870_, _01868_, _01865_);
  or (_01871_, _01870_, _01864_);
  or (_01872_, _01871_, _01858_);
  or (_01873_, _01872_, _01829_);
  and (_01874_, _01814_, _01734_);
  and (_01875_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01876_, _01813_, _11960_);
  and (_01877_, _01815_, _01876_);
  and (_01878_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01879_, _01878_, _01875_);
  or (_01880_, _01879_, _01873_);
  or (_01881_, _01880_, _01811_);
  nand (_01882_, _01874_, _12172_);
  nand (_01883_, _01877_, _06613_);
  and (_01884_, _01883_, _01882_);
  nand (_01885_, _01825_, _06471_);
  nand (_01886_, _01885_, _01884_);
  nand (_01887_, _01886_, _05151_);
  nand (_01888_, _01877_, _06617_);
  and (_01889_, _01772_, _06150_);
  nand (_01890_, _01889_, _12082_);
  and (_01891_, _01890_, _01888_);
  and (_01892_, _01891_, _12340_);
  and (_01893_, _01892_, _01887_);
  and (_01894_, _01893_, _01881_);
  nor (_01895_, _01877_, _01874_);
  nand (_01896_, _01813_, _01726_);
  nor (_01897_, _01825_, _01731_);
  nor (_01898_, _01819_, _01816_);
  and (_01899_, _01898_, _01897_);
  and (_01900_, _01899_, _01896_);
  and (_01901_, _01900_, _01895_);
  nor (_01902_, _01744_, _01739_);
  nand (_01903_, _01733_, _11918_);
  or (_01904_, _01903_, _11958_);
  not (_01906_, _01742_);
  or (_01907_, _12330_, _12228_);
  or (_01909_, _01907_, _01906_);
  or (_01910_, _01909_, _01904_);
  nand (_01912_, _01724_, _01736_);
  or (_01913_, _01912_, _01904_);
  and (_01915_, _01913_, _01910_);
  and (_01916_, _01915_, _01902_);
  or (_01918_, _12071_, _12020_);
  or (_01919_, _01918_, _11920_);
  or (_01921_, _01919_, _11958_);
  not (_01922_, _01736_);
  or (_01923_, _12328_, _12228_);
  or (_01924_, _01923_, _01922_);
  or (_01925_, _01924_, _01921_);
  or (_01926_, _01771_, _01922_);
  or (_01927_, _01926_, _01904_);
  and (_01928_, _01927_, _01925_);
  nor (_01929_, _01777_, _01774_);
  and (_01930_, _01929_, _01928_);
  and (_01932_, _01930_, _01916_);
  or (_01933_, _01922_, _01907_);
  or (_01935_, _01921_, _01933_);
  or (_01936_, _01926_, _01921_);
  and (_01938_, _01936_, _01935_);
  nor (_01939_, _01790_, _01788_);
  and (_01941_, _01939_, _01938_);
  nor (_01942_, _01806_, _01803_);
  nor (_01943_, _01798_, _01796_);
  and (_01944_, _01943_, _01942_);
  and (_01945_, _01944_, _01941_);
  and (_01946_, _01945_, _01932_);
  nand (_01947_, _01946_, _01901_);
  nand (_01948_, _01947_, _01893_);
  and (_01949_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_01950_, _01949_, _01894_);
  or (_01951_, _01950_, _01732_);
  nand (_01952_, _01732_, _07028_);
  and (_01953_, _01952_, _05110_);
  and (_02423_, _01953_, _01951_);
  and (_01954_, _00523_, _10209_);
  nand (_01955_, _00523_, _10208_);
  and (_01956_, _01955_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_01957_, _01956_, _01954_);
  and (_01958_, _01957_, _05794_);
  and (_01959_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_01960_, _00531_, _07235_);
  or (_01961_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01962_, _01961_, _05806_);
  and (_01963_, _01962_, _01960_);
  or (_01964_, _01963_, _01959_);
  or (_01965_, _01964_, _01958_);
  and (_02463_, _01965_, _05110_);
  and (_01966_, _00523_, _08272_);
  nand (_01967_, _01966_, _05872_);
  or (_01968_, _01966_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01969_, _01968_, _05794_);
  and (_01970_, _01969_, _01967_);
  and (_01971_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01972_, _00550_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_01973_, _00550_, _06512_);
  or (_01974_, _01973_, _01972_);
  and (_01975_, _01974_, _05806_);
  or (_01976_, _01975_, _01971_);
  or (_01977_, _01976_, _01970_);
  and (_02466_, _01977_, _05110_);
  and (_02472_, _11976_, _05110_);
  or (_01978_, _01732_, rst);
  nor (_02476_, _01978_, _01893_);
  and (_01979_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_01980_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_02503_, _01980_, _01979_);
  and (_01981_, _06625_, _06122_);
  and (_01982_, _01981_, _08133_);
  nand (_01983_, _01982_, _05872_);
  or (_01984_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01985_, _01984_, _05794_);
  and (_01986_, _01985_, _01983_);
  and (_01987_, _06128_, _05992_);
  not (_01988_, _01987_);
  nor (_01989_, _01988_, _06054_);
  and (_01990_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_01991_, _01990_, _01989_);
  and (_01992_, _01991_, _05806_);
  and (_01993_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_01994_, _01993_, rst);
  or (_01995_, _01994_, _01992_);
  or (_02518_, _01995_, _01986_);
  and (_01996_, _10154_, _05789_);
  and (_01997_, _01996_, _05488_);
  nand (_01998_, _01997_, _05872_);
  or (_01999_, _01997_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02000_, _01999_, _05794_);
  and (_02001_, _02000_, _01998_);
  and (_02002_, _08252_, _05992_);
  nand (_02003_, _02002_, _05841_);
  or (_02004_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02005_, _02004_, _05806_);
  and (_02006_, _02005_, _02003_);
  and (_02007_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_02008_, _02007_, rst);
  or (_02009_, _02008_, _02006_);
  or (_02520_, _02009_, _02001_);
  and (_02011_, _01996_, _08272_);
  nand (_02012_, _02011_, _05872_);
  or (_02013_, _02011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02014_, _02013_, _05794_);
  and (_02015_, _02014_, _02012_);
  nand (_02016_, _02002_, _05938_);
  or (_02017_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02018_, _02017_, _05806_);
  and (_02019_, _02018_, _02016_);
  and (_02020_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_02021_, _02020_, rst);
  or (_02022_, _02021_, _02019_);
  or (_02522_, _02022_, _02015_);
  nand (_02023_, _01174_, _11559_);
  and (_02024_, _02023_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02025_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02026_, _02025_, _08245_);
  and (_02027_, _02026_, _01174_);
  or (_02028_, _02027_, _02024_);
  and (_02029_, _02028_, _05794_);
  nand (_02030_, _01180_, _06229_);
  or (_02031_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02032_, _02031_, _05806_);
  and (_02033_, _02032_, _02030_);
  and (_02034_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02035_, _02034_, rst);
  or (_02036_, _02035_, _02033_);
  or (_02525_, _02036_, _02029_);
  nor (_02037_, _08056_, _06054_);
  and (_02038_, _08117_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_02039_, _02038_, _02037_);
  and (_02543_, _02039_, _05110_);
  and (_02040_, _10154_, _06122_);
  and (_02041_, _02040_, _10208_);
  nand (_02042_, _02041_, _05872_);
  or (_02043_, _02041_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_02044_, _02043_, _05794_);
  and (_02045_, _02044_, _02042_);
  and (_02046_, _06145_, _05992_);
  not (_02047_, _02046_);
  nor (_02049_, _02047_, _05334_);
  and (_02050_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02051_, _02050_, _02049_);
  and (_02052_, _02051_, _05806_);
  and (_02053_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02054_, _02053_, rst);
  or (_02055_, _02054_, _02052_);
  or (_02547_, _02055_, _02045_);
  and (_02056_, _01981_, _10208_);
  nand (_02057_, _02056_, _05872_);
  or (_02058_, _02056_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_02059_, _02058_, _05794_);
  and (_02060_, _02059_, _02057_);
  nor (_02061_, _01988_, _05334_);
  and (_02062_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_02063_, _02062_, _02061_);
  and (_02064_, _02063_, _05806_);
  and (_02065_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_02066_, _02065_, rst);
  or (_02067_, _02066_, _02064_);
  or (_02549_, _02067_, _02060_);
  and (_02068_, _01996_, _08133_);
  nand (_02069_, _02068_, _05872_);
  or (_02070_, _02068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02071_, _02070_, _05794_);
  and (_02072_, _02071_, _02069_);
  nand (_02073_, _02002_, _06054_);
  or (_02074_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02075_, _02074_, _05806_);
  and (_02076_, _02075_, _02073_);
  and (_02077_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_02078_, _02077_, rst);
  or (_02079_, _02078_, _02076_);
  or (_02553_, _02079_, _02072_);
  not (_02080_, _02002_);
  or (_02081_, _02080_, _05782_);
  or (_02082_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_02083_, _02082_, _05794_);
  and (_02084_, _02083_, _02081_);
  nand (_02085_, _02002_, _06798_);
  and (_02087_, _02082_, _05806_);
  and (_02088_, _02087_, _02085_);
  not (_02089_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_02090_, _05793_, _02089_);
  or (_02091_, _02090_, rst);
  or (_02092_, _02091_, _02088_);
  or (_02555_, _02092_, _02084_);
  and (_02093_, _01996_, _06631_);
  nand (_02094_, _02093_, _05872_);
  or (_02095_, _02093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02096_, _02095_, _05794_);
  and (_02097_, _02096_, _02094_);
  nand (_02098_, _02002_, _06088_);
  or (_02099_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02100_, _02099_, _05806_);
  and (_02101_, _02100_, _02098_);
  and (_02102_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_02103_, _02102_, rst);
  or (_02104_, _02103_, _02101_);
  or (_02557_, _02104_, _02097_);
  and (_02105_, _01174_, _05488_);
  nand (_02106_, _02105_, _05872_);
  or (_02107_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02108_, _02107_, _05794_);
  and (_02109_, _02108_, _02106_);
  nand (_02110_, _01180_, _05841_);
  or (_02111_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02112_, _02111_, _05806_);
  and (_02113_, _02112_, _02110_);
  and (_02114_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_02115_, _02114_, rst);
  or (_02116_, _02115_, _02113_);
  or (_02559_, _02116_, _02109_);
  and (_02117_, _05804_, _05996_);
  nand (_02118_, _02117_, _05872_);
  or (_02119_, _02117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02120_, _02119_, _05794_);
  and (_02121_, _02120_, _02118_);
  nand (_02122_, _01180_, _05938_);
  or (_02123_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02124_, _02123_, _05806_);
  and (_02125_, _02124_, _02122_);
  and (_02126_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_02127_, _02126_, rst);
  or (_02128_, _02127_, _02125_);
  or (_02562_, _02128_, _02121_);
  and (_02129_, _01174_, _10208_);
  nand (_02130_, _02129_, _05872_);
  or (_02131_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02132_, _02131_, _05794_);
  and (_02133_, _02132_, _02130_);
  nand (_02134_, _01180_, _05334_);
  or (_02135_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02136_, _02135_, _05806_);
  and (_02137_, _02136_, _02134_);
  and (_02138_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_02139_, _02138_, rst);
  or (_02140_, _02139_, _02137_);
  or (_02565_, _02140_, _02133_);
  nand (_02141_, _06560_, _06054_);
  or (_02142_, _06560_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_02143_, _02142_, _05110_);
  and (_02578_, _02143_, _02141_);
  or (_02144_, _07141_, _07125_);
  and (_02145_, _02144_, _05474_);
  and (_02146_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02147_, _02146_, _07150_);
  or (_02148_, _02147_, _02145_);
  and (_02587_, _02148_, _05110_);
  and (_02602_, _11954_, _05110_);
  and (_02149_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02150_, _02149_, _07149_);
  and (_02151_, _02150_, _05110_);
  and (_02152_, _07116_, _06277_);
  or (_02153_, _06868_, _07065_);
  or (_02154_, _02153_, _07134_);
  or (_02155_, _02154_, _02152_);
  and (_02156_, _02155_, _06842_);
  or (_02607_, _02156_, _02151_);
  not (_02157_, _08253_);
  and (_02158_, _08243_, _05867_);
  or (_02159_, _02158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_02160_, _02159_, _02157_);
  nand (_02161_, _02158_, _05872_);
  and (_02162_, _02161_, _02160_);
  nor (_02163_, _02157_, _05901_);
  or (_02164_, _02163_, _02162_);
  and (_02626_, _02164_, _05110_);
  and (_02165_, _01981_, _06631_);
  nand (_02166_, _02165_, _05872_);
  or (_02167_, _02165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_02168_, _02167_, _05794_);
  and (_02169_, _02168_, _02166_);
  nor (_02170_, _01988_, _06088_);
  and (_02171_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_02172_, _02171_, _02170_);
  and (_02173_, _02172_, _05806_);
  and (_02174_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_02175_, _02174_, rst);
  or (_02176_, _02175_, _02173_);
  or (_02655_, _02176_, _02169_);
  and (_02177_, _01981_, _06472_);
  nand (_02178_, _02177_, _05872_);
  or (_02179_, _02177_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_02180_, _02179_, _05794_);
  and (_02181_, _02180_, _02178_);
  nor (_02182_, _01988_, _06229_);
  and (_02183_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02184_, _02183_, _02182_);
  and (_02185_, _02184_, _05806_);
  and (_02186_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02187_, _02186_, rst);
  or (_02188_, _02187_, _02185_);
  or (_02656_, _02188_, _02181_);
  and (_02189_, _01981_, _08272_);
  nand (_02190_, _02189_, _05872_);
  or (_02191_, _02189_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_02192_, _02191_, _05794_);
  and (_02193_, _02192_, _02190_);
  nor (_02194_, _01988_, _05938_);
  and (_02195_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_02196_, _02195_, _02194_);
  and (_02197_, _02196_, _05806_);
  and (_02198_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_02199_, _02198_, rst);
  or (_02200_, _02199_, _02197_);
  or (_02666_, _02200_, _02193_);
  and (_02201_, _02040_, _06472_);
  nand (_02202_, _02201_, _05872_);
  or (_02203_, _02201_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_02204_, _02203_, _05794_);
  and (_02205_, _02204_, _02202_);
  nor (_02206_, _02047_, _06229_);
  and (_02208_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02209_, _02208_, _02206_);
  and (_02210_, _02209_, _05806_);
  and (_02211_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02212_, _02211_, rst);
  or (_02213_, _02212_, _02210_);
  or (_02668_, _02213_, _02205_);
  and (_02214_, _02040_, _08272_);
  nand (_02215_, _02214_, _05872_);
  or (_02216_, _02214_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_02217_, _02216_, _05794_);
  and (_02219_, _02217_, _02215_);
  nor (_02220_, _02047_, _05938_);
  and (_02221_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_02223_, _02221_, _02220_);
  and (_02224_, _02223_, _05806_);
  and (_02225_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_02226_, _02225_, rst);
  or (_02227_, _02226_, _02224_);
  or (_02671_, _02227_, _02219_);
  and (_02228_, _02040_, _05488_);
  nand (_02229_, _02228_, _05872_);
  or (_02230_, _02228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_02231_, _02230_, _05794_);
  and (_02232_, _02231_, _02229_);
  nor (_02233_, _02047_, _05841_);
  and (_02234_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02235_, _02234_, _02233_);
  and (_02236_, _02235_, _05806_);
  and (_02237_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02238_, _02237_, rst);
  or (_02239_, _02238_, _02236_);
  or (_02677_, _02239_, _02232_);
  or (_02240_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_02241_, _02240_, _05110_);
  nand (_02242_, _08257_, _05901_);
  and (_02688_, _02242_, _02241_);
  nand (_02243_, _01174_, _05805_);
  or (_02244_, _02243_, _05782_);
  or (_02245_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_02246_, _02245_, _05794_);
  and (_02247_, _02246_, _02244_);
  nand (_02248_, _01180_, _06798_);
  and (_02249_, _02245_, _05806_);
  and (_02250_, _02249_, _02248_);
  not (_02251_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_02252_, _05793_, _02251_);
  or (_02253_, _02252_, rst);
  or (_02254_, _02253_, _02250_);
  or (_02690_, _02254_, _02247_);
  and (_02256_, _01174_, _08133_);
  nand (_02257_, _02256_, _05872_);
  or (_02258_, _02256_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_02259_, _02258_, _05794_);
  and (_02260_, _02259_, _02257_);
  nand (_02261_, _01180_, _06054_);
  or (_02262_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_02263_, _02262_, _05806_);
  and (_02264_, _02263_, _02261_);
  and (_02265_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_02266_, _02265_, rst);
  or (_02267_, _02266_, _02264_);
  or (_02692_, _02267_, _02260_);
  and (_02268_, _01174_, _06631_);
  nand (_02269_, _02268_, _05872_);
  or (_02270_, _02268_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02271_, _02270_, _05794_);
  and (_02272_, _02271_, _02269_);
  nand (_02273_, _01180_, _06088_);
  or (_02274_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02275_, _02274_, _05806_);
  and (_02276_, _02275_, _02273_);
  and (_02277_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_02278_, _02277_, rst);
  or (_02279_, _02278_, _02276_);
  or (_02694_, _02279_, _02272_);
  or (_02280_, _01988_, _05782_);
  or (_02281_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_02282_, _02281_, _05794_);
  and (_02283_, _02282_, _02280_);
  and (_02284_, _01987_, _06799_);
  not (_02285_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_02286_, _01987_, _02285_);
  or (_02287_, _02286_, _02284_);
  and (_02288_, _02287_, _05806_);
  nor (_02289_, _05793_, _02285_);
  or (_02290_, _02289_, rst);
  or (_02291_, _02290_, _02288_);
  or (_02696_, _02291_, _02283_);
  and (_02292_, _01996_, _10208_);
  nand (_02293_, _02292_, _05872_);
  or (_02294_, _02292_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02295_, _02294_, _05794_);
  and (_02296_, _02295_, _02293_);
  nand (_02297_, _02002_, _05334_);
  or (_02298_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02299_, _02298_, _05806_);
  and (_02300_, _02299_, _02297_);
  and (_02301_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_02302_, _02301_, rst);
  or (_02303_, _02302_, _02300_);
  or (_02698_, _02303_, _02296_);
  and (_02304_, _01996_, _06472_);
  nand (_02305_, _02304_, _05872_);
  or (_02306_, _02304_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02307_, _02306_, _05794_);
  and (_02308_, _02307_, _02305_);
  nand (_02309_, _02002_, _06229_);
  or (_02310_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_02311_, _02310_, _05806_);
  and (_02312_, _02311_, _02309_);
  and (_02313_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_02314_, _02313_, rst);
  or (_02315_, _02314_, _02312_);
  or (_02700_, _02315_, _02308_);
  nand (_02316_, _02040_, _05805_);
  or (_02317_, _02316_, _05782_);
  or (_02318_, _02046_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_02319_, _02318_, _05794_);
  and (_02320_, _02319_, _02317_);
  nand (_02321_, _02046_, _06798_);
  and (_02322_, _02318_, _05806_);
  and (_02323_, _02322_, _02321_);
  not (_02324_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_02325_, _05793_, _02324_);
  or (_02326_, _02325_, rst);
  or (_02327_, _02326_, _02323_);
  or (_02702_, _02327_, _02320_);
  and (_02328_, _01981_, _05488_);
  nand (_02329_, _02328_, _05872_);
  or (_02330_, _02328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_02331_, _02330_, _05794_);
  and (_02332_, _02331_, _02329_);
  nor (_02333_, _01988_, _05841_);
  and (_02334_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02335_, _02334_, _02333_);
  and (_02336_, _02335_, _05806_);
  and (_02337_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02338_, _02337_, rst);
  or (_02339_, _02338_, _02336_);
  or (_02704_, _02339_, _02332_);
  and (_02340_, _02040_, _08133_);
  nand (_02341_, _02340_, _05872_);
  or (_02342_, _02340_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_02343_, _02342_, _05794_);
  and (_02344_, _02343_, _02341_);
  nor (_02345_, _02047_, _06054_);
  and (_02346_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_02347_, _02346_, _02345_);
  and (_02348_, _02347_, _05806_);
  and (_02349_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_02350_, _02349_, rst);
  or (_02351_, _02350_, _02348_);
  or (_02707_, _02351_, _02344_);
  and (_02352_, _02040_, _06631_);
  nand (_02353_, _02352_, _05872_);
  or (_02354_, _02352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_02355_, _02354_, _05794_);
  and (_02356_, _02355_, _02353_);
  nor (_02357_, _02047_, _06088_);
  and (_02358_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_02359_, _02358_, _02357_);
  and (_02360_, _02359_, _05806_);
  and (_02361_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_02362_, _02361_, rst);
  or (_02363_, _02362_, _02360_);
  or (_02709_, _02363_, _02356_);
  and (_02364_, _07034_, _05997_);
  nand (_02365_, _05997_, _05337_);
  and (_02366_, _02365_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_02367_, _02366_, _02364_);
  and (_02738_, _02367_, _05110_);
  and (_02368_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_02369_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_02370_, pc_log_change, _02369_);
  or (_02371_, _02370_, _02368_);
  and (_02755_, _02371_, _05110_);
  or (_02372_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not (_02373_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_02374_, pc_log_change, _02373_);
  and (_02375_, _02374_, _05110_);
  and (_02759_, _02375_, _02372_);
  or (_02376_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not (_02377_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_02378_, pc_log_change, _02377_);
  and (_02379_, _02378_, _05110_);
  and (_02762_, _02379_, _02376_);
  and (_02380_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_02381_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_02382_, pc_log_change, _02381_);
  or (_02383_, _02382_, _02380_);
  and (_02763_, _02383_, _05110_);
  and (_02384_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_02385_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_02386_, pc_log_change, _02385_);
  or (_02387_, _02386_, _02384_);
  and (_02771_, _02387_, _05110_);
  or (_02388_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_02389_, pc_log_change, _05264_);
  and (_02390_, _02389_, _05110_);
  and (_02774_, _02390_, _02388_);
  and (_02392_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_02393_, pc_log_change, _06162_);
  or (_02394_, _02393_, _02392_);
  and (_02776_, _02394_, _05110_);
  and (_02395_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_02396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_02397_, pc_log_change, _02396_);
  or (_02398_, _02397_, _02395_);
  and (_02780_, _02398_, _05110_);
  or (_02399_, _01668_, _07093_);
  and (_02400_, _06463_, _06434_);
  or (_02401_, _07052_, _02400_);
  or (_02402_, _02401_, _02399_);
  or (_02403_, _06849_, _06435_);
  and (_02404_, _11727_, _06464_);
  or (_02405_, _02404_, _02403_);
  and (_02406_, _07139_, _11802_);
  or (_02408_, _02406_, _12156_);
  and (_02409_, _07107_, _06852_);
  and (_02410_, _11729_, _06464_);
  or (_02411_, _02410_, _02409_);
  or (_02412_, _02411_, _02408_);
  or (_02413_, _02412_, _02405_);
  or (_02414_, _02413_, _02402_);
  or (_02415_, _13078_, _12134_);
  or (_02416_, _01664_, _06439_);
  or (_02417_, _02416_, _01648_);
  or (_02418_, _02417_, _02415_);
  or (_02419_, _07126_, _07089_);
  or (_02420_, _02419_, _07041_);
  or (_02421_, _07131_, _07106_);
  or (_02422_, _02421_, _02420_);
  or (_02424_, _01665_, _06867_);
  or (_02425_, _01670_, _01712_);
  or (_02426_, _02425_, _02424_);
  or (_02427_, _02426_, _01650_);
  or (_02428_, _02427_, _02422_);
  or (_02429_, _02428_, _02418_);
  or (_02430_, _02429_, _02414_);
  and (_02431_, _02430_, _05474_);
  and (_02432_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_02433_, _00489_);
  and (_02434_, _02433_, _06240_);
  or (_02435_, _07056_, _02434_);
  or (_02436_, _02435_, _02432_);
  or (_02437_, _02436_, _02431_);
  and (_02812_, _02437_, _05110_);
  or (_02438_, _06453_, _06435_);
  or (_02439_, _02438_, _07139_);
  or (_02440_, _07108_, _07041_);
  or (_02441_, _02440_, _02439_);
  or (_02442_, _02441_, _01650_);
  or (_02443_, _11756_, _11297_);
  and (_02444_, _13086_, _06827_);
  and (_02445_, _12149_, _06448_);
  or (_02446_, _02445_, _02444_);
  or (_02447_, _02446_, _02443_);
  or (_02448_, _02447_, _02402_);
  or (_02449_, _02448_, _02442_);
  or (_02450_, _02449_, _02418_);
  and (_02451_, _02450_, _05474_);
  and (_02452_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02453_, _02452_, _02435_);
  or (_02454_, _02453_, _02451_);
  and (_02814_, _02454_, _05110_);
  and (_02455_, _06901_, _08224_);
  and (_02456_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_02457_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_02458_, _02457_, _06011_);
  or (_02459_, _02458_, _02456_);
  or (_02460_, _02459_, _02455_);
  and (_02820_, _02460_, _05110_);
  or (_02461_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not (_02462_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_02464_, pc_log_change, _02462_);
  and (_02465_, _02464_, _05110_);
  and (_02825_, _02465_, _02461_);
  and (_02467_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_02468_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_02469_, pc_log_change, _02468_);
  or (_02470_, _02469_, _02467_);
  and (_02828_, _02470_, _05110_);
  or (_02471_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand (_02473_, _06205_, _07553_);
  and (_02474_, _02473_, _05110_);
  and (_02834_, _02474_, _02471_);
  and (_02475_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_02477_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_02478_, pc_log_change, _02477_);
  or (_02479_, _02478_, _02475_);
  and (_02837_, _02479_, _05110_);
  and (_02480_, _06807_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_02481_, _06825_, _06448_);
  or (_02482_, _02481_, _01645_);
  or (_02483_, _02482_, _11738_);
  or (_02484_, _02483_, _06951_);
  and (_02485_, _06820_, _06448_);
  or (_02486_, _02485_, _06939_);
  or (_02487_, _11742_, _11754_);
  or (_02488_, _02487_, _02486_);
  or (_02489_, _07045_, _06458_);
  or (_02490_, _02489_, _02404_);
  and (_02491_, _11727_, _06448_);
  and (_02492_, _07044_, _06276_);
  or (_02493_, _02492_, _02491_);
  or (_02494_, _02493_, _02490_);
  and (_02495_, _11727_, _06431_);
  or (_02496_, _02495_, _07041_);
  or (_02497_, _07111_, _07052_);
  or (_02498_, _02497_, _02496_);
  or (_02499_, _02498_, _02494_);
  or (_02500_, _02499_, _02488_);
  or (_02501_, _02500_, _02484_);
  and (_02502_, _02501_, _06842_);
  or (_02848_, _02502_, _02480_);
  and (_02504_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not (_02505_, pc_log_change);
  and (_02506_, _02505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02507_, _02506_, _02504_);
  and (_02850_, _02507_, _05110_);
  or (_02508_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not (_02509_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_02510_, pc_log_change, _02509_);
  and (_02511_, _02510_, _05110_);
  and (_02861_, _02511_, _02508_);
  and (_02512_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_02513_, pc_log_change, _02509_);
  or (_02514_, _02513_, _02512_);
  and (_02863_, _02514_, _05110_);
  or (_02515_, _06461_, _06457_);
  or (_02516_, _07081_, _06465_);
  or (_02517_, _02516_, _02515_);
  or (_02519_, _11293_, _06449_);
  or (_02521_, _02519_, _02517_);
  and (_02523_, _07080_, _06460_);
  or (_02524_, _01668_, _01645_);
  nor (_02526_, _02524_, _02523_);
  nand (_02527_, _02526_, _01836_);
  or (_02528_, _02527_, _02521_);
  or (_02529_, _02491_, _02485_);
  or (_02530_, _02410_, _12156_);
  or (_02531_, _02530_, _02529_);
  or (_02532_, _02531_, _07091_);
  or (_02533_, _02532_, _02405_);
  or (_02534_, _02533_, _02528_);
  and (_02535_, _02534_, _06842_);
  nor (_02536_, _06870_, rst);
  and (_02537_, _02536_, _06435_);
  and (_02538_, _06807_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_02539_, _02538_, _02537_);
  or (_02875_, _02539_, _02535_);
  nand (_02540_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02541_, _02540_, _08274_);
  and (_02542_, _08274_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_02544_, _02542_, _02541_);
  and (_02878_, _02544_, _05110_);
  nand (_02545_, _01836_, _11299_);
  or (_02546_, _01667_, _07092_);
  or (_02548_, _02546_, _02415_);
  or (_02550_, _02548_, _02545_);
  and (_02551_, _07038_, _06448_);
  or (_02552_, _02489_, _01649_);
  or (_02554_, _02552_, _02551_);
  or (_02556_, _07052_, _06828_);
  or (_02558_, _11737_, _07097_);
  or (_02560_, _02558_, _02556_);
  or (_02561_, _02560_, _02554_);
  or (_02563_, _01664_, _07121_);
  or (_02564_, _02563_, _02481_);
  or (_02566_, _02564_, _06822_);
  or (_02567_, _02566_, _02561_);
  or (_02568_, _02567_, _02550_);
  and (_02569_, _02568_, _05474_);
  and (_02570_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_02571_, _06435_, _05151_);
  or (_02572_, _02571_, _02570_);
  or (_02573_, _02572_, _02569_);
  and (_02881_, _02573_, _05110_);
  and (_02574_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_02575_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_02576_, _02575_, _02574_);
  and (_02885_, _02576_, _05110_);
  and (_02577_, _06807_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  or (_02579_, _06460_, _06448_);
  and (_02580_, _02579_, _06814_);
  or (_02581_, _02546_, _02487_);
  or (_02582_, _02581_, _02580_);
  or (_02583_, _01649_, _06462_);
  and (_02584_, _06946_, _06810_);
  or (_02585_, _01647_, _02584_);
  or (_02586_, _02585_, _02583_);
  or (_02588_, _12089_, _06439_);
  or (_02589_, _01665_, _07139_);
  or (_02590_, _02589_, _02588_);
  or (_02591_, _02590_, _06819_);
  or (_02592_, _02591_, _02586_);
  or (_02593_, _02592_, _02564_);
  or (_02594_, _02593_, _02582_);
  or (_02595_, _06439_, _05473_);
  nor (_02596_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and (_02597_, _02596_, _02595_);
  and (_02598_, _02597_, _02594_);
  or (_02894_, _02598_, _02577_);
  or (_02599_, _09328_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_02600_, _09328_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02601_, _02600_, _02599_);
  nand (_02603_, _02601_, _05110_);
  nor (_02897_, _02603_, _08274_);
  nor (_02604_, _05901_, _06010_);
  and (_02605_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_02606_, _02605_, _05995_);
  or (_02608_, _02606_, _02604_);
  or (_02609_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02610_, _02609_, _05110_);
  and (_02906_, _02610_, _02608_);
  nand (_02611_, _06673_, _05901_);
  or (_02612_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02613_, _02612_, _05110_);
  and (_02917_, _02613_, _02611_);
  and (_02614_, _01996_, _05867_);
  nand (_02615_, _02614_, _05872_);
  or (_02616_, _02614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_02617_, _02616_, _05794_);
  and (_02618_, _02617_, _02615_);
  nand (_02619_, _02002_, _05901_);
  or (_02620_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_02621_, _02620_, _05806_);
  and (_02622_, _02621_, _02619_);
  and (_02623_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_02624_, _02623_, rst);
  or (_02625_, _02624_, _02622_);
  or (_02921_, _02625_, _02618_);
  nand (_02627_, _06673_, _05841_);
  or (_02628_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02629_, _02628_, _05110_);
  and (_02925_, _02629_, _02627_);
  and (_02630_, _06807_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_02631_, _02556_, _11738_);
  or (_02632_, _02631_, _02482_);
  or (_02633_, _12134_, _11761_);
  or (_02634_, _13072_, _02491_);
  or (_02635_, _02634_, _02633_);
  or (_02636_, _02635_, _07050_);
  or (_02637_, _02636_, _02488_);
  or (_02638_, _02637_, _02632_);
  and (_02639_, _02638_, _06842_);
  or (_02940_, _02639_, _02630_);
  or (_02640_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_02641_, _06205_, _12002_);
  and (_02642_, _02641_, _05110_);
  and (_02946_, _02642_, _02640_);
  and (_02948_, _01725_, _05110_);
  nand (_02643_, _06560_, _06088_);
  or (_02644_, _06560_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_02645_, _02644_, _05110_);
  and (_02954_, _02645_, _02643_);
  and (_02646_, _06901_, _12894_);
  and (_02647_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_02648_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_02649_, _02648_, _06011_);
  or (_02650_, _02649_, _02647_);
  or (_02651_, _02650_, _02646_);
  and (_02963_, _02651_, _05110_);
  and (_02652_, _08056_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_02653_, _08056_, _05901_);
  or (_02654_, _02653_, _02652_);
  and (_02970_, _02654_, _05110_);
  or (_02657_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_02658_, _06205_, _13066_);
  and (_02659_, _02658_, _05110_);
  and (_03001_, _02659_, _02657_);
  and (_02660_, _08056_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_02661_, _07034_, _06001_);
  or (_02662_, _02661_, _02660_);
  and (_03033_, _02662_, _05110_);
  nor (_02663_, _01320_, _05841_);
  and (_02664_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_02665_, _02664_, _02663_);
  and (_03057_, _02665_, _05110_);
  and (_02667_, _12841_, _08280_);
  and (_02669_, _08286_, _12828_);
  and (_02670_, _02669_, _12841_);
  not (_02672_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_02673_, _08286_, _02672_);
  or (_02674_, _02673_, _02670_);
  and (_02675_, _02674_, _08282_);
  nand (_02676_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02678_, _02676_, _08281_);
  nor (_02679_, _02678_, _02675_);
  nor (_02680_, _02679_, _08280_);
  or (_02681_, _02680_, _02667_);
  nand (_02682_, _02681_, _05110_);
  nor (_03059_, _02682_, _08274_);
  and (_03064_, _11832_, _05110_);
  and (_03073_, _12252_, _05110_);
  and (_03075_, _12220_, _05110_);
  nand (_02683_, _02670_, _08281_);
  nand (_02684_, _02683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02685_, _02684_, _02667_);
  or (_02686_, _02685_, _08274_);
  and (_03085_, _02686_, _05110_);
  and (_03089_, _12291_, _05110_);
  nor (_03101_, _12014_, rst);
  and (_02687_, _10641_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_03108_, _02687_, _10460_);
  and (_02689_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_02691_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_03112_, _02691_, _02689_);
  not (_02693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  and (_02695_, _01326_, _02693_);
  and (_02697_, _02695_, _08752_);
  or (_02699_, _02697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not (_02701_, rxd_i);
  nand (_02703_, _02697_, _02701_);
  and (_02705_, _02703_, _05110_);
  and (_03114_, _02705_, _02699_);
  and (_02706_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_02708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05850_);
  nor (_02710_, _02708_, _05987_);
  not (_02711_, _02710_);
  and (_02712_, _02711_, _06099_);
  or (_02713_, _02712_, _05986_);
  or (_02714_, _02713_, _02706_);
  or (_02715_, _02710_, _06137_);
  and (_02716_, _02715_, _05110_);
  and (_03130_, _02716_, _02714_);
  and (_02717_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_02718_, _08235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02719_, _02718_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_02720_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02721_, _02720_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_02722_, _02693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02723_, _02722_, _02721_);
  and (_02724_, _02723_, _08745_);
  nor (_02725_, _02724_, _02719_);
  nor (_02726_, _02725_, _01050_);
  nor (_02727_, _02723_, _01325_);
  and (_02728_, _08742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02729_, _08235_, _01057_);
  and (_02730_, _02729_, _02728_);
  nor (_02731_, _02730_, _08745_);
  not (_02732_, _02731_);
  nor (_02733_, _02732_, _08748_);
  nor (_02734_, _02733_, _02727_);
  not (_02735_, _02719_);
  nand (_02736_, _02735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor (_02737_, _02736_, _02734_);
  or (_02739_, _02737_, _02726_);
  and (_02740_, _02739_, _09325_);
  or (_03135_, _02740_, _02717_);
  not (_02741_, _02725_);
  and (_02742_, _02741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand (_02743_, _02735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_02744_, _02743_, _02734_);
  or (_02745_, _02744_, _02742_);
  and (_02746_, _02745_, _09325_);
  or (_03143_, _02746_, _09324_);
  and (_02747_, _02741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02748_, _02727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_02749_, _08748_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02750_, _02749_, _02731_);
  or (_02751_, _02750_, _02748_);
  and (_02752_, _02751_, _02735_);
  or (_02753_, _02752_, _02747_);
  and (_02754_, _02753_, _09325_);
  or (_03145_, _02754_, _01065_);
  or (_02756_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_02757_, _02756_, _02734_);
  or (_02758_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02760_, _02758_, _09325_);
  and (_02761_, _02760_, _02757_);
  or (_03147_, _02761_, _01195_);
  or (_02764_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_02765_, _02764_, _02734_);
  or (_02766_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02767_, _02766_, _09325_);
  and (_02768_, _02767_, _02765_);
  or (_03149_, _02768_, _01197_);
  or (_02769_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_02770_, _02769_, _02734_);
  or (_02772_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_02773_, _02772_, _09325_);
  and (_02775_, _02773_, _02770_);
  or (_03151_, _02775_, _01199_);
  or (_02777_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_02778_, _02777_, _02734_);
  or (_02779_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02781_, _02779_, _09325_);
  and (_02782_, _02781_, _02778_);
  or (_03153_, _02782_, _01979_);
  not (_02783_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_02784_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not (_02785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_02786_, _05846_, _02785_);
  or (_02787_, _02786_, _11265_);
  nor (_02788_, _02787_, _02784_);
  nand (_02789_, _02788_, _02783_);
  nor (_02790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_02791_, _02790_, _02788_);
  nand (_02792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_02793_, _02792_, _02791_);
  and (_02794_, _02793_, _05110_);
  and (_03155_, _02794_, _02789_);
  or (_02795_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_02796_, _02795_, _02734_);
  or (_02797_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02798_, _02797_, _09325_);
  and (_02799_, _02798_, _02796_);
  or (_03165_, _02799_, _02689_);
  or (_02800_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02801_, _02800_, _02734_);
  and (_02802_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02803_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_02804_, _02803_, _09325_);
  or (_02805_, _02804_, _02802_);
  and (_03167_, _02805_, _02801_);
  or (_02806_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02807_, _02806_, _02734_);
  and (_02808_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02809_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  and (_02810_, _02809_, _09325_);
  or (_02811_, _02810_, _02808_);
  and (_03170_, _02811_, _02807_);
  or (_02813_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02815_, _02813_, _02734_);
  and (_02816_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02817_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and (_02818_, _02817_, _09325_);
  or (_02819_, _02818_, _02816_);
  and (_03173_, _02819_, _02815_);
  and (_03186_, _02791_, _05110_);
  nor (_02821_, _02734_, _01050_);
  and (_02822_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  or (_02823_, _02822_, rxd_i);
  or (_02824_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and (_02826_, _02824_, _02724_);
  or (_02827_, _02826_, _02719_);
  and (_02829_, _02827_, _02823_);
  or (_02830_, _02829_, _02821_);
  nand (_02831_, _02719_, _02701_);
  and (_02832_, _02831_, _09325_);
  and (_02833_, _02832_, _02830_);
  and (_02835_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_03191_, _02835_, _02833_);
  and (_02836_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_03193_, _02836_, _02717_);
  or (_02838_, _12171_, _05782_);
  nor (_02839_, _12172_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_02840_, _02839_, _10157_);
  and (_02841_, _02840_, _02838_);
  or (_02842_, _02841_, _10162_);
  and (_02843_, _12083_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_02844_, _02843_, _01548_);
  and (_02845_, _02844_, _10157_);
  or (_02846_, _02845_, _02842_);
  nand (_02847_, _10162_, _05901_);
  and (_02849_, _02847_, _05110_);
  and (_03196_, _02849_, _02846_);
  and (_03198_, _12049_, _05110_);
  and (_03203_, _11909_, _05110_);
  and (_02851_, _07204_, _06613_);
  nor (_02852_, _10208_, _05142_);
  or (_02853_, _02852_, _10209_);
  and (_02854_, _06638_, _08132_);
  nand (_02855_, _02854_, _02853_);
  nor (_02856_, _07235_, _06622_);
  and (_02857_, _12179_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_02858_, _02857_, _02856_);
  nand (_02859_, _02858_, _02855_);
  and (_02860_, _02859_, _06637_);
  or (_02862_, _02860_, _02851_);
  and (_03309_, _02862_, _05110_);
  and (_02864_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_02865_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_02866_, _02865_, _06011_);
  and (_02867_, _06799_, _06901_);
  or (_02868_, _02867_, _02866_);
  or (_02869_, _02868_, _02864_);
  and (_03316_, _02869_, _05110_);
  or (_02870_, _01327_, _08750_);
  and (_02871_, _02870_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_02872_, _02871_, _02697_);
  and (_03532_, _02872_, _05110_);
  and (_02873_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_02874_, _08617_, _06183_);
  or (_02876_, _02874_, _02873_);
  and (_03534_, _02876_, _05110_);
  not (_02877_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_02879_, _02722_, _08753_);
  and (_02880_, _02879_, _08752_);
  nor (_02882_, _02880_, _02877_);
  and (_02883_, _02880_, rxd_i);
  or (_02884_, _02883_, _02882_);
  and (_03571_, _02884_, _05110_);
  and (_02886_, _01981_, _05867_);
  nand (_02887_, _02886_, _05872_);
  or (_02888_, _02886_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_02889_, _02888_, _05794_);
  and (_02890_, _02889_, _02887_);
  nor (_02891_, _01988_, _05901_);
  and (_02892_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_02893_, _02892_, _02891_);
  and (_02895_, _02893_, _05806_);
  and (_02896_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_02898_, _02896_, rst);
  or (_02899_, _02898_, _02895_);
  or (_03593_, _02899_, _02890_);
  and (_02900_, _02040_, _05867_);
  nand (_02901_, _02900_, _05872_);
  or (_02902_, _02900_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_02903_, _02902_, _05794_);
  and (_02904_, _02903_, _02901_);
  nor (_02905_, _02047_, _05901_);
  and (_02907_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_02908_, _02907_, _02905_);
  and (_02909_, _02908_, _05806_);
  and (_02910_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_02911_, _02910_, rst);
  or (_02912_, _02911_, _02909_);
  or (_03596_, _02912_, _02904_);
  not (_02913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_02914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_02915_, _02914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not (_02916_, _02915_);
  nor (_02918_, _08235_, _08741_);
  and (_02919_, _02918_, _02916_);
  and (_02920_, _02919_, _01325_);
  nor (_02922_, _02920_, _02913_);
  and (_02923_, _02920_, rxd_i);
  or (_02924_, _02923_, rst);
  or (_03599_, _02924_, _02922_);
  nor (_02926_, _08235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_02927_, _02926_, _08745_);
  nor (_02928_, _02724_, _08741_);
  or (_02929_, _02928_, _02927_);
  and (_02930_, _02929_, _02735_);
  nand (_02931_, _02741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_02932_, _02931_, _09325_);
  or (_03659_, _02932_, _02930_);
  or (_02933_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand (_02934_, pc_log_change, _00990_);
  and (_02935_, _02934_, _05110_);
  and (_03660_, _02935_, _02933_);
  and (_02936_, _08617_, _08224_);
  nor (_02937_, _06004_, _05995_);
  or (_02938_, _02937_, _08614_);
  and (_02939_, _02938_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_02941_, _02939_, _02936_);
  and (_03663_, _02941_, _05110_);
  and (_02942_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_02944_, pc_log_change, _02943_);
  or (_02945_, _02944_, _02942_);
  and (_03670_, _02945_, _05110_);
  and (_02947_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_02949_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_02950_, _02949_, _02947_);
  and (_02951_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_02952_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_02953_, _02952_, _02951_);
  or (_02955_, _02953_, _02950_);
  and (_02956_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_02957_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_02958_, _02957_, _02956_);
  and (_02959_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_02960_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_02961_, _02960_, _02959_);
  or (_02962_, _02961_, _02958_);
  or (_02964_, _02962_, _02955_);
  and (_02965_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_02966_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_02967_, _02966_, _02965_);
  and (_02968_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02969_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_02971_, _02969_, _02968_);
  or (_02972_, _02971_, _02967_);
  and (_02973_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_02974_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_02975_, _02974_, _02973_);
  and (_02976_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_02977_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_02978_, _02977_, _02976_);
  or (_02979_, _02978_, _02975_);
  or (_02980_, _02979_, _02972_);
  or (_02981_, _02980_, _02964_);
  and (_02982_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02983_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_02984_, _02983_, _02982_);
  and (_02985_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_02986_, _01819_, _12029_);
  or (_02987_, _02986_, _02985_);
  or (_02988_, _02987_, _02984_);
  or (_02989_, _01846_, p2_in[6]);
  or (_02990_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_02991_, _02990_, _02989_);
  and (_02992_, _02991_, _01853_);
  or (_02993_, _01846_, p3_in[6]);
  or (_02994_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_02995_, _02994_, _02993_);
  and (_02996_, _02995_, _01830_);
  or (_02997_, _02996_, _02992_);
  or (_02998_, _01846_, p1_in[6]);
  or (_02999_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03000_, _02999_, _02998_);
  and (_03002_, _03000_, _01865_);
  or (_03003_, _01846_, p0_in[6]);
  or (_03004_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03005_, _03004_, _03003_);
  and (_03006_, _03005_, _01859_);
  or (_03007_, _03006_, _03002_);
  or (_03008_, _03007_, _02997_);
  or (_03009_, _03008_, _02988_);
  and (_03010_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03011_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_03012_, _03011_, _03010_);
  or (_03013_, _03012_, _03009_);
  or (_03014_, _03013_, _02981_);
  and (_03015_, _03014_, _01893_);
  and (_03016_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_03017_, _03016_, _03015_);
  or (_03018_, _03017_, _01732_);
  nand (_03019_, _01732_, _06780_);
  and (_03020_, _03019_, _05110_);
  and (_03684_, _03020_, _03018_);
  or (_03021_, _02913_, rxd_i);
  nand (_03022_, _03021_, _08746_);
  or (_03023_, _08748_, _08743_);
  and (_03024_, _03023_, _03022_);
  or (_03025_, _02732_, _02718_);
  or (_03026_, _03025_, _03024_);
  and (_03686_, _03026_, _09325_);
  not (_03027_, _06239_);
  and (_03028_, _12095_, _03027_);
  or (_03029_, _11730_, _07111_);
  or (_03030_, _03029_, _11761_);
  or (_03031_, _03030_, _02487_);
  or (_03032_, _03031_, _11740_);
  and (_03034_, _03032_, _06870_);
  or (_03035_, _03034_, _03028_);
  and (_03704_, _03035_, _05110_);
  nor (_03036_, _01722_, rst);
  nand (_03037_, _01721_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03038_, _01721_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03039_, _03038_, _03037_);
  and (_03706_, _03039_, _03036_);
  nor (_03040_, _06229_, _05465_);
  and (_03041_, _08329_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_03042_, _03041_, _03040_);
  and (_03709_, _03042_, _05110_);
  nor (_03724_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  nand (_03043_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_03044_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_03045_, _03044_, _03043_);
  or (_03046_, _01910_, _11600_);
  or (_03047_, _01913_, _06897_);
  and (_03048_, _03047_, _03046_);
  and (_03049_, _03048_, _03045_);
  or (_03050_, _01927_, _11628_);
  or (_03051_, _01925_, _05904_);
  and (_03052_, _03051_, _03050_);
  nand (_03053_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand (_03054_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_03055_, _03054_, _03053_);
  and (_03056_, _03055_, _03052_);
  and (_03058_, _03056_, _03049_);
  or (_03060_, _01936_, _13275_);
  or (_03061_, _01935_, _00059_);
  and (_03062_, _03061_, _03060_);
  nand (_03063_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_03065_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_03066_, _03065_, _03063_);
  and (_03067_, _03066_, _03062_);
  nand (_03068_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_03069_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_03070_, _03069_, _03068_);
  nand (_03071_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_03072_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_03074_, _03072_, _03071_);
  and (_03076_, _03074_, _03070_);
  and (_03077_, _03076_, _03067_);
  and (_03078_, _03077_, _03058_);
  nand (_03079_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_03080_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_03081_, _03080_, _03079_);
  nand (_03082_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_03083_, _12324_);
  nand (_03084_, _01819_, _03083_);
  and (_03086_, _03084_, _03082_);
  and (_03087_, _03086_, _03081_);
  nor (_03088_, _01846_, p3_in[0]);
  and (_03090_, _01846_, _02324_);
  nor (_03091_, _03090_, _03088_);
  nand (_03092_, _03091_, _01830_);
  nor (_03093_, _01846_, p2_in[0]);
  and (_03094_, _01846_, _02285_);
  nor (_03095_, _03094_, _03093_);
  nand (_03096_, _03095_, _01853_);
  and (_03097_, _03096_, _03092_);
  nor (_03098_, _01846_, p0_in[0]);
  and (_03100_, _01846_, _02251_);
  nor (_03102_, _03100_, _03098_);
  nand (_03103_, _03102_, _01859_);
  nor (_03104_, _01846_, p1_in[0]);
  and (_03105_, _01846_, _02089_);
  nor (_03106_, _03105_, _03104_);
  nand (_03107_, _03106_, _01865_);
  and (_03109_, _03107_, _03103_);
  and (_03110_, _03109_, _03097_);
  and (_03111_, _03110_, _03087_);
  and (_03113_, _12179_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_03115_, _06622_, _06512_);
  nor (_03116_, _03115_, _03113_);
  and (_03117_, _03116_, _06637_);
  nor (_03118_, _08272_, _05269_);
  or (_03119_, _03118_, _00998_);
  nand (_03120_, _03119_, _02854_);
  nand (_03121_, _03120_, _03117_);
  or (_03122_, _07364_, _06637_);
  nand (_03123_, _03122_, _03121_);
  nand (_03124_, _03123_, _08312_);
  or (_03125_, _03123_, _08312_);
  nand (_03126_, _03125_, _03124_);
  not (_03127_, _08155_);
  nand (_03128_, _03127_, _06672_);
  or (_03129_, _03127_, _06672_);
  and (_03131_, _03129_, _03128_);
  nand (_03132_, _03131_, _03126_);
  or (_03133_, _03131_, _03126_);
  nand (_03134_, _03133_, _03132_);
  nor (_03136_, _06784_, _06746_);
  nand (_03137_, _08144_, _03136_);
  or (_03138_, _08144_, _03136_);
  and (_03139_, _03138_, _03137_);
  nand (_03140_, _03139_, _03134_);
  or (_03141_, _03139_, _03134_);
  and (_03142_, _03141_, _03140_);
  or (_03144_, _02862_, _07032_);
  nand (_03146_, _02862_, _07032_);
  and (_03148_, _03146_, _03144_);
  nand (_03150_, _03148_, _03142_);
  or (_03152_, _03148_, _03142_);
  nand (_03154_, _03152_, _03150_);
  nand (_03156_, _03154_, _01874_);
  nand (_03157_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_03158_, _03157_, _03156_);
  and (_03159_, _03158_, _03111_);
  nand (_03160_, _03159_, _03078_);
  and (_03161_, _03160_, _01893_);
  and (_03162_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_03163_, _03162_, _01732_);
  or (_03164_, _03163_, _03161_);
  nand (_03166_, _01732_, _07418_);
  and (_03168_, _03166_, _05110_);
  and (_03748_, _03168_, _03164_);
  and (_03169_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_03171_, _08617_, _12874_);
  or (_03172_, _03171_, _03169_);
  and (_03755_, _03172_, _05110_);
  and (_03174_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_03175_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03176_, _03175_, _03174_);
  and (_03177_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_03178_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_03179_, _03178_, _03177_);
  or (_03180_, _03179_, _03176_);
  and (_03181_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_03182_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_03183_, _03182_, _03181_);
  and (_03184_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_03185_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03187_, _03185_, _03184_);
  or (_03188_, _03187_, _03183_);
  or (_03189_, _03188_, _03180_);
  and (_03190_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_03192_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_03194_, _03192_, _03190_);
  and (_03195_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_03197_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_03199_, _03197_, _03195_);
  or (_03200_, _03199_, _03194_);
  and (_03201_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_03202_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03204_, _03202_, _03201_);
  and (_03205_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_03206_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_03207_, _03206_, _03205_);
  or (_03208_, _03207_, _03204_);
  or (_03209_, _03208_, _03200_);
  or (_03210_, _03209_, _03189_);
  and (_03211_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03212_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_03213_, _03212_, _03211_);
  and (_03214_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_03215_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_03216_, _03215_, _03214_);
  and (_03217_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_03218_, _01819_, _12194_);
  or (_03219_, _03218_, _03217_);
  or (_03220_, _03219_, _03216_);
  or (_03221_, _01846_, p3_in[1]);
  or (_03223_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03224_, _03223_, _03221_);
  and (_03225_, _03224_, _01830_);
  or (_03226_, _01846_, p2_in[1]);
  or (_03227_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03228_, _03227_, _03226_);
  and (_03229_, _03228_, _01853_);
  or (_03230_, _03229_, _03225_);
  or (_03231_, _01846_, p1_in[1]);
  or (_03232_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03233_, _03232_, _03231_);
  and (_03234_, _03233_, _01865_);
  or (_03235_, _01846_, p0_in[1]);
  or (_03236_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03237_, _03236_, _03235_);
  and (_03238_, _03237_, _01859_);
  or (_03239_, _03238_, _03234_);
  or (_03240_, _03239_, _03230_);
  or (_03241_, _03240_, _03220_);
  or (_03242_, _03241_, _03213_);
  or (_03243_, _03242_, _03210_);
  and (_03244_, _03243_, _01893_);
  and (_03245_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_03246_, _03245_, _03244_);
  or (_03247_, _03246_, _01732_);
  nand (_03248_, _01732_, _06512_);
  and (_03249_, _03248_, _05110_);
  and (_03766_, _03249_, _03247_);
  or (_03250_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_03251_, _01721_, rst);
  and (_03769_, _03251_, _03250_);
  and (_03252_, _11871_, _11960_);
  and (_03253_, _01815_, _03252_);
  and (_03254_, _03253_, _06617_);
  nor (_03255_, _03254_, _12086_);
  and (_03256_, _01748_, _06183_);
  or (_03257_, _03256_, _12268_);
  and (_03258_, _01737_, _12874_);
  and (_03259_, _01762_, _12894_);
  and (_03260_, _01724_, _08224_);
  or (_03261_, _03260_, _03259_);
  or (_03262_, _03261_, _03258_);
  or (_03263_, _03262_, _03257_);
  and (_03264_, _01748_, _06559_);
  or (_03265_, _03264_, _12270_);
  and (_03266_, _01737_, _06799_);
  and (_03267_, _01762_, _06194_);
  and (_03268_, _01724_, _06230_);
  or (_03269_, _03268_, _03267_);
  or (_03270_, _03269_, _03266_);
  or (_03271_, _03270_, _03265_);
  nand (_03272_, _03271_, _03263_);
  nor (_03273_, _03272_, _03255_);
  or (_03274_, _11873_, _11960_);
  or (_03275_, _03274_, _01903_);
  or (_03276_, _03154_, _12270_);
  or (_03277_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03278_, _03277_, _01737_);
  and (_03279_, _03278_, _03276_);
  and (_03280_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03281_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_03282_, _03281_, _03280_);
  and (_03283_, _03282_, _12270_);
  and (_03284_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_03285_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03286_, _03285_, _03284_);
  and (_03287_, _03286_, _01762_);
  and (_03288_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03289_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03290_, _03289_, _03288_);
  and (_03291_, _03290_, _12268_);
  or (_03292_, _03291_, _03287_);
  or (_03293_, _03292_, _03283_);
  nor (_03294_, _03293_, _03279_);
  nor (_03295_, _03294_, _03275_);
  and (_03296_, _01769_, _11871_);
  or (_03297_, _01846_, p3_in[5]);
  or (_03298_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03299_, _03298_, _03297_);
  and (_03300_, _03299_, _12270_);
  and (_03301_, _03224_, _12268_);
  or (_03302_, _03301_, _03300_);
  and (_03303_, _03302_, _01748_);
  and (_03304_, _01850_, _12270_);
  or (_03305_, _01846_, p3_in[3]);
  or (_03306_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03307_, _03306_, _03305_);
  and (_03308_, _03307_, _12268_);
  or (_03310_, _03308_, _03304_);
  and (_03311_, _03310_, _01762_);
  or (_03312_, _01846_, p3_in[4]);
  or (_03313_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03314_, _03313_, _03312_);
  and (_03315_, _03314_, _12270_);
  and (_03317_, _03091_, _12268_);
  or (_03318_, _03317_, _03315_);
  and (_03319_, _03318_, _01737_);
  and (_03320_, _02995_, _12270_);
  or (_03321_, _01846_, p3_in[2]);
  or (_03322_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03323_, _03322_, _03321_);
  and (_03324_, _03323_, _12268_);
  or (_03325_, _03324_, _03320_);
  and (_03326_, _03325_, _01724_);
  or (_03327_, _03326_, _03319_);
  or (_03328_, _03327_, _03311_);
  or (_03329_, _03328_, _03303_);
  and (_03330_, _03329_, _11958_);
  and (_03331_, _01856_, _12270_);
  or (_03332_, _01846_, p2_in[3]);
  or (_03333_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03334_, _03333_, _03332_);
  and (_03335_, _03334_, _12268_);
  or (_03336_, _03335_, _03331_);
  and (_03337_, _03336_, _01762_);
  or (_03338_, _01846_, p2_in[2]);
  or (_03339_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03340_, _03339_, _03338_);
  or (_03341_, _03340_, _12270_);
  or (_03342_, _02991_, _12268_);
  and (_03343_, _03342_, _03341_);
  and (_03344_, _03343_, _01724_);
  or (_03345_, _01846_, p2_in[4]);
  or (_03346_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03347_, _03346_, _03345_);
  and (_03348_, _03347_, _12270_);
  and (_03349_, _03095_, _12268_);
  or (_03350_, _03349_, _03348_);
  and (_03351_, _03350_, _01737_);
  or (_03352_, _03351_, _03344_);
  or (_03353_, _01846_, p2_in[5]);
  or (_03354_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03355_, _03354_, _03353_);
  and (_03356_, _03355_, _12270_);
  and (_03357_, _03228_, _12268_);
  or (_03358_, _03357_, _03356_);
  and (_03359_, _03358_, _01748_);
  or (_03360_, _03359_, _03352_);
  or (_03361_, _03360_, _03337_);
  and (_03362_, _03361_, _11960_);
  nor (_03363_, _03362_, _03330_);
  nand (_03364_, _03363_, _03296_);
  and (_03365_, _01815_, _11871_);
  nand (_03366_, _03252_, _01727_);
  nand (_03367_, _03275_, _03366_);
  nor (_03368_, _03367_, _03365_);
  nand (_03369_, _01794_, _11871_);
  and (_03370_, _11918_, _12071_);
  and (_03371_, _11873_, _01725_);
  and (_03372_, _03371_, _11960_);
  and (_03373_, _03372_, _03370_);
  or (_03374_, _01918_, _11871_);
  nand (_03375_, _03374_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_03376_, _03375_, _03373_);
  and (_03377_, _03376_, _03369_);
  and (_03378_, _03377_, _03368_);
  or (_03379_, _03378_, _03296_);
  and (_03380_, _03379_, _03364_);
  and (_03381_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03382_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_03383_, _03382_, _03381_);
  and (_03384_, _03383_, _01737_);
  and (_03385_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03386_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_03387_, _03386_, _03385_);
  and (_03388_, _03387_, _01762_);
  or (_03389_, _03388_, _03384_);
  and (_03390_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03391_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03392_, _03391_, _03390_);
  and (_03393_, _03392_, _01724_);
  and (_03394_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_03395_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03396_, _03395_, _03394_);
  and (_03397_, _03396_, _01748_);
  or (_03398_, _03397_, _03393_);
  or (_03399_, _03398_, _03389_);
  and (_03400_, _03399_, _01728_);
  and (_03401_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_03402_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03403_, _03402_, _03401_);
  and (_03404_, _03403_, _01737_);
  and (_03405_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_03406_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_03407_, _03406_, _03405_);
  and (_03408_, _03407_, _01748_);
  or (_03409_, _03408_, _03404_);
  and (_03410_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03411_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03412_, _03411_, _03410_);
  and (_03413_, _03412_, _01724_);
  and (_03414_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03415_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_03416_, _03415_, _03414_);
  and (_03417_, _03416_, _01762_);
  or (_03418_, _03417_, _03413_);
  or (_03419_, _03418_, _03409_);
  and (_03420_, _03419_, _01776_);
  or (_03421_, _03420_, _03400_);
  and (_03422_, _03421_, _11873_);
  and (_03423_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_03424_, _03423_, _12268_);
  and (_03425_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03426_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_03427_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_03428_, _03427_, _03426_);
  or (_03429_, _03428_, _03425_);
  or (_03430_, _03429_, _03424_);
  and (_03431_, _03365_, _11958_);
  and (_03432_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_03433_, _03432_, _12270_);
  and (_03434_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_03435_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_03436_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03437_, _03436_, _03435_);
  or (_03438_, _03437_, _03434_);
  or (_03439_, _03438_, _03433_);
  and (_03440_, _03439_, _03431_);
  and (_03441_, _03440_, _03430_);
  and (_03442_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03443_, _03442_, _12270_);
  and (_03444_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_03445_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_03446_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03447_, _03446_, _03445_);
  or (_03448_, _03447_, _03444_);
  or (_03449_, _03448_, _03443_);
  and (_03450_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03451_, _03450_, _12268_);
  and (_03452_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03453_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03454_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03455_, _03454_, _03453_);
  or (_03456_, _03455_, _03452_);
  or (_03457_, _03456_, _03451_);
  and (_03458_, _03457_, _03253_);
  and (_03459_, _03458_, _03449_);
  or (_03460_, _03459_, _03441_);
  or (_03461_, _03460_, _03422_);
  and (_03462_, _03106_, _01737_);
  or (_03463_, _03462_, _12270_);
  or (_03464_, _01846_, p1_in[3]);
  or (_03465_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03466_, _03465_, _03464_);
  and (_03467_, _03466_, _01762_);
  or (_03468_, _01846_, p1_in[2]);
  or (_03469_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03470_, _03469_, _03468_);
  and (_03471_, _03470_, _01724_);
  and (_03472_, _03233_, _01748_);
  or (_03473_, _03472_, _03471_);
  or (_03474_, _03473_, _03467_);
  or (_03475_, _03474_, _03463_);
  and (_03476_, _03000_, _01724_);
  or (_03477_, _03476_, _12268_);
  or (_03478_, _01846_, p1_in[4]);
  or (_03479_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03480_, _03479_, _03478_);
  and (_03481_, _03480_, _01737_);
  or (_03482_, _01846_, p1_in[5]);
  or (_03483_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03484_, _03483_, _03482_);
  and (_03485_, _03484_, _01748_);
  and (_03486_, _01868_, _01762_);
  or (_03487_, _03486_, _03485_);
  or (_03488_, _03487_, _03481_);
  or (_03489_, _03488_, _03477_);
  and (_03490_, _03489_, _03475_);
  or (_03491_, _03490_, _11873_);
  and (_03492_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03493_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03494_, _03493_, _03492_);
  and (_03495_, _03494_, _01724_);
  and (_03496_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_03497_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_03498_, _03497_, _03496_);
  and (_03499_, _03498_, _01737_);
  or (_03500_, _03499_, _03495_);
  and (_03501_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_03502_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03503_, _03502_, _03501_);
  and (_03504_, _03503_, _01762_);
  or (_03505_, _03504_, _03500_);
  and (_03506_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_03507_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03508_, _03507_, _03506_);
  and (_03509_, _03508_, _01748_);
  or (_03510_, _03509_, _11871_);
  or (_03511_, _03510_, _03505_);
  and (_03512_, _03511_, _01794_);
  and (_03513_, _03512_, _03491_);
  nand (_03514_, _12338_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_03515_, _01770_, _11873_);
  and (_03516_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_03517_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_03518_, _03517_, _03516_);
  and (_03519_, _03518_, _01737_);
  and (_03520_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_03521_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03522_, _03521_, _03520_);
  and (_03523_, _03522_, _01748_);
  or (_03524_, _03523_, _03519_);
  and (_03525_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03526_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03527_, _03526_, _03525_);
  and (_03528_, _03527_, _01724_);
  and (_03529_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03530_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03531_, _03530_, _03529_);
  and (_03533_, _03531_, _01762_);
  or (_03535_, _03533_, _03528_);
  or (_03536_, _03535_, _03524_);
  and (_03537_, _03536_, _03515_);
  and (_03538_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_03539_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03540_, _03539_, _03538_);
  and (_03541_, _03540_, _01724_);
  and (_03542_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_03543_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03544_, _03543_, _03542_);
  and (_03545_, _03544_, _01748_);
  or (_03546_, _03545_, _03541_);
  and (_03547_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03548_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_03549_, _03548_, _03547_);
  and (_03550_, _03549_, _01737_);
  and (_03551_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03552_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_03553_, _03552_, _03551_);
  and (_03554_, _03553_, _01762_);
  or (_03555_, _03554_, _03550_);
  or (_03556_, _03555_, _03546_);
  and (_03557_, _03556_, _03373_);
  or (_03558_, _01846_, p0_in[4]);
  or (_03559_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03560_, _03559_, _03558_);
  and (_03561_, _03560_, _12270_);
  and (_03562_, _03102_, _12268_);
  or (_03563_, _03562_, _03561_);
  and (_03564_, _03563_, _01737_);
  and (_03565_, _01863_, _12270_);
  or (_03566_, _01846_, p0_in[3]);
  or (_03567_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03568_, _03567_, _03566_);
  and (_03569_, _03568_, _12268_);
  or (_03570_, _03569_, _03565_);
  and (_03572_, _03570_, _01762_);
  or (_03573_, _03572_, _03564_);
  and (_03574_, _03005_, _12270_);
  or (_03575_, _01846_, p0_in[2]);
  or (_03576_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03577_, _03576_, _03575_);
  and (_03578_, _03577_, _12268_);
  or (_03579_, _03578_, _03574_);
  and (_03580_, _03579_, _01724_);
  or (_03581_, _01846_, p0_in[5]);
  or (_03582_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03583_, _03582_, _03581_);
  and (_03584_, _03583_, _12270_);
  and (_03585_, _03237_, _12268_);
  or (_03586_, _03585_, _03584_);
  and (_03587_, _03586_, _01748_);
  or (_03588_, _03587_, _03580_);
  nor (_03589_, _03588_, _03573_);
  nor (_03590_, _03589_, _03366_);
  or (_03591_, _03590_, _03557_);
  nor (_03592_, _03591_, _03537_);
  nand (_03594_, _03592_, _03514_);
  or (_03595_, _03594_, _03513_);
  or (_03597_, _03595_, _03461_);
  or (_03598_, _03597_, _03380_);
  or (_03600_, _03598_, _03295_);
  or (_03601_, _03514_, _05782_);
  and (_03602_, _03601_, _03255_);
  and (_03603_, _03602_, _03600_);
  or (_03604_, _03603_, _03273_);
  and (_03797_, _03604_, _05110_);
  and (_03605_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_03606_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or (_03607_, _03606_, _03605_);
  and (_03834_, _03607_, _05110_);
  or (_03608_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_03609_, _06205_, _12984_);
  and (_03610_, _03609_, _05110_);
  and (_03849_, _03610_, _03608_);
  and (_03611_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_03612_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or (_03613_, _03612_, _03611_);
  and (_03857_, _03613_, _05110_);
  nor (_03614_, _01721_, _01720_);
  or (_03615_, _03614_, _01722_);
  and (_03616_, _03037_, _05110_);
  and (_03866_, _03616_, _03615_);
  and (_03617_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_03618_, pc_log_change, _01639_);
  or (_03619_, _03618_, _03617_);
  and (_03868_, _03619_, _05110_);
  nor (_03877_, _03123_, rst);
  or (_03620_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_03621_, _06205_, _13092_);
  and (_03622_, _03621_, _05110_);
  and (_03895_, _03622_, _03620_);
  and (_03623_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_03624_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  or (_03625_, _03624_, _03623_);
  and (_03899_, _03625_, _05110_);
  and (_03626_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_03627_, _07034_, _06002_);
  or (_03628_, _03627_, _03626_);
  and (_03907_, _03628_, _05110_);
  and (_03629_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_03630_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or (_03631_, _03630_, _03629_);
  and (_03910_, _03631_, _05110_);
  and (_03632_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_03633_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or (_03634_, _03633_, _03632_);
  and (_03912_, _03634_, _05110_);
  or (_03635_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_03636_, _06205_, _12904_);
  and (_03637_, _03636_, _05110_);
  and (_03914_, _03637_, _03635_);
  nand (_03638_, _06798_, _06673_);
  or (_03639_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03640_, _03639_, _03638_);
  and (_03919_, _03640_, _05110_);
  nand (_03641_, _00531_, _07028_);
  or (_03642_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03643_, _03642_, _05806_);
  and (_03644_, _03643_, _03641_);
  and (_03645_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03646_, _00523_, _05867_);
  nand (_03647_, _03646_, _05872_);
  or (_03648_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03649_, _03648_, _05794_);
  and (_03650_, _03649_, _03647_);
  or (_03651_, _03650_, _03645_);
  or (_03652_, _03651_, _03644_);
  and (_03929_, _03652_, _05110_);
  nor (_03653_, _08056_, _05841_);
  and (_03654_, _08117_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_03655_, _03654_, _03653_);
  and (_03972_, _03655_, _05110_);
  nor (_03656_, _01320_, _05334_);
  and (_03657_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_03658_, _03657_, _03656_);
  and (_03985_, _03658_, _05110_);
  and (_03661_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_03662_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_03664_, _03662_, _03661_);
  and (_03665_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_03666_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_03667_, _03666_, _03665_);
  or (_03668_, _03667_, _03664_);
  and (_03669_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03671_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_03672_, _03671_, _03669_);
  and (_03673_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03674_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03675_, _03674_, _03673_);
  or (_03676_, _03675_, _03672_);
  or (_03677_, _03676_, _03668_);
  and (_03678_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_03679_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_03680_, _03679_, _03678_);
  and (_03681_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_03682_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_03683_, _03682_, _03681_);
  or (_03685_, _03683_, _03680_);
  and (_03687_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_03688_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03689_, _03688_, _03687_);
  and (_03690_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_03691_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_03692_, _03691_, _03690_);
  or (_03693_, _03692_, _03689_);
  or (_03694_, _03693_, _03685_);
  or (_03695_, _03694_, _03677_);
  and (_03696_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_03697_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03698_, _03697_, _03696_);
  and (_03699_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_03700_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_03701_, _03700_, _03699_);
  and (_03702_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_03703_, _11866_);
  and (_03705_, _01819_, _03703_);
  or (_03707_, _03705_, _03702_);
  or (_03708_, _03707_, _03701_);
  and (_03710_, _03334_, _01853_);
  and (_03711_, _03307_, _01830_);
  or (_03712_, _03711_, _03710_);
  and (_03713_, _03466_, _01865_);
  and (_03714_, _03568_, _01859_);
  or (_03715_, _03714_, _03713_);
  or (_03716_, _03715_, _03712_);
  or (_03717_, _03716_, _03708_);
  or (_03718_, _03717_, _03698_);
  or (_03719_, _03718_, _03695_);
  and (_03720_, _03719_, _01893_);
  and (_03721_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_03722_, _03721_, _03720_);
  or (_03723_, _03722_, _01732_);
  nand (_03725_, _01732_, _06668_);
  and (_03726_, _03725_, _05110_);
  and (_03992_, _03726_, _03723_);
  or (_03727_, _08750_, _02720_);
  or (_03728_, _08752_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_03729_, _03728_, _05110_);
  and (_03994_, _03729_, _03727_);
  and (_03730_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_03731_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_03732_, _03731_, _03730_);
  and (_03733_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_03734_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_03735_, _03734_, _03733_);
  or (_03736_, _03735_, _03732_);
  and (_03737_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_03738_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03739_, _03738_, _03737_);
  and (_03740_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_03741_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03742_, _03741_, _03740_);
  or (_03743_, _03742_, _03739_);
  or (_03744_, _03743_, _03736_);
  and (_03745_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_03746_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_03747_, _03746_, _03745_);
  and (_03749_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_03750_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_03751_, _03750_, _03749_);
  or (_03752_, _03751_, _03747_);
  and (_03753_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_03754_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_03756_, _03754_, _03753_);
  and (_03757_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_03758_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_03759_, _03758_, _03757_);
  or (_03760_, _03759_, _03756_);
  or (_03761_, _03760_, _03752_);
  or (_03762_, _03761_, _03744_);
  and (_03763_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_03764_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03765_, _03764_, _03763_);
  and (_03767_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_03768_, _01819_, _12262_);
  or (_03770_, _03768_, _03767_);
  and (_03771_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_03772_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_03773_, _03772_, _03771_);
  or (_03774_, _03773_, _03770_);
  and (_03775_, _03340_, _01853_);
  and (_03776_, _03323_, _01830_);
  or (_03777_, _03776_, _03775_);
  and (_03778_, _03577_, _01859_);
  and (_03779_, _03470_, _01865_);
  or (_03780_, _03779_, _03778_);
  or (_03781_, _03780_, _03777_);
  or (_03782_, _03781_, _03774_);
  or (_03783_, _03782_, _03765_);
  or (_03784_, _03783_, _03762_);
  and (_03785_, _03784_, _01893_);
  and (_03786_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or (_03787_, _03786_, _03785_);
  or (_03788_, _03787_, _01732_);
  nand (_03789_, _01732_, _07337_);
  and (_03790_, _03789_, _05110_);
  and (_03996_, _03790_, _03788_);
  and (_03791_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_03792_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or (_03793_, _03792_, _03791_);
  and (_03999_, _03793_, _05110_);
  and (_03794_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_03795_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or (_03796_, _03795_, _03794_);
  and (_04001_, _03796_, _05110_);
  or (_03798_, _01892_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_03799_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_03800_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_03801_, _03800_, _03799_);
  and (_03802_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_03803_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_03804_, _03803_, _03802_);
  or (_03805_, _03804_, _03801_);
  and (_03806_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_03807_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03808_, _03807_, _03806_);
  and (_03809_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_03810_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_03811_, _03810_, _03809_);
  or (_03812_, _03811_, _03808_);
  or (_03813_, _03812_, _03805_);
  and (_03814_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_03815_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_03816_, _03815_, _03814_);
  and (_03817_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_03818_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_03819_, _03818_, _03817_);
  or (_03820_, _03819_, _03816_);
  and (_03821_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_03822_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_03823_, _03822_, _03821_);
  and (_03824_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_03825_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_03826_, _03825_, _03824_);
  or (_03827_, _03826_, _03823_);
  or (_03828_, _03827_, _03820_);
  or (_03829_, _03828_, _03813_);
  and (_03830_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_03831_, _01819_, _11890_);
  or (_03833_, _03831_, _03830_);
  and (_03835_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_03836_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_03837_, _03836_, _03835_);
  or (_03838_, _03837_, _03833_);
  and (_03839_, _03299_, _01830_);
  and (_03840_, _03355_, _01853_);
  or (_03841_, _03840_, _03839_);
  and (_03842_, _03484_, _01865_);
  and (_03843_, _03583_, _01859_);
  or (_03844_, _03843_, _03842_);
  or (_03845_, _03844_, _03841_);
  or (_03846_, _03845_, _03838_);
  and (_03847_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03848_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_03850_, _03848_, _03847_);
  or (_03851_, _03850_, _03846_);
  or (_03852_, _03851_, _03829_);
  and (_03853_, _03852_, _01887_);
  and (_03854_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_03855_, _03854_, _03853_);
  and (_03856_, _03855_, _03798_);
  or (_03858_, _03856_, _01732_);
  nand (_03859_, _01732_, _06548_);
  and (_03860_, _03859_, _05110_);
  and (_04003_, _03860_, _03858_);
  and (_03861_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03862_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_03863_, _03862_, _03861_);
  and (_03864_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_03865_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_03867_, _03865_, _03864_);
  or (_03869_, _03867_, _03863_);
  and (_03870_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03871_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_03872_, _03871_, _03870_);
  and (_03873_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_03874_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_03875_, _03874_, _03873_);
  or (_03876_, _03875_, _03872_);
  or (_03878_, _03876_, _03869_);
  and (_03879_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_03880_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_03881_, _03880_, _03879_);
  and (_03882_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_03883_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_03884_, _03883_, _03882_);
  or (_03885_, _03884_, _03881_);
  and (_03886_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_03887_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_03888_, _03887_, _03886_);
  and (_03889_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_03890_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_03891_, _03890_, _03889_);
  or (_03892_, _03891_, _03888_);
  or (_03893_, _03892_, _03885_);
  or (_03894_, _03893_, _03878_);
  and (_03896_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03897_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_03898_, _03897_, _03896_);
  and (_03900_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03901_, _01819_, _11954_);
  or (_03902_, _03901_, _03900_);
  and (_03903_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_03904_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_03905_, _03904_, _03903_);
  or (_03906_, _03905_, _03902_);
  and (_03908_, _03347_, _01853_);
  and (_03909_, _03314_, _01830_);
  or (_03911_, _03909_, _03908_);
  and (_03913_, _03560_, _01859_);
  and (_03915_, _03480_, _01865_);
  or (_03916_, _03915_, _03913_);
  or (_03917_, _03916_, _03911_);
  or (_03918_, _03917_, _03906_);
  or (_03920_, _03918_, _03898_);
  or (_03921_, _03920_, _03894_);
  and (_03922_, _03921_, _01893_);
  and (_03923_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_03924_, _03923_, _03922_);
  or (_03925_, _03924_, _01732_);
  nand (_03926_, _01732_, _07235_);
  and (_03927_, _03926_, _05110_);
  and (_04065_, _03927_, _03925_);
  and (_03928_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_03930_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or (_03931_, _03930_, _03928_);
  and (_04067_, _03931_, _05110_);
  and (_03932_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_03933_, pc_log_change, _02462_);
  or (_03934_, _03933_, _03932_);
  and (_04070_, _03934_, _05110_);
  and (_03935_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_03936_, pc_log_change, _02373_);
  or (_03937_, _03936_, _03935_);
  and (_04112_, _03937_, _05110_);
  and (_03938_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_03939_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or (_03940_, _03939_, _03938_);
  and (_04114_, _03940_, _05110_);
  and (_03941_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_03942_, pc_log_change, _02377_);
  or (_03943_, _03942_, _03941_);
  and (_04166_, _03943_, _05110_);
  not (_03944_, cy_reg);
  and (_03945_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_03946_, _03945_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_03947_, _03946_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand (_03948_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_03949_, _03948_, _05482_);
  or (_03951_, _03949_, _00664_);
  and (_03952_, _03951_, _03947_);
  or (_03953_, _03952_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_03954_, _03945_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_03955_, _03954_, _03949_);
  and (_03956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _07627_);
  not (_03957_, _03956_);
  and (_03958_, _03957_, _03955_);
  nand (_03959_, _03958_, _03953_);
  not (_03960_, _03955_);
  or (_03961_, _03952_, _07604_);
  nand (_03962_, _03952_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand (_03963_, _03962_, _03961_);
  nand (_03964_, _03963_, _03960_);
  nand (_03965_, _03964_, _03959_);
  nor (_03966_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand (_03967_, _03966_, _03965_);
  or (_03968_, _03952_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_03969_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02468_);
  or (_03970_, _00664_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_03971_, _03970_, _03969_);
  and (_03973_, _03971_, _03968_);
  nand (_03974_, _03951_, _03947_);
  or (_03975_, _03974_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_03976_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_03977_, _03976_, _03945_);
  and (_03978_, _03977_, _03975_);
  or (_03979_, _03978_, _03973_);
  and (_03980_, _03979_, _03955_);
  or (_03981_, _03952_, _07666_);
  nand (_03982_, _03952_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_03983_, _03982_, _03981_);
  and (_03984_, _03983_, _03946_);
  not (_03986_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_03987_, _03952_, _03986_);
  or (_03988_, _03974_, _08206_);
  nand (_03989_, _03988_, _03987_);
  not (_03990_, _03969_);
  nor (_03991_, _03990_, _03955_);
  and (_03993_, _03991_, _03989_);
  or (_03995_, _03993_, _03984_);
  nor (_03997_, _03995_, _03980_);
  and (_03998_, _02381_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_04000_, _03974_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_04002_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_04004_, _04002_);
  and (_04005_, _04004_, _03955_);
  nand (_04006_, _04005_, _04000_);
  or (_04007_, _03952_, _07638_);
  nand (_04008_, _03952_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand (_04009_, _04008_, _04007_);
  nand (_04010_, _04009_, _03960_);
  nand (_04011_, _04010_, _04006_);
  nand (_04012_, _04011_, _03998_);
  and (_04013_, _04012_, _03997_);
  and (_04014_, _04013_, _03967_);
  and (_04015_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04016_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_04017_, _04016_, _04015_);
  and (_04018_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_04019_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_04020_, _04019_, _04018_);
  and (_04021_, _04020_, _04017_);
  and (_04022_, _04021_, _03960_);
  and (_04023_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04024_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_04025_, _04024_, _04023_);
  and (_04026_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_04027_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_04028_, _04027_, _04026_);
  and (_04029_, _04028_, _04025_);
  and (_04030_, _04029_, _03955_);
  or (_04031_, _04030_, _03952_);
  nor (_04032_, _04031_, _04022_);
  and (_04033_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04034_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_04035_, _04034_, _04033_);
  and (_04036_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_04037_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_04038_, _04037_, _04036_);
  and (_04039_, _04038_, _04035_);
  nor (_04040_, _04039_, _03955_);
  and (_04041_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04042_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_04043_, _04042_, _04041_);
  and (_04044_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_04045_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_04046_, _04045_, _04044_);
  and (_04047_, _04046_, _04043_);
  nor (_04048_, _04047_, _03960_);
  or (_04049_, _04048_, _04040_);
  and (_04050_, _04049_, _03952_);
  nor (_04051_, _04050_, _04032_);
  nor (_04052_, _04051_, _04014_);
  and (_04053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04054_, _04053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04055_, _04054_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_04056_, _04055_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_04057_, _04056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_04058_, _04057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_04059_, _04058_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_04060_, _04059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_04061_, _04060_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_04062_, _04061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_04063_, _04062_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_04064_, _04063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_04066_, _04064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04068_, _04064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04069_, _04068_, _04066_);
  and (_04071_, _04069_, _04052_);
  nor (_04072_, _04063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_04073_, _04072_, _04064_);
  and (_04074_, _04073_, _04052_);
  nor (_04075_, _04073_, _04052_);
  nor (_04076_, _04075_, _04074_);
  not (_04077_, _04076_);
  nor (_04078_, _04061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04079_, _04078_, _04062_);
  and (_04080_, _04079_, _04052_);
  nor (_04081_, _04060_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_04082_, _04081_, _04061_);
  and (_04083_, _04082_, _04052_);
  and (_04084_, _04083_, _13096_);
  nor (_04085_, _04084_, _04080_);
  nor (_04086_, _04079_, _04052_);
  nor (_04087_, _04086_, _04080_);
  not (_04088_, _04087_);
  nor (_04089_, _04082_, _04052_);
  nor (_04090_, _04089_, _04083_);
  nor (_04091_, _04059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_04092_, _04091_, _04060_);
  and (_04093_, _04092_, _04052_);
  nor (_04094_, _04058_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_04095_, _04094_, _04059_);
  and (_04096_, _04095_, _04052_);
  nor (_04097_, _04096_, _04093_);
  nor (_04098_, _04092_, _04052_);
  nor (_04099_, _04098_, _04093_);
  not (_04100_, _04099_);
  nor (_04101_, _04057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_04102_, _04101_, _04058_);
  and (_04103_, _04102_, _04052_);
  nor (_04104_, _04102_, _04052_);
  and (_04105_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_04106_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_04107_, _04106_, _04105_);
  and (_04108_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_04109_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_04110_, _04109_, _04108_);
  and (_04111_, _04110_, _04107_);
  and (_04113_, _04111_, _03960_);
  and (_04115_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04116_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_04117_, _04116_, _04115_);
  and (_04118_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04119_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_04120_, _04119_, _04118_);
  and (_04121_, _04120_, _04117_);
  and (_04122_, _04121_, _03955_);
  or (_04123_, _04122_, _03952_);
  nor (_04124_, _04123_, _04113_);
  and (_04125_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_04126_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_04127_, _04126_, _04125_);
  and (_04128_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_04129_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_04130_, _04129_, _04128_);
  and (_04131_, _04130_, _04127_);
  and (_04132_, _04131_, _03960_);
  and (_04133_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04134_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_04135_, _04134_, _04133_);
  and (_04136_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_04137_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_04138_, _04137_, _04136_);
  and (_04139_, _04138_, _04135_);
  and (_04140_, _04139_, _03955_);
  or (_04141_, _04140_, _03974_);
  nor (_04142_, _04141_, _04132_);
  nor (_04143_, _04142_, _04124_);
  nor (_04144_, _04143_, _04014_);
  nor (_04145_, _04056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_04146_, _04145_, _04057_);
  and (_04147_, _04146_, _04144_);
  nor (_04148_, _04146_, _04144_);
  nor (_04149_, _04148_, _04147_);
  and (_04150_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_04151_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_04152_, _04151_, _04150_);
  and (_04153_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_04154_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_04155_, _04154_, _04153_);
  and (_04156_, _04155_, _04152_);
  and (_04157_, _04156_, _03960_);
  and (_04158_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_04159_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_04160_, _04159_, _04158_);
  and (_04161_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_04162_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_04163_, _04162_, _04161_);
  and (_04164_, _04163_, _04160_);
  and (_04165_, _04164_, _03955_);
  or (_04167_, _04165_, _03952_);
  nor (_04168_, _04167_, _04157_);
  and (_04169_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_04170_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_04171_, _04170_, _04169_);
  and (_04172_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_04173_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_04174_, _04173_, _04172_);
  and (_04175_, _04174_, _04171_);
  and (_04176_, _04175_, _03960_);
  and (_04177_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_04178_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_04179_, _04178_, _04177_);
  and (_04180_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_04181_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_04182_, _04181_, _04180_);
  and (_04183_, _04182_, _04179_);
  and (_04184_, _04183_, _03955_);
  or (_04186_, _04184_, _03974_);
  nor (_04187_, _04186_, _04176_);
  nor (_04188_, _04187_, _04168_);
  nor (_04189_, _04188_, _04014_);
  nor (_04190_, _04055_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_04191_, _04190_, _04056_);
  and (_04192_, _04191_, _04189_);
  nor (_04193_, _04191_, _04189_);
  nor (_04194_, _04193_, _04192_);
  and (_04195_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_04196_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_04197_, _04196_, _04195_);
  and (_04198_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_04199_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_04200_, _04199_, _04198_);
  and (_04201_, _04200_, _04197_);
  and (_04202_, _04201_, _03960_);
  and (_04203_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_04204_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_04205_, _04204_, _04203_);
  and (_04206_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_04207_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_04208_, _04207_, _04206_);
  and (_04209_, _04208_, _04205_);
  and (_04210_, _04209_, _03955_);
  or (_04211_, _04210_, _03952_);
  nor (_04212_, _04211_, _04202_);
  and (_04213_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04214_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_04215_, _04214_, _04213_);
  and (_04216_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04217_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_04218_, _04217_, _04216_);
  and (_04219_, _04218_, _04215_);
  and (_04220_, _04219_, _03955_);
  and (_04221_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04222_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_04223_, _04222_, _04221_);
  and (_04224_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_04225_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_04226_, _04225_, _04224_);
  and (_04227_, _04226_, _04223_);
  and (_04228_, _04227_, _03960_);
  nor (_04229_, _04228_, _04220_);
  and (_04230_, _04229_, _03952_);
  nor (_04231_, _04230_, _04212_);
  nor (_04232_, _04231_, _04014_);
  nor (_04233_, _04054_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_04234_, _04233_, _04055_);
  and (_04235_, _04234_, _04232_);
  and (_04236_, _04235_, _04194_);
  nor (_04237_, _04236_, _04192_);
  and (_04238_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_04239_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_04240_, _04239_, _04238_);
  and (_04241_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_04242_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_04243_, _04242_, _04241_);
  and (_04244_, _04243_, _04240_);
  and (_04245_, _04244_, _03960_);
  and (_04246_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_04247_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_04248_, _04247_, _04246_);
  and (_04249_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_04250_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_04251_, _04250_, _04249_);
  and (_04252_, _04251_, _04248_);
  and (_04253_, _04252_, _03955_);
  or (_04254_, _04253_, _03952_);
  nor (_04255_, _04254_, _04245_);
  and (_04256_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_04257_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_04258_, _04257_, _04256_);
  and (_04259_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_04260_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_04261_, _04260_, _04259_);
  and (_04262_, _04261_, _04258_);
  nor (_04263_, _04262_, _03955_);
  and (_04264_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_04265_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_04266_, _04265_, _04264_);
  and (_04267_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_04268_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_04269_, _04268_, _04267_);
  and (_04270_, _04269_, _04266_);
  nor (_04271_, _04270_, _03960_);
  or (_04272_, _04271_, _04263_);
  and (_04273_, _04272_, _03952_);
  nor (_04274_, _04273_, _04255_);
  nor (_04275_, _04274_, _04014_);
  nor (_04276_, _04053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04277_, _04276_, _04054_);
  nand (_04278_, _04277_, _04275_);
  or (_04279_, _04277_, _04275_);
  and (_04280_, _04279_, _04278_);
  not (_04281_, _04280_);
  and (_04282_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _05482_);
  and (_04283_, _02468_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04284_, _04283_, _04282_);
  not (_04285_, _04284_);
  and (_04286_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_04287_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_04288_, _04287_, _04286_);
  and (_04289_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_04290_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_04291_, _04290_, _04289_);
  and (_04292_, _04291_, _04288_);
  and (_04293_, _04292_, _03960_);
  and (_04294_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_04295_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_04297_, _04295_, _04294_);
  and (_04298_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_04299_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_04300_, _04299_, _04298_);
  and (_04301_, _04300_, _04297_);
  and (_04302_, _04301_, _03955_);
  or (_04303_, _04302_, _03952_);
  nor (_04304_, _04303_, _04293_);
  and (_04305_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_04306_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_04307_, _04306_, _04305_);
  and (_04308_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_04309_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_04310_, _04309_, _04308_);
  and (_04311_, _04310_, _04307_);
  nor (_04312_, _04311_, _03955_);
  and (_04313_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_04314_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_04315_, _04314_, _04313_);
  and (_04316_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_04317_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_04318_, _04317_, _04316_);
  and (_04319_, _04318_, _04315_);
  nor (_04320_, _04319_, _03960_);
  or (_04321_, _04320_, _04312_);
  and (_04322_, _04321_, _03952_);
  nor (_04323_, _04322_, _04304_);
  nor (_04324_, _04323_, _04014_);
  nand (_04325_, _04324_, _04285_);
  not (_04326_, _04014_);
  and (_04327_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_04328_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_04329_, _04328_, _04327_);
  and (_04330_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_04331_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_04332_, _04331_, _04330_);
  and (_04333_, _04332_, _04329_);
  and (_04334_, _04333_, _03955_);
  nand (_04335_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand (_04336_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_04337_, _04336_, _04335_);
  and (_04338_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_04339_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_04340_, _04339_, _04338_);
  and (_04341_, _04340_, _04337_);
  nand (_04342_, _04341_, _03960_);
  nand (_04343_, _04342_, _03952_);
  or (_04344_, _04343_, _04334_);
  and (_04345_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_04346_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_04347_, _04346_, _04345_);
  and (_04348_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_04349_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_04350_, _04349_, _04348_);
  and (_04351_, _04350_, _04347_);
  and (_04352_, _04351_, _03955_);
  nand (_04353_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nand (_04354_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_04355_, _04354_, _04353_);
  and (_04356_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_04357_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_04358_, _04357_, _04356_);
  and (_04359_, _04358_, _04355_);
  nand (_04360_, _04359_, _03960_);
  nand (_04361_, _04360_, _03974_);
  or (_04362_, _04361_, _04352_);
  nand (_04363_, _04362_, _04344_);
  and (_04364_, _04363_, _04326_);
  nand (_04365_, _04364_, _02468_);
  and (_04366_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_04367_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_04368_, _04367_, _04366_);
  and (_04369_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_04370_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_04371_, _04370_, _04369_);
  and (_04372_, _04371_, _04368_);
  and (_04373_, _04372_, _03960_);
  and (_04374_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_04375_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_04376_, _04375_, _04374_);
  and (_04378_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_04379_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_04380_, _04379_, _04378_);
  and (_04381_, _04380_, _04376_);
  and (_04382_, _04381_, _03955_);
  or (_04383_, _04382_, _03952_);
  nor (_04384_, _04383_, _04373_);
  and (_04385_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04386_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_04387_, _04386_, _04385_);
  and (_04388_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_04389_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_04390_, _04389_, _04388_);
  and (_04391_, _04390_, _04387_);
  and (_04392_, _04391_, _03960_);
  and (_04393_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_04394_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_04395_, _04394_, _04393_);
  and (_04396_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04397_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_04398_, _04397_, _04396_);
  and (_04399_, _04398_, _04395_);
  and (_04400_, _04399_, _03955_);
  or (_04401_, _04400_, _03974_);
  nor (_04402_, _04401_, _04392_);
  nor (_04403_, _04402_, _04384_);
  nor (_04404_, _04403_, _04014_);
  and (_04405_, _04404_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_04406_, _04364_, _02468_);
  nand (_04407_, _04406_, _04365_);
  not (_04408_, _04407_);
  nand (_04409_, _04408_, _04405_);
  and (_04410_, _04409_, _04365_);
  or (_04411_, _04324_, _04285_);
  and (_04412_, _04411_, _04325_);
  not (_04413_, _04412_);
  or (_04414_, _04413_, _04410_);
  and (_04415_, _04414_, _04325_);
  or (_04416_, _04415_, _04281_);
  nand (_04417_, _04416_, _04278_);
  nor (_04418_, _04234_, _04232_);
  nor (_04419_, _04418_, _04235_);
  and (_04420_, _04419_, _04194_);
  nand (_04421_, _04420_, _04417_);
  nand (_04422_, _04421_, _04237_);
  and (_04423_, _04422_, _04149_);
  nor (_04424_, _04423_, _04147_);
  nor (_04425_, _04424_, _04104_);
  or (_04426_, _04425_, _04103_);
  nor (_04427_, _04095_, _04052_);
  nor (_04428_, _04427_, _04096_);
  nand (_04429_, _04428_, _04426_);
  or (_04430_, _04429_, _04100_);
  nand (_04431_, _04430_, _04097_);
  nand (_04432_, _04431_, _04090_);
  or (_04433_, _04432_, _04088_);
  nand (_04434_, _04433_, _04085_);
  nor (_04435_, _04062_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04436_, _04435_, _04063_);
  and (_04437_, _04436_, _04052_);
  nor (_04438_, _04436_, _04052_);
  nor (_04439_, _04438_, _04437_);
  nand (_04440_, _04439_, _04434_);
  or (_04441_, _04440_, _04077_);
  and (_04442_, _04437_, _02369_);
  nor (_04443_, _04442_, _04074_);
  nand (_04444_, _04443_, _04441_);
  nor (_04445_, _04069_, _04052_);
  nor (_04446_, _04445_, _04071_);
  and (_04447_, _04446_, _04444_);
  nor (_04448_, _04447_, _04071_);
  or (_04449_, _04066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand (_04450_, _04066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_04451_, _04450_, _04449_);
  nor (_04452_, _04451_, _04052_);
  and (_04453_, _04451_, _04052_);
  nor (_04454_, _04453_, _04452_);
  or (_04455_, _04454_, _04448_);
  nand (_04456_, _04454_, _04448_);
  and (_04457_, _04456_, _04455_);
  and (_04458_, _04457_, _03944_);
  nor (_04459_, _04451_, _03944_);
  or (_04460_, _04459_, _04458_);
  nor (_04461_, _04460_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_04462_, _04460_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_04463_, _04439_, _04434_);
  nor (_04464_, _04463_, _04437_);
  nand (_04465_, _04464_, _04077_);
  or (_04466_, _04464_, _04077_);
  nand (_04467_, _04466_, _04465_);
  and (_04468_, _04467_, _03944_);
  nor (_04469_, _04073_, _03944_);
  nor (_04470_, _04469_, _04468_);
  nor (_04471_, _04470_, _02385_);
  and (_04472_, _04470_, _02385_);
  nor (_04473_, _04079_, _03944_);
  and (_04474_, _04431_, _04090_);
  nor (_04475_, _04474_, _04083_);
  nand (_04476_, _04475_, _04088_);
  or (_04477_, _04475_, _04088_);
  nand (_04478_, _04477_, _04476_);
  and (_04479_, _04478_, _03944_);
  nor (_04480_, _04479_, _04473_);
  nor (_04481_, _04480_, _12879_);
  and (_04482_, _04480_, _12879_);
  and (_04483_, _04092_, cy_reg);
  and (_04484_, _04428_, _04426_);
  nor (_04485_, _04484_, _04096_);
  nand (_04486_, _04485_, _04099_);
  or (_04487_, _04485_, _04099_);
  nand (_04488_, _04487_, _04486_);
  and (_04489_, _04488_, _03944_);
  nor (_04490_, _04489_, _04483_);
  nor (_04491_, _04490_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_04492_, _04490_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_04493_, _04428_, _04426_);
  nand (_04494_, _04493_, _04429_);
  and (_04495_, _04494_, _03944_);
  nor (_04496_, _04095_, _03944_);
  nor (_04497_, _04496_, _04495_);
  nor (_04498_, _04497_, _02462_);
  and (_04499_, _04497_, _02462_);
  nor (_04500_, _04102_, _03944_);
  nor (_04501_, _04103_, _04104_);
  nand (_04502_, _04501_, _04424_);
  or (_04503_, _04501_, _04424_);
  and (_04504_, _04503_, _03944_);
  and (_04505_, _04504_, _04502_);
  or (_04506_, _04505_, _04500_);
  nor (_04507_, _04506_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_04508_, _04422_, _04149_);
  or (_04509_, _04508_, _04423_);
  and (_04510_, _04509_, _03944_);
  nor (_04511_, _04146_, _03944_);
  or (_04512_, _04511_, _04510_);
  nor (_04513_, _04512_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_04514_, _04235_);
  nand (_04515_, _04419_, _04417_);
  nand (_04516_, _04515_, _04514_);
  nand (_04517_, _04516_, _04194_);
  or (_04518_, _04516_, _04194_);
  nand (_04519_, _04518_, _04517_);
  and (_04520_, _04519_, _03944_);
  nor (_04521_, _04191_, _03944_);
  or (_04522_, _04521_, _04520_);
  nor (_04523_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_04524_, _04234_, cy_reg);
  or (_04525_, _04419_, _04417_);
  and (_04526_, _04525_, _04515_);
  and (_04527_, _04526_, _03944_);
  or (_04528_, _04527_, _04524_);
  and (_04529_, _04528_, _02377_);
  and (_04530_, _04277_, cy_reg);
  nand (_04531_, _04415_, _04281_);
  and (_04532_, _04531_, _04416_);
  and (_04533_, _04532_, _03944_);
  nor (_04534_, _04533_, _04530_);
  nor (_04535_, _04534_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04536_, _04284_, _03944_);
  nand (_04537_, _04413_, _04410_);
  and (_04538_, _04537_, _04414_);
  and (_04539_, _04538_, _03944_);
  nor (_04540_, _04539_, _04536_);
  nor (_04541_, _04540_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04542_, _04404_, _03944_);
  nor (_04543_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04544_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04545_, _04544_, _04543_);
  nand (_04546_, _04545_, _04542_);
  or (_04547_, _04545_, _04542_);
  and (_04548_, _04547_, _04546_);
  or (_04549_, _04548_, _04541_);
  or (_04550_, _04549_, _04535_);
  or (_04551_, _04550_, _04529_);
  or (_04552_, _04551_, _04523_);
  or (_04553_, _04552_, _04513_);
  and (_04554_, _04506_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_04555_, _04512_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_04556_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_04557_, _04528_, _02377_);
  and (_04558_, _04534_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04559_, _04540_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04560_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or (_04561_, _04408_, _04405_);
  nand (_04562_, _04561_, _04409_);
  and (_04563_, _04562_, _03944_);
  or (_04564_, _04563_, _04560_);
  nor (_04565_, _04564_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04566_, _04564_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04567_, _04566_, _04565_);
  or (_04568_, _04567_, _04559_);
  or (_04569_, _04568_, _04558_);
  or (_04570_, _04569_, _04557_);
  or (_04571_, _04570_, _04556_);
  or (_04572_, _04571_, _04555_);
  or (_04573_, _04572_, _04554_);
  or (_04574_, _04573_, _04553_);
  or (_04575_, _04574_, _04507_);
  or (_04576_, _04575_, _04499_);
  or (_04577_, _04576_, _04498_);
  or (_04578_, _04577_, _04492_);
  or (_04579_, _04578_, _04491_);
  and (_04580_, _04082_, cy_reg);
  or (_04581_, _04431_, _04090_);
  and (_04582_, _04581_, _04432_);
  and (_04583_, _04582_, _03944_);
  or (_04584_, _04583_, _04580_);
  nor (_04585_, _04584_, _02509_);
  and (_04586_, _04584_, _02509_);
  or (_04587_, _04586_, _04585_);
  or (_04588_, _04587_, _04579_);
  or (_04589_, _04588_, _04482_);
  or (_04590_, _04589_, _04481_);
  and (_04591_, _04436_, cy_reg);
  or (_04592_, _04439_, _04434_);
  and (_04593_, _04592_, _04440_);
  and (_04594_, _04593_, _03944_);
  or (_04595_, _04594_, _04591_);
  nor (_04596_, _04595_, _01639_);
  and (_04597_, _04595_, _01639_);
  or (_04598_, _04597_, _04596_);
  or (_04599_, _04598_, _04590_);
  or (_04600_, _04599_, _04472_);
  or (_04601_, _04600_, _04471_);
  and (_04602_, _04069_, cy_reg);
  nor (_04603_, _04446_, _04444_);
  nor (_04604_, _04603_, _04447_);
  and (_04605_, _04604_, _03944_);
  or (_04606_, _04605_, _04602_);
  nor (_04607_, _04606_, _00990_);
  and (_04608_, _04606_, _00990_);
  or (_04609_, _04608_, _04607_);
  or (_04610_, _04609_, _04601_);
  or (_04611_, _04610_, _04462_);
  or (_04612_, _04611_, _04461_);
  nor (_04613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_04614_, _04613_, _02396_);
  nor (_04615_, _04614_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04616_, _04614_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04617_, _04616_, _04615_);
  or (_04618_, _01339_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_04619_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04620_, _04619_, _04618_);
  or (_04621_, _04620_, _04617_);
  and (_04622_, _04613_, _02396_);
  nor (_04623_, _04622_, _04614_);
  or (_04624_, _01339_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_04625_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_04626_, _04625_, _04624_);
  and (_04627_, _04626_, _04617_);
  nor (_04628_, _04627_, _04623_);
  and (_04629_, _04628_, _04621_);
  and (_04630_, _04617_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_04631_, _02477_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_04632_, _04631_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04633_, _04632_, _04630_);
  and (_04634_, _04617_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_04635_, _02477_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_04636_, _04635_, _01339_);
  or (_04637_, _04636_, _04634_);
  and (_04638_, _04637_, _04623_);
  and (_04639_, _04638_, _04633_);
  or (_04640_, _04639_, _04629_);
  and (_04641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04642_, _04641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_04643_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_04644_, _04643_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_04645_, _04644_, _04642_);
  not (_04646_, _04645_);
  nor (_04647_, _04642_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04648_, _04642_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04649_, _04648_, _04647_);
  or (_04650_, _04649_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_04651_, _02477_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_04652_, _04651_, _04650_);
  or (_04653_, _04652_, _04646_);
  nand (_04654_, _04649_, _08206_);
  or (_04655_, _04649_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_04656_, _04655_, _04654_);
  or (_04657_, _04656_, _04645_);
  and (_04658_, _04657_, _04653_);
  or (_04659_, _04658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_04660_, _04649_, _07666_);
  and (_04661_, _04649_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_04662_, _04661_, _04660_);
  and (_04663_, _04662_, _04646_);
  or (_04664_, _04649_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_04665_, _02477_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_04666_, _04665_, _04645_);
  and (_04667_, _04666_, _04664_);
  or (_04668_, _04667_, _01339_);
  or (_04669_, _04668_, _04663_);
  or (_04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_04671_, _02477_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_04672_, _04671_, _04670_);
  or (_04673_, _04672_, _02396_);
  or (_04674_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_04675_, _02477_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_04676_, _04675_, _04674_);
  or (_04677_, _04676_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04678_, _04677_, _04673_);
  and (_04679_, _04678_, _04643_);
  and (_04680_, _01339_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_04681_, _02477_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_04682_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_04683_, _04682_, _04681_);
  or (_04684_, _04683_, _02396_);
  or (_04685_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_04686_, _02477_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_04687_, _04686_, _04685_);
  or (_04688_, _04687_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04689_, _04688_, _04684_);
  and (_04690_, _04689_, _04680_);
  or (_04691_, _04690_, _04679_);
  and (_04692_, _04678_, _01339_);
  and (_04693_, _02396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04694_, _04693_, _04683_);
  or (_04695_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_04696_, _02477_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04697_, _04696_, _04641_);
  and (_04698_, _04697_, _04695_);
  or (_04699_, _04698_, _04694_);
  or (_04700_, _04699_, _04692_);
  and (_04701_, _04700_, _04691_);
  and (_04702_, _04701_, _04669_);
  and (_04703_, _04702_, _04659_);
  and (_04704_, _04703_, _04640_);
  and (_04705_, _04617_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_04706_, _02477_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_04707_, _04706_, _04623_);
  or (_04708_, _04707_, _04705_);
  and (_04709_, _04708_, _01339_);
  nor (_04710_, _04617_, _07638_);
  and (_04711_, _04617_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_04712_, _04711_, _04710_);
  or (_04713_, _04712_, _04623_);
  and (_04714_, _04713_, _04709_);
  or (_04715_, _04714_, _04699_);
  and (_04716_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_04717_, _02477_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_04718_, _04717_, _04716_);
  and (_04719_, _04718_, _02396_);
  and (_04720_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_04721_, _04720_, _04631_);
  and (_04722_, _04721_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_04723_, _04722_, _04719_);
  and (_04724_, _04723_, _01339_);
  or (_04725_, _04649_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_04726_, _04681_, _04645_);
  and (_04727_, _04726_, _04725_);
  not (_04728_, _04649_);
  or (_04729_, _04728_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_04730_, _04649_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04731_, _04730_, _04646_);
  and (_04732_, _04731_, _04729_);
  or (_04733_, _04732_, _04727_);
  and (_04734_, _04733_, _04724_);
  or (_04735_, _04649_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_04736_, _04671_, _04645_);
  and (_04737_, _04736_, _04735_);
  or (_04738_, _04728_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_04739_, _04649_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_04740_, _04739_, _04646_);
  and (_04741_, _04740_, _04738_);
  or (_04742_, _04741_, _04737_);
  and (_04743_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_04744_, _04635_, _02396_);
  or (_04745_, _04744_, _04743_);
  or (_04746_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_04747_, _02477_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_04748_, _04747_, _04746_);
  or (_04749_, _04748_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04750_, _04749_, _04745_);
  and (_04751_, _04750_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04752_, _04721_, _04693_);
  or (_04753_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_04754_, _02477_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04755_, _04754_, _04641_);
  and (_04756_, _04755_, _04753_);
  or (_04757_, _04756_, _04752_);
  and (_04758_, _04757_, _04751_);
  and (_04759_, _04758_, _04742_);
  or (_04760_, _04759_, _04734_);
  or (_04761_, _04757_, _04750_);
  and (_04762_, _04761_, _02943_);
  and (_04763_, _04762_, _04760_);
  and (_04764_, _04763_, _04715_);
  or (_04765_, _04764_, _04704_);
  not (_04766_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_04767_, _03966_, _05482_);
  nor (_04768_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04769_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04770_, _04769_, _04768_);
  nand (_04771_, _04770_, _04766_);
  nor (_04772_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04773_, _04772_, _02381_);
  nor (_04774_, _04773_, _04767_);
  or (_04775_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_04776_, _04775_, _04774_);
  and (_04777_, _04776_, _04771_);
  not (_04778_, _04774_);
  and (_04779_, _04770_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_04780_, _04770_, _03986_);
  or (_04781_, _04780_, _04779_);
  and (_04782_, _04781_, _04778_);
  or (_04783_, _04782_, _04777_);
  and (_04784_, _04783_, _03945_);
  nand (_04785_, _04770_, _07627_);
  or (_04786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_04787_, _04786_, _04774_);
  and (_04788_, _04787_, _04785_);
  and (_04789_, _04770_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_04790_, _04770_, _07604_);
  or (_04791_, _04790_, _04789_);
  and (_04792_, _04791_, _04778_);
  or (_04793_, _04792_, _04788_);
  and (_04794_, _04793_, _03998_);
  or (_04795_, _04794_, _04784_);
  nand (_04796_, _04770_, _07647_);
  and (_04797_, _04774_, _04004_);
  and (_04798_, _04797_, _04796_);
  and (_04799_, _04770_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_04800_, _04770_, _07638_);
  or (_04801_, _04800_, _04799_);
  and (_04802_, _04801_, _04778_);
  or (_04803_, _04802_, _04798_);
  and (_04804_, _04803_, _03966_);
  nand (_04805_, _04770_, _07675_);
  and (_04806_, _04774_, _03976_);
  and (_04807_, _04806_, _04805_);
  and (_04808_, _04770_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_04809_, _04770_, _07666_);
  or (_04810_, _04809_, _04808_);
  and (_04811_, _04810_, _04778_);
  or (_04812_, _04811_, _04807_);
  and (_04813_, _04812_, _03969_);
  or (_04814_, _04813_, _04804_);
  or (_04815_, _04814_, _04795_);
  or (_04816_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand (_04817_, _04816_, _03969_);
  or (_04818_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand (_04819_, _04818_, _03998_);
  and (_04820_, _04819_, _04817_);
  or (_04821_, _03948_, _09288_);
  nand (_04822_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_04823_, _04822_, _04821_);
  and (_04824_, _04823_, _04820_);
  nand (_04825_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  or (_04826_, _03948_, _07721_);
  and (_04827_, _04826_, _04825_);
  nor (_04828_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  or (_04829_, _04828_, _03948_);
  nand (_04830_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_04831_, _04830_, _04829_);
  and (_04832_, _04831_, _04827_);
  and (_04833_, _04832_, _04824_);
  nand (_04834_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_04835_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  or (_04836_, _04835_, _03948_);
  and (_04837_, _04836_, _04834_);
  or (_04838_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_04839_, _04838_, _03969_);
  or (_04840_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand (_04841_, _04840_, _03998_);
  and (_04842_, _04841_, _04839_);
  and (_04843_, _04842_, _04837_);
  or (_04844_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand (_04845_, _04844_, _03966_);
  or (_04846_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand (_04847_, _04846_, _03966_);
  and (_04848_, _04847_, _04845_);
  nand (_04849_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nand (_04850_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_04851_, _04850_, _04849_);
  and (_04852_, _04851_, _04848_);
  and (_04853_, _04852_, _04843_);
  and (_04854_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04855_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or (_04856_, _04855_, _04854_);
  and (_04857_, _03945_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04858_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or (_04859_, _04858_, _04857_);
  or (_04860_, _04859_, _04856_);
  and (_04861_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_04862_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or (_04863_, _04862_, _04861_);
  and (_04864_, _03945_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_04865_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  or (_04866_, _04865_, _04864_);
  or (_04867_, _04866_, _04863_);
  and (_04868_, _04867_, _04860_);
  and (_04869_, _04868_, _04853_);
  and (_04870_, _04869_, _04833_);
  or (_04871_, _04870_, _05482_);
  or (_04872_, _03948_, _07716_);
  nand (_04873_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_04874_, _04873_, _04872_);
  nor (_04875_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  or (_04876_, _04875_, _03948_);
  or (_04877_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand (_04878_, _04877_, _03966_);
  and (_04879_, _04878_, _04876_);
  and (_04880_, _04879_, _04874_);
  nand (_04881_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or (_04882_, _03948_, _08830_);
  and (_04883_, _04882_, _04881_);
  or (_04884_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand (_04885_, _04884_, _03969_);
  or (_04886_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand (_04887_, _04886_, _03998_);
  and (_04888_, _04887_, _04885_);
  and (_04889_, _04888_, _04883_);
  and (_04890_, _04889_, _04880_);
  nand (_04891_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_04892_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  or (_04893_, _04892_, _03948_);
  and (_04894_, _04893_, _04891_);
  or (_04895_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_04896_, _04895_, _03969_);
  or (_04897_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand (_04898_, _04897_, _03998_);
  and (_04899_, _04898_, _04896_);
  and (_04900_, _04899_, _04894_);
  nand (_04901_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or (_04902_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand (_04903_, _04902_, _03966_);
  and (_04904_, _04903_, _04901_);
  nand (_04905_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_04906_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_04907_, _04906_, _04905_);
  and (_04908_, _04907_, _04904_);
  and (_04909_, _04908_, _04900_);
  and (_04910_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_04911_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or (_04912_, _04911_, _04910_);
  and (_04913_, _03945_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_04914_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or (_04915_, _04914_, _04913_);
  or (_04916_, _04915_, _04912_);
  and (_04917_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_04918_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or (_04919_, _04918_, _04917_);
  and (_04920_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_04921_, _03945_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  or (_04922_, _04921_, _04920_);
  or (_04923_, _04922_, _04919_);
  and (_04924_, _04923_, _04916_);
  and (_04925_, _04924_, _04909_);
  and (_04926_, _04925_, _04890_);
  or (_04927_, _04926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04928_, _04927_, _04871_);
  or (_04929_, _04928_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04930_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04931_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or (_04932_, _04931_, _04930_);
  and (_04933_, _03945_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_04934_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or (_04935_, _04934_, _04933_);
  or (_04936_, _04935_, _04932_);
  and (_04937_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_04938_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or (_04939_, _04938_, _04937_);
  and (_04940_, _03945_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_04941_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or (_04942_, _04941_, _04940_);
  or (_04943_, _04942_, _04939_);
  nand (_04944_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  or (_04945_, _03948_, _09716_);
  and (_04946_, _04945_, _04944_);
  nand (_04947_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_04948_, _04947_, _04946_);
  and (_04949_, _04948_, _04943_);
  and (_04950_, _04949_, _04936_);
  nor (_04951_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_04952_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand (_04953_, _04952_, _04951_);
  nand (_04954_, _04953_, _03998_);
  not (_04955_, _03966_);
  nor (_04956_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_04957_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_04958_, _04957_, _04956_);
  or (_04959_, _04958_, _04955_);
  nor (_04960_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_04961_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand (_04962_, _04961_, _04960_);
  nand (_04963_, _04962_, _03969_);
  and (_04964_, _04963_, _04959_);
  and (_04965_, _04964_, _04954_);
  nand (_04966_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_04967_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_04968_, _04967_, _04966_);
  or (_04969_, _03948_, _07691_);
  nand (_04970_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_04971_, _04970_, _04969_);
  and (_04972_, _04971_, _04968_);
  nor (_04973_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_04974_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_04975_, _04974_, _04973_);
  or (_04976_, _04975_, _03948_);
  nand (_04977_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_04978_, _04977_, _05482_);
  and (_04979_, _04978_, _04976_);
  and (_04980_, _04979_, _04972_);
  and (_04981_, _04980_, _04965_);
  and (_04982_, _04981_, _04950_);
  and (_04983_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04984_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or (_04985_, _04984_, _04983_);
  and (_04986_, _03945_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04987_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or (_04988_, _04987_, _04986_);
  or (_04989_, _04988_, _04985_);
  and (_04990_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_04991_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or (_04992_, _04991_, _04990_);
  and (_04993_, _03945_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04994_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or (_04995_, _04994_, _04993_);
  or (_04996_, _04995_, _04992_);
  nand (_04997_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_04998_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_04999_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_05000_, _04999_, _04998_);
  and (_05001_, _05000_, _04997_);
  and (_05002_, _05001_, _04996_);
  and (_05003_, _05002_, _04989_);
  nor (_05004_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_05005_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand (_05006_, _05005_, _05004_);
  nand (_05007_, _05006_, _03969_);
  nor (_05008_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_05009_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_05010_, _05009_, _05008_);
  or (_05011_, _05010_, _04955_);
  nor (_05012_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_05013_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_05014_, _05013_, _05012_);
  nand (_05015_, _05014_, _03998_);
  and (_05016_, _05015_, _05011_);
  and (_05017_, _05016_, _05007_);
  nand (_05018_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  or (_05019_, _03948_, _10131_);
  and (_05020_, _05019_, _05018_);
  or (_05021_, _03948_, _07684_);
  nand (_05022_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_05023_, _05022_, _05021_);
  and (_05024_, _05023_, _05020_);
  nor (_05025_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_05026_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_05027_, _05026_, _05025_);
  or (_05028_, _05027_, _03948_);
  nand (_05029_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_05030_, _05029_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05031_, _05030_, _05028_);
  and (_05032_, _05031_, _05024_);
  and (_05033_, _05032_, _05017_);
  and (_05034_, _05033_, _05003_);
  or (_05035_, _05034_, _00664_);
  or (_05036_, _05035_, _04982_);
  and (_05037_, _04775_, _03970_);
  or (_05038_, _05037_, _05482_);
  or (_05039_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05040_, _00664_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05041_, _05040_, _05039_);
  or (_05042_, _05041_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05043_, _05042_, _05038_);
  and (_05044_, _05043_, _02468_);
  or (_05045_, _00664_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05046_, _05045_, _03976_);
  and (_05047_, _05046_, _04282_);
  or (_05048_, _00664_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05049_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05050_, _05049_, _04053_);
  and (_05051_, _05050_, _05048_);
  or (_05052_, _05051_, _05047_);
  or (_05053_, _05052_, _05044_);
  and (_05054_, _05053_, _02381_);
  or (_05055_, _00664_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_05056_, _04002_, _05482_);
  and (_05057_, _05056_, _05055_);
  or (_05058_, _00664_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05060_, _05059_, _05482_);
  and (_05061_, _05060_, _05058_);
  or (_05062_, _05061_, _05057_);
  and (_05063_, _05062_, _03969_);
  or (_05064_, _00664_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05065_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05066_, _05065_, _05064_);
  and (_05067_, _05066_, _03946_);
  and (_05068_, _03945_, _05482_);
  and (_05069_, _04786_, _03957_);
  and (_05070_, _05069_, _05068_);
  or (_05071_, _05070_, _05067_);
  or (_05072_, _05071_, _05063_);
  and (_05073_, _05062_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05074_, _05069_, _04283_);
  or (_05075_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05076_, _00664_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05077_, _05076_, _05075_);
  and (_05078_, _05077_, _04772_);
  or (_05079_, _05078_, _02381_);
  or (_05080_, _05079_, _05074_);
  or (_05081_, _05080_, _05073_);
  and (_05082_, _05081_, _05072_);
  or (_05083_, _05082_, _05054_);
  and (_05084_, _05043_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05085_, _05046_, _04283_);
  and (_05086_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05087_, _00664_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05088_, _05087_, _05086_);
  and (_05089_, _05088_, _04772_);
  or (_05090_, _05089_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_05091_, _05090_, _05085_);
  or (_05092_, _05091_, _05084_);
  nor (_05093_, _02505_, first_instr);
  and (_05094_, _05093_, _05092_);
  and (_05095_, _05094_, _05083_);
  and (_05096_, _05095_, _05036_);
  and (_05097_, _05096_, _04929_);
  and (_05098_, _05097_, _04326_);
  and (_05099_, _05098_, _04815_);
  and (_05100_, _05099_, _04765_);
  and (property_invalid_jnc, _05100_, _04612_);
  and (_05101_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_05102_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or (_05103_, _05102_, _05101_);
  and (_04185_, _05103_, _05110_);
  or (_05104_, pc_log_change_r, _03944_);
  nand (_05105_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_00000_, _05105_, _05104_);
  and (_05106_, _02505_, first_instr);
  or (_00001_, _05106_, rst);
  dff (cy_reg, _00000_);
  dff (pc_log_change_r, pc_log_change);
  dff (first_instr, _00001_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _08906_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _08909_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _08913_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _08916_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _08920_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _08923_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _08926_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _06039_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _08823_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _08826_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _08829_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _08832_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _08835_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _08839_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _08843_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _08846_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _13437_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _13438_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _13439_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _08744_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _13440_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _13441_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _13442_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _13443_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _08636_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _08640_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _08645_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _08650_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _13433_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _13434_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _13435_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _13436_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _08550_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _08552_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _08556_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _08559_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _08562_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _08566_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _08568_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _08571_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _08465_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _08468_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _08472_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _08475_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _08477_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _08479_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _08482_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _08485_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _08374_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _08377_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _08382_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _08386_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _08389_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _08392_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _08396_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _08399_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _13449_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _08271_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _08275_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _08279_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _08284_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _08289_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _08295_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _08299_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _08171_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _08175_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _13444_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _13445_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _13446_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _13447_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _13448_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _08185_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _08077_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _08080_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _08084_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _08089_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _08091_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _08094_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _08098_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _08103_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _07991_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _07994_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _07997_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _08000_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _08003_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _08006_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _08009_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _08012_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _07573_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _07577_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _07581_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _07584_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _07587_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _07590_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _07593_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _07597_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _07468_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _07472_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _07476_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _07481_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _07484_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _07488_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _07491_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _07495_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _07792_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _07795_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _07798_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _07803_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _07807_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _07812_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _07817_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _07822_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _07686_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _07689_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _07692_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _07697_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _07700_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _07703_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _07708_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _07713_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _07911_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _07915_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _07919_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _07922_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _07924_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _07928_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _07932_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _07934_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _06060_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _06090_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _06133_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _06181_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _06236_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _06299_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _06361_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _06441_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _06527_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _06614_);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _06715_);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _06806_);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _06900_);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _06995_);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _07112_);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _06013_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _05695_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _05698_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _05701_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _05704_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _05706_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _05709_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _05712_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _05565_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _10979_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _05721_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _05724_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _05727_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _05730_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _05733_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _12746_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _05745_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _05748_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _05750_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _12081_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _05757_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _05569_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _11725_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12506_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _11704_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _12511_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _05342_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _11694_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _05315_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _11718_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _05525_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _09737_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09877_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09900_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09902_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09897_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09905_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _02086_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _11679_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _02048_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _01001_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _02391_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05179_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _02587_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _02607_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05205_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _02812_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _02814_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05208_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _02848_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05331_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _02875_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _02881_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _02894_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _05477_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _02940_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05430_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _05513_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03919_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _02218_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _11913_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _03950_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _05107_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _04296_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _02925_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _02917_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _02738_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _02207_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _07166_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _02222_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _04377_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _01746_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _01905_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _02906_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03907_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _03222_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _05108_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _02954_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03985_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _02578_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _03057_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _01604_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03033_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _06408_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _06372_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _06192_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _06684_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _02543_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _03972_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _02970_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _03316_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _08933_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _10862_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _00018_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _00921_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _05289_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _02820_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _02963_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _13169_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _07653_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _00648_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _07648_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _03755_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _03534_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _03663_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _01577_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _05173_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _07639_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _03709_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _07665_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _05161_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _10144_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01540_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _07102_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _05428_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _12941_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _13173_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _12945_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _12614_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _12886_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _06855_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _11392_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _01561_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _01531_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _00824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _00590_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _10714_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _03670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _01646_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _02780_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _02837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _04166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _02776_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _04112_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _04070_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02774_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _02863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _11004_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _03868_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _02771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _00915_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _13027_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02828_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _06919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _00377_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _02762_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _06782_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _10427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _02759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _02825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _02850_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _02861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _11702_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _02010_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _02755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _03660_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _13022_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _10724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _10883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _11198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _02834_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _02255_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _13108_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _11991_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _08747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _08380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _12124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _03849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _03001_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _11980_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _10720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _03895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _03914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03912_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _03910_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _03899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _12019_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _04185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _04114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _04067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _04001_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _03999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _12015_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _10717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _10880_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _10935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _03834_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _03857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _02885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _02948_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _03089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _03075_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _03073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03064_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _12047_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _03203_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _03198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _10712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _12055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03101_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _12593_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _10813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _10803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _00796_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _00792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _00785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _00769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _00767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _12143_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _00933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _00931_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _00884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _00871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12139_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _10697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _00483_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _00467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _00462_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _10789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _00253_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _00306_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _00302_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _00273_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _12157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _10679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _11164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _11210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _12202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _00004_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _00038_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _00035_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _00028_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _10784_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _10517_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _10562_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _10567_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12107_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _12079_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12076_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12069_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _12685_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _12644_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _10558_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _11739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _10539_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _10663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11534_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11531_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _11522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _12600_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _12582_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _12721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _11496_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _10654_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _10641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _10620_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _11514_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _11509_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _11126_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03099_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _11624_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _11121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _11229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11270_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11649_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _11643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _11115_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11659_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _11112_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _11224_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11674_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11668_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _11697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _11095_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _11221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _11267_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _11291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _11364_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _11390_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11375_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11244_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11318_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _11154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _11278_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _11413_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _10400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03108_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _10460_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _11285_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _11947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _11940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _10472_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _02407_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _03724_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _03769_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _03866_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _03706_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _03797_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _02476_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _03748_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _03766_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _03996_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _03992_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _04065_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _04003_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03684_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _02423_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _03704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _06484_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _03877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _07042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _03832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _03309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _06474_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _05109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _05360_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _13347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _02466_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _13360_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _13357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _02463_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _13307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _13293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _05691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _05688_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _05680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _05657_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _05665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _01636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _05775_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _01593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07867_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _05780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _05772_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _01615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _05783_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _01669_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _08294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _01574_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _01571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _01479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _01590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _01581_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _01478_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _01520_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _08055_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _01475_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _03130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _07918_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _01527_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _01756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _10256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _01759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _01471_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _10385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _01763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _01767_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _09243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _07655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _07357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _01522_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _01567_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _01565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _07249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _01795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _01465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _01801_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _01799_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _01463_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _01516_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _01804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _01812_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _01460_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _01826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _01822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _01459_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _01494_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _01845_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _10406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _02525_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _02565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _02559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _01488_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _02522_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _02557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _02698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _02553_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02520_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _02921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _02696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02666_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _02656_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _02655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _02549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02518_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _02704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _03593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02671_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _02668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _02547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _02677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _09234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _01741_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _09629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _09639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _09636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _09633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03196_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _12852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _12846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _12842_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _12840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _02602_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _12781_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _12774_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _02472_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _13155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00411_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00422_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _12133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _12136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _12116_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _12113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _12110_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _12122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _12085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _00415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _12152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _12155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _12170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _12161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _12164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _12238_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _00419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _00417_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _00383_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12199_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _12196_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12251_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _12244_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _12247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _00387_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _12320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _12331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _12335_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _12296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _12293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _00385_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _00399_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12375_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _12366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _12372_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _12391_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _12383_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _12388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00395_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01940_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01931_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _05216_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _12309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _12306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _12302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _12299_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _07864_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _12342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _12271_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _12267_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _07878_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _11138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _12206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _07900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _12218_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _01752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _09843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _10730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _10755_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _10746_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _10739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _10736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _10660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _10649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _10645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _12226_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _10684_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _10709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _10705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _10524_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _12261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _10600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _10597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _10587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _10585_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _10582_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _03173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _03170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _03167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _03165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _03153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _03151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _03149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _03147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _03145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _03143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _03135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _03191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _09231_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _10104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _01600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _03686_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _03659_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _03599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _03114_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _03571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _03994_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _07758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01619_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _03532_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _03112_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _02503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01513_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01500_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01498_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01447_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _08247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _03193_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _03186_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _03155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _03085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _03059_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _07189_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _07175_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _08250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02897_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _10942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _07036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _10974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _10966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _11006_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _10985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _11161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _11073_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _12398_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _11983_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _02878_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _00031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _12951_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _00263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _00128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _06965_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _00472_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _00451_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _02688_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01043_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _00929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _06961_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01468_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01453_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _07022_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _07047_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02626_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [8], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [9], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [10], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [11], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [12], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [13], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [14], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [15], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [16], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [0], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [1], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [2], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [3], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [4], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [5], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [6], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [7], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [0], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [1], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [2], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [3], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [4], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [5], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [6], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [7], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.mulOv , ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [0], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [1], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [2], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [3], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [4], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [5], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [6], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [7], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_alu1.divOv , ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.ABINPUT000 [0], ABINPUT000[0]);
  buf(\oc8051_top_1.ABINPUT000 [1], ABINPUT000[1]);
  buf(\oc8051_top_1.ABINPUT000 [2], ABINPUT000[2]);
  buf(\oc8051_top_1.ABINPUT000 [3], ABINPUT000[3]);
  buf(\oc8051_top_1.ABINPUT000 [4], ABINPUT000[4]);
  buf(\oc8051_top_1.ABINPUT000 [5], ABINPUT000[5]);
  buf(\oc8051_top_1.ABINPUT000 [6], ABINPUT000[6]);
  buf(\oc8051_top_1.ABINPUT000 [7], ABINPUT000[7]);
  buf(\oc8051_top_1.ABINPUT000 [8], ABINPUT000[8]);
  buf(\oc8051_top_1.ABINPUT000 [9], ABINPUT000[9]);
  buf(\oc8051_top_1.ABINPUT000 [10], ABINPUT000[10]);
  buf(\oc8051_top_1.ABINPUT000 [11], ABINPUT000[11]);
  buf(\oc8051_top_1.ABINPUT000 [12], ABINPUT000[12]);
  buf(\oc8051_top_1.ABINPUT000 [13], ABINPUT000[13]);
  buf(\oc8051_top_1.ABINPUT000 [14], ABINPUT000[14]);
  buf(\oc8051_top_1.ABINPUT000 [15], ABINPUT000[15]);
  buf(\oc8051_top_1.ABINPUT000 [16], ABINPUT000[16]);
  buf(\oc8051_top_1.ABINPUT000000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.ABINPUT000000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.ABINPUT000000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.ABINPUT000000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.ABINPUT000000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.ABINPUT000000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.ABINPUT000000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.ABINPUT000000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.ABINPUT000000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.ABINPUT000000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.ABINPUT000000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.ABINPUT000000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.ABINPUT000000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.ABINPUT000000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.ABINPUT000000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.ABINPUT000000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.ABINPUT000000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
